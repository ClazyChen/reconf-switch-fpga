module Parser(
  input         clock,
  input  [7:0]  io_pipe_phv_in_data_0,
  input  [7:0]  io_pipe_phv_in_data_1,
  input  [7:0]  io_pipe_phv_in_data_2,
  input  [7:0]  io_pipe_phv_in_data_3,
  input  [7:0]  io_pipe_phv_in_data_4,
  input  [7:0]  io_pipe_phv_in_data_5,
  input  [7:0]  io_pipe_phv_in_data_6,
  input  [7:0]  io_pipe_phv_in_data_7,
  input  [7:0]  io_pipe_phv_in_data_8,
  input  [7:0]  io_pipe_phv_in_data_9,
  input  [7:0]  io_pipe_phv_in_data_10,
  input  [7:0]  io_pipe_phv_in_data_11,
  input  [7:0]  io_pipe_phv_in_data_12,
  input  [7:0]  io_pipe_phv_in_data_13,
  input  [7:0]  io_pipe_phv_in_data_14,
  input  [7:0]  io_pipe_phv_in_data_15,
  input  [7:0]  io_pipe_phv_in_data_16,
  input  [7:0]  io_pipe_phv_in_data_17,
  input  [7:0]  io_pipe_phv_in_data_18,
  input  [7:0]  io_pipe_phv_in_data_19,
  input  [7:0]  io_pipe_phv_in_data_20,
  input  [7:0]  io_pipe_phv_in_data_21,
  input  [7:0]  io_pipe_phv_in_data_22,
  input  [7:0]  io_pipe_phv_in_data_23,
  input  [7:0]  io_pipe_phv_in_data_24,
  input  [7:0]  io_pipe_phv_in_data_25,
  input  [7:0]  io_pipe_phv_in_data_26,
  input  [7:0]  io_pipe_phv_in_data_27,
  input  [7:0]  io_pipe_phv_in_data_28,
  input  [7:0]  io_pipe_phv_in_data_29,
  input  [7:0]  io_pipe_phv_in_data_30,
  input  [7:0]  io_pipe_phv_in_data_31,
  input  [7:0]  io_pipe_phv_in_data_32,
  input  [7:0]  io_pipe_phv_in_data_33,
  input  [7:0]  io_pipe_phv_in_data_34,
  input  [7:0]  io_pipe_phv_in_data_35,
  input  [7:0]  io_pipe_phv_in_data_36,
  input  [7:0]  io_pipe_phv_in_data_37,
  input  [7:0]  io_pipe_phv_in_data_38,
  input  [7:0]  io_pipe_phv_in_data_39,
  input  [7:0]  io_pipe_phv_in_data_40,
  input  [7:0]  io_pipe_phv_in_data_41,
  input  [7:0]  io_pipe_phv_in_data_42,
  input  [7:0]  io_pipe_phv_in_data_43,
  input  [7:0]  io_pipe_phv_in_data_44,
  input  [7:0]  io_pipe_phv_in_data_45,
  input  [7:0]  io_pipe_phv_in_data_46,
  input  [7:0]  io_pipe_phv_in_data_47,
  input  [7:0]  io_pipe_phv_in_data_48,
  input  [7:0]  io_pipe_phv_in_data_49,
  input  [7:0]  io_pipe_phv_in_data_50,
  input  [7:0]  io_pipe_phv_in_data_51,
  input  [7:0]  io_pipe_phv_in_data_52,
  input  [7:0]  io_pipe_phv_in_data_53,
  input  [7:0]  io_pipe_phv_in_data_54,
  input  [7:0]  io_pipe_phv_in_data_55,
  input  [7:0]  io_pipe_phv_in_data_56,
  input  [7:0]  io_pipe_phv_in_data_57,
  input  [7:0]  io_pipe_phv_in_data_58,
  input  [7:0]  io_pipe_phv_in_data_59,
  input  [7:0]  io_pipe_phv_in_data_60,
  input  [7:0]  io_pipe_phv_in_data_61,
  input  [7:0]  io_pipe_phv_in_data_62,
  input  [7:0]  io_pipe_phv_in_data_63,
  input  [7:0]  io_pipe_phv_in_data_64,
  input  [7:0]  io_pipe_phv_in_data_65,
  input  [7:0]  io_pipe_phv_in_data_66,
  input  [7:0]  io_pipe_phv_in_data_67,
  input  [7:0]  io_pipe_phv_in_data_68,
  input  [7:0]  io_pipe_phv_in_data_69,
  input  [7:0]  io_pipe_phv_in_data_70,
  input  [7:0]  io_pipe_phv_in_data_71,
  input  [7:0]  io_pipe_phv_in_data_72,
  input  [7:0]  io_pipe_phv_in_data_73,
  input  [7:0]  io_pipe_phv_in_data_74,
  input  [7:0]  io_pipe_phv_in_data_75,
  input  [7:0]  io_pipe_phv_in_data_76,
  input  [7:0]  io_pipe_phv_in_data_77,
  input  [7:0]  io_pipe_phv_in_data_78,
  input  [7:0]  io_pipe_phv_in_data_79,
  input  [7:0]  io_pipe_phv_in_data_80,
  input  [7:0]  io_pipe_phv_in_data_81,
  input  [7:0]  io_pipe_phv_in_data_82,
  input  [7:0]  io_pipe_phv_in_data_83,
  input  [7:0]  io_pipe_phv_in_data_84,
  input  [7:0]  io_pipe_phv_in_data_85,
  input  [7:0]  io_pipe_phv_in_data_86,
  input  [7:0]  io_pipe_phv_in_data_87,
  input  [7:0]  io_pipe_phv_in_data_88,
  input  [7:0]  io_pipe_phv_in_data_89,
  input  [7:0]  io_pipe_phv_in_data_90,
  input  [7:0]  io_pipe_phv_in_data_91,
  input  [7:0]  io_pipe_phv_in_data_92,
  input  [7:0]  io_pipe_phv_in_data_93,
  input  [7:0]  io_pipe_phv_in_data_94,
  input  [7:0]  io_pipe_phv_in_data_95,
  input  [7:0]  io_pipe_phv_in_data_96,
  input  [7:0]  io_pipe_phv_in_data_97,
  input  [7:0]  io_pipe_phv_in_data_98,
  input  [7:0]  io_pipe_phv_in_data_99,
  input  [7:0]  io_pipe_phv_in_data_100,
  input  [7:0]  io_pipe_phv_in_data_101,
  input  [7:0]  io_pipe_phv_in_data_102,
  input  [7:0]  io_pipe_phv_in_data_103,
  input  [7:0]  io_pipe_phv_in_data_104,
  input  [7:0]  io_pipe_phv_in_data_105,
  input  [7:0]  io_pipe_phv_in_data_106,
  input  [7:0]  io_pipe_phv_in_data_107,
  input  [7:0]  io_pipe_phv_in_data_108,
  input  [7:0]  io_pipe_phv_in_data_109,
  input  [7:0]  io_pipe_phv_in_data_110,
  input  [7:0]  io_pipe_phv_in_data_111,
  input  [7:0]  io_pipe_phv_in_data_112,
  input  [7:0]  io_pipe_phv_in_data_113,
  input  [7:0]  io_pipe_phv_in_data_114,
  input  [7:0]  io_pipe_phv_in_data_115,
  input  [7:0]  io_pipe_phv_in_data_116,
  input  [7:0]  io_pipe_phv_in_data_117,
  input  [7:0]  io_pipe_phv_in_data_118,
  input  [7:0]  io_pipe_phv_in_data_119,
  input  [7:0]  io_pipe_phv_in_data_120,
  input  [7:0]  io_pipe_phv_in_data_121,
  input  [7:0]  io_pipe_phv_in_data_122,
  input  [7:0]  io_pipe_phv_in_data_123,
  input  [7:0]  io_pipe_phv_in_data_124,
  input  [7:0]  io_pipe_phv_in_data_125,
  input  [7:0]  io_pipe_phv_in_data_126,
  input  [7:0]  io_pipe_phv_in_data_127,
  input  [7:0]  io_pipe_phv_in_data_128,
  input  [7:0]  io_pipe_phv_in_data_129,
  input  [7:0]  io_pipe_phv_in_data_130,
  input  [7:0]  io_pipe_phv_in_data_131,
  input  [7:0]  io_pipe_phv_in_data_132,
  input  [7:0]  io_pipe_phv_in_data_133,
  input  [7:0]  io_pipe_phv_in_data_134,
  input  [7:0]  io_pipe_phv_in_data_135,
  input  [7:0]  io_pipe_phv_in_data_136,
  input  [7:0]  io_pipe_phv_in_data_137,
  input  [7:0]  io_pipe_phv_in_data_138,
  input  [7:0]  io_pipe_phv_in_data_139,
  input  [7:0]  io_pipe_phv_in_data_140,
  input  [7:0]  io_pipe_phv_in_data_141,
  input  [7:0]  io_pipe_phv_in_data_142,
  input  [7:0]  io_pipe_phv_in_data_143,
  input  [7:0]  io_pipe_phv_in_data_144,
  input  [7:0]  io_pipe_phv_in_data_145,
  input  [7:0]  io_pipe_phv_in_data_146,
  input  [7:0]  io_pipe_phv_in_data_147,
  input  [7:0]  io_pipe_phv_in_data_148,
  input  [7:0]  io_pipe_phv_in_data_149,
  input  [7:0]  io_pipe_phv_in_data_150,
  input  [7:0]  io_pipe_phv_in_data_151,
  input  [7:0]  io_pipe_phv_in_data_152,
  input  [7:0]  io_pipe_phv_in_data_153,
  input  [7:0]  io_pipe_phv_in_data_154,
  input  [7:0]  io_pipe_phv_in_data_155,
  input  [7:0]  io_pipe_phv_in_data_156,
  input  [7:0]  io_pipe_phv_in_data_157,
  input  [7:0]  io_pipe_phv_in_data_158,
  input  [7:0]  io_pipe_phv_in_data_159,
  input  [7:0]  io_pipe_phv_in_data_160,
  input  [7:0]  io_pipe_phv_in_data_161,
  input  [7:0]  io_pipe_phv_in_data_162,
  input  [7:0]  io_pipe_phv_in_data_163,
  input  [7:0]  io_pipe_phv_in_data_164,
  input  [7:0]  io_pipe_phv_in_data_165,
  input  [7:0]  io_pipe_phv_in_data_166,
  input  [7:0]  io_pipe_phv_in_data_167,
  input  [7:0]  io_pipe_phv_in_data_168,
  input  [7:0]  io_pipe_phv_in_data_169,
  input  [7:0]  io_pipe_phv_in_data_170,
  input  [7:0]  io_pipe_phv_in_data_171,
  input  [7:0]  io_pipe_phv_in_data_172,
  input  [7:0]  io_pipe_phv_in_data_173,
  input  [7:0]  io_pipe_phv_in_data_174,
  input  [7:0]  io_pipe_phv_in_data_175,
  input  [7:0]  io_pipe_phv_in_data_176,
  input  [7:0]  io_pipe_phv_in_data_177,
  input  [7:0]  io_pipe_phv_in_data_178,
  input  [7:0]  io_pipe_phv_in_data_179,
  input  [7:0]  io_pipe_phv_in_data_180,
  input  [7:0]  io_pipe_phv_in_data_181,
  input  [7:0]  io_pipe_phv_in_data_182,
  input  [7:0]  io_pipe_phv_in_data_183,
  input  [7:0]  io_pipe_phv_in_data_184,
  input  [7:0]  io_pipe_phv_in_data_185,
  input  [7:0]  io_pipe_phv_in_data_186,
  input  [7:0]  io_pipe_phv_in_data_187,
  input  [7:0]  io_pipe_phv_in_data_188,
  input  [7:0]  io_pipe_phv_in_data_189,
  input  [7:0]  io_pipe_phv_in_data_190,
  input  [7:0]  io_pipe_phv_in_data_191,
  input  [7:0]  io_pipe_phv_in_data_192,
  input  [7:0]  io_pipe_phv_in_data_193,
  input  [7:0]  io_pipe_phv_in_data_194,
  input  [7:0]  io_pipe_phv_in_data_195,
  input  [7:0]  io_pipe_phv_in_data_196,
  input  [7:0]  io_pipe_phv_in_data_197,
  input  [7:0]  io_pipe_phv_in_data_198,
  input  [7:0]  io_pipe_phv_in_data_199,
  input  [7:0]  io_pipe_phv_in_data_200,
  input  [7:0]  io_pipe_phv_in_data_201,
  input  [7:0]  io_pipe_phv_in_data_202,
  input  [7:0]  io_pipe_phv_in_data_203,
  input  [7:0]  io_pipe_phv_in_data_204,
  input  [7:0]  io_pipe_phv_in_data_205,
  input  [7:0]  io_pipe_phv_in_data_206,
  input  [7:0]  io_pipe_phv_in_data_207,
  input  [7:0]  io_pipe_phv_in_data_208,
  input  [7:0]  io_pipe_phv_in_data_209,
  input  [7:0]  io_pipe_phv_in_data_210,
  input  [7:0]  io_pipe_phv_in_data_211,
  input  [7:0]  io_pipe_phv_in_data_212,
  input  [7:0]  io_pipe_phv_in_data_213,
  input  [7:0]  io_pipe_phv_in_data_214,
  input  [7:0]  io_pipe_phv_in_data_215,
  input  [7:0]  io_pipe_phv_in_data_216,
  input  [7:0]  io_pipe_phv_in_data_217,
  input  [7:0]  io_pipe_phv_in_data_218,
  input  [7:0]  io_pipe_phv_in_data_219,
  input  [7:0]  io_pipe_phv_in_data_220,
  input  [7:0]  io_pipe_phv_in_data_221,
  input  [7:0]  io_pipe_phv_in_data_222,
  input  [7:0]  io_pipe_phv_in_data_223,
  input  [7:0]  io_pipe_phv_in_data_224,
  input  [7:0]  io_pipe_phv_in_data_225,
  input  [7:0]  io_pipe_phv_in_data_226,
  input  [7:0]  io_pipe_phv_in_data_227,
  input  [7:0]  io_pipe_phv_in_data_228,
  input  [7:0]  io_pipe_phv_in_data_229,
  input  [7:0]  io_pipe_phv_in_data_230,
  input  [7:0]  io_pipe_phv_in_data_231,
  input  [7:0]  io_pipe_phv_in_data_232,
  input  [7:0]  io_pipe_phv_in_data_233,
  input  [7:0]  io_pipe_phv_in_data_234,
  input  [7:0]  io_pipe_phv_in_data_235,
  input  [7:0]  io_pipe_phv_in_data_236,
  input  [7:0]  io_pipe_phv_in_data_237,
  input  [7:0]  io_pipe_phv_in_data_238,
  input  [7:0]  io_pipe_phv_in_data_239,
  input  [7:0]  io_pipe_phv_in_data_240,
  input  [7:0]  io_pipe_phv_in_data_241,
  input  [7:0]  io_pipe_phv_in_data_242,
  input  [7:0]  io_pipe_phv_in_data_243,
  input  [7:0]  io_pipe_phv_in_data_244,
  input  [7:0]  io_pipe_phv_in_data_245,
  input  [7:0]  io_pipe_phv_in_data_246,
  input  [7:0]  io_pipe_phv_in_data_247,
  input  [7:0]  io_pipe_phv_in_data_248,
  input  [7:0]  io_pipe_phv_in_data_249,
  input  [7:0]  io_pipe_phv_in_data_250,
  input  [7:0]  io_pipe_phv_in_data_251,
  input  [7:0]  io_pipe_phv_in_data_252,
  input  [7:0]  io_pipe_phv_in_data_253,
  input  [7:0]  io_pipe_phv_in_data_254,
  input  [7:0]  io_pipe_phv_in_data_255,
  input  [15:0] io_pipe_phv_in_header_0,
  input  [15:0] io_pipe_phv_in_header_1,
  input  [15:0] io_pipe_phv_in_header_2,
  input  [15:0] io_pipe_phv_in_header_3,
  input  [15:0] io_pipe_phv_in_header_4,
  input  [15:0] io_pipe_phv_in_header_5,
  input  [15:0] io_pipe_phv_in_header_6,
  input  [15:0] io_pipe_phv_in_header_7,
  input  [15:0] io_pipe_phv_in_header_8,
  input  [15:0] io_pipe_phv_in_header_9,
  input  [15:0] io_pipe_phv_in_header_10,
  input  [15:0] io_pipe_phv_in_header_11,
  input  [15:0] io_pipe_phv_in_header_12,
  input  [15:0] io_pipe_phv_in_header_13,
  input  [15:0] io_pipe_phv_in_header_14,
  input  [15:0] io_pipe_phv_in_header_15,
  input  [7:0]  io_pipe_phv_in_parse_current_state,
  input  [7:0]  io_pipe_phv_in_parse_current_offset,
  input  [15:0] io_pipe_phv_in_parse_transition_field,
  input  [2:0]  io_pipe_phv_in_next_processor_id,
  input         io_pipe_phv_in_next_config_id,
  input         io_pipe_phv_in_is_valid_processor,
  output [7:0]  io_pipe_phv_out_data_0,
  output [7:0]  io_pipe_phv_out_data_1,
  output [7:0]  io_pipe_phv_out_data_2,
  output [7:0]  io_pipe_phv_out_data_3,
  output [7:0]  io_pipe_phv_out_data_4,
  output [7:0]  io_pipe_phv_out_data_5,
  output [7:0]  io_pipe_phv_out_data_6,
  output [7:0]  io_pipe_phv_out_data_7,
  output [7:0]  io_pipe_phv_out_data_8,
  output [7:0]  io_pipe_phv_out_data_9,
  output [7:0]  io_pipe_phv_out_data_10,
  output [7:0]  io_pipe_phv_out_data_11,
  output [7:0]  io_pipe_phv_out_data_12,
  output [7:0]  io_pipe_phv_out_data_13,
  output [7:0]  io_pipe_phv_out_data_14,
  output [7:0]  io_pipe_phv_out_data_15,
  output [7:0]  io_pipe_phv_out_data_16,
  output [7:0]  io_pipe_phv_out_data_17,
  output [7:0]  io_pipe_phv_out_data_18,
  output [7:0]  io_pipe_phv_out_data_19,
  output [7:0]  io_pipe_phv_out_data_20,
  output [7:0]  io_pipe_phv_out_data_21,
  output [7:0]  io_pipe_phv_out_data_22,
  output [7:0]  io_pipe_phv_out_data_23,
  output [7:0]  io_pipe_phv_out_data_24,
  output [7:0]  io_pipe_phv_out_data_25,
  output [7:0]  io_pipe_phv_out_data_26,
  output [7:0]  io_pipe_phv_out_data_27,
  output [7:0]  io_pipe_phv_out_data_28,
  output [7:0]  io_pipe_phv_out_data_29,
  output [7:0]  io_pipe_phv_out_data_30,
  output [7:0]  io_pipe_phv_out_data_31,
  output [7:0]  io_pipe_phv_out_data_32,
  output [7:0]  io_pipe_phv_out_data_33,
  output [7:0]  io_pipe_phv_out_data_34,
  output [7:0]  io_pipe_phv_out_data_35,
  output [7:0]  io_pipe_phv_out_data_36,
  output [7:0]  io_pipe_phv_out_data_37,
  output [7:0]  io_pipe_phv_out_data_38,
  output [7:0]  io_pipe_phv_out_data_39,
  output [7:0]  io_pipe_phv_out_data_40,
  output [7:0]  io_pipe_phv_out_data_41,
  output [7:0]  io_pipe_phv_out_data_42,
  output [7:0]  io_pipe_phv_out_data_43,
  output [7:0]  io_pipe_phv_out_data_44,
  output [7:0]  io_pipe_phv_out_data_45,
  output [7:0]  io_pipe_phv_out_data_46,
  output [7:0]  io_pipe_phv_out_data_47,
  output [7:0]  io_pipe_phv_out_data_48,
  output [7:0]  io_pipe_phv_out_data_49,
  output [7:0]  io_pipe_phv_out_data_50,
  output [7:0]  io_pipe_phv_out_data_51,
  output [7:0]  io_pipe_phv_out_data_52,
  output [7:0]  io_pipe_phv_out_data_53,
  output [7:0]  io_pipe_phv_out_data_54,
  output [7:0]  io_pipe_phv_out_data_55,
  output [7:0]  io_pipe_phv_out_data_56,
  output [7:0]  io_pipe_phv_out_data_57,
  output [7:0]  io_pipe_phv_out_data_58,
  output [7:0]  io_pipe_phv_out_data_59,
  output [7:0]  io_pipe_phv_out_data_60,
  output [7:0]  io_pipe_phv_out_data_61,
  output [7:0]  io_pipe_phv_out_data_62,
  output [7:0]  io_pipe_phv_out_data_63,
  output [7:0]  io_pipe_phv_out_data_64,
  output [7:0]  io_pipe_phv_out_data_65,
  output [7:0]  io_pipe_phv_out_data_66,
  output [7:0]  io_pipe_phv_out_data_67,
  output [7:0]  io_pipe_phv_out_data_68,
  output [7:0]  io_pipe_phv_out_data_69,
  output [7:0]  io_pipe_phv_out_data_70,
  output [7:0]  io_pipe_phv_out_data_71,
  output [7:0]  io_pipe_phv_out_data_72,
  output [7:0]  io_pipe_phv_out_data_73,
  output [7:0]  io_pipe_phv_out_data_74,
  output [7:0]  io_pipe_phv_out_data_75,
  output [7:0]  io_pipe_phv_out_data_76,
  output [7:0]  io_pipe_phv_out_data_77,
  output [7:0]  io_pipe_phv_out_data_78,
  output [7:0]  io_pipe_phv_out_data_79,
  output [7:0]  io_pipe_phv_out_data_80,
  output [7:0]  io_pipe_phv_out_data_81,
  output [7:0]  io_pipe_phv_out_data_82,
  output [7:0]  io_pipe_phv_out_data_83,
  output [7:0]  io_pipe_phv_out_data_84,
  output [7:0]  io_pipe_phv_out_data_85,
  output [7:0]  io_pipe_phv_out_data_86,
  output [7:0]  io_pipe_phv_out_data_87,
  output [7:0]  io_pipe_phv_out_data_88,
  output [7:0]  io_pipe_phv_out_data_89,
  output [7:0]  io_pipe_phv_out_data_90,
  output [7:0]  io_pipe_phv_out_data_91,
  output [7:0]  io_pipe_phv_out_data_92,
  output [7:0]  io_pipe_phv_out_data_93,
  output [7:0]  io_pipe_phv_out_data_94,
  output [7:0]  io_pipe_phv_out_data_95,
  output [7:0]  io_pipe_phv_out_data_96,
  output [7:0]  io_pipe_phv_out_data_97,
  output [7:0]  io_pipe_phv_out_data_98,
  output [7:0]  io_pipe_phv_out_data_99,
  output [7:0]  io_pipe_phv_out_data_100,
  output [7:0]  io_pipe_phv_out_data_101,
  output [7:0]  io_pipe_phv_out_data_102,
  output [7:0]  io_pipe_phv_out_data_103,
  output [7:0]  io_pipe_phv_out_data_104,
  output [7:0]  io_pipe_phv_out_data_105,
  output [7:0]  io_pipe_phv_out_data_106,
  output [7:0]  io_pipe_phv_out_data_107,
  output [7:0]  io_pipe_phv_out_data_108,
  output [7:0]  io_pipe_phv_out_data_109,
  output [7:0]  io_pipe_phv_out_data_110,
  output [7:0]  io_pipe_phv_out_data_111,
  output [7:0]  io_pipe_phv_out_data_112,
  output [7:0]  io_pipe_phv_out_data_113,
  output [7:0]  io_pipe_phv_out_data_114,
  output [7:0]  io_pipe_phv_out_data_115,
  output [7:0]  io_pipe_phv_out_data_116,
  output [7:0]  io_pipe_phv_out_data_117,
  output [7:0]  io_pipe_phv_out_data_118,
  output [7:0]  io_pipe_phv_out_data_119,
  output [7:0]  io_pipe_phv_out_data_120,
  output [7:0]  io_pipe_phv_out_data_121,
  output [7:0]  io_pipe_phv_out_data_122,
  output [7:0]  io_pipe_phv_out_data_123,
  output [7:0]  io_pipe_phv_out_data_124,
  output [7:0]  io_pipe_phv_out_data_125,
  output [7:0]  io_pipe_phv_out_data_126,
  output [7:0]  io_pipe_phv_out_data_127,
  output [7:0]  io_pipe_phv_out_data_128,
  output [7:0]  io_pipe_phv_out_data_129,
  output [7:0]  io_pipe_phv_out_data_130,
  output [7:0]  io_pipe_phv_out_data_131,
  output [7:0]  io_pipe_phv_out_data_132,
  output [7:0]  io_pipe_phv_out_data_133,
  output [7:0]  io_pipe_phv_out_data_134,
  output [7:0]  io_pipe_phv_out_data_135,
  output [7:0]  io_pipe_phv_out_data_136,
  output [7:0]  io_pipe_phv_out_data_137,
  output [7:0]  io_pipe_phv_out_data_138,
  output [7:0]  io_pipe_phv_out_data_139,
  output [7:0]  io_pipe_phv_out_data_140,
  output [7:0]  io_pipe_phv_out_data_141,
  output [7:0]  io_pipe_phv_out_data_142,
  output [7:0]  io_pipe_phv_out_data_143,
  output [7:0]  io_pipe_phv_out_data_144,
  output [7:0]  io_pipe_phv_out_data_145,
  output [7:0]  io_pipe_phv_out_data_146,
  output [7:0]  io_pipe_phv_out_data_147,
  output [7:0]  io_pipe_phv_out_data_148,
  output [7:0]  io_pipe_phv_out_data_149,
  output [7:0]  io_pipe_phv_out_data_150,
  output [7:0]  io_pipe_phv_out_data_151,
  output [7:0]  io_pipe_phv_out_data_152,
  output [7:0]  io_pipe_phv_out_data_153,
  output [7:0]  io_pipe_phv_out_data_154,
  output [7:0]  io_pipe_phv_out_data_155,
  output [7:0]  io_pipe_phv_out_data_156,
  output [7:0]  io_pipe_phv_out_data_157,
  output [7:0]  io_pipe_phv_out_data_158,
  output [7:0]  io_pipe_phv_out_data_159,
  output [7:0]  io_pipe_phv_out_data_160,
  output [7:0]  io_pipe_phv_out_data_161,
  output [7:0]  io_pipe_phv_out_data_162,
  output [7:0]  io_pipe_phv_out_data_163,
  output [7:0]  io_pipe_phv_out_data_164,
  output [7:0]  io_pipe_phv_out_data_165,
  output [7:0]  io_pipe_phv_out_data_166,
  output [7:0]  io_pipe_phv_out_data_167,
  output [7:0]  io_pipe_phv_out_data_168,
  output [7:0]  io_pipe_phv_out_data_169,
  output [7:0]  io_pipe_phv_out_data_170,
  output [7:0]  io_pipe_phv_out_data_171,
  output [7:0]  io_pipe_phv_out_data_172,
  output [7:0]  io_pipe_phv_out_data_173,
  output [7:0]  io_pipe_phv_out_data_174,
  output [7:0]  io_pipe_phv_out_data_175,
  output [7:0]  io_pipe_phv_out_data_176,
  output [7:0]  io_pipe_phv_out_data_177,
  output [7:0]  io_pipe_phv_out_data_178,
  output [7:0]  io_pipe_phv_out_data_179,
  output [7:0]  io_pipe_phv_out_data_180,
  output [7:0]  io_pipe_phv_out_data_181,
  output [7:0]  io_pipe_phv_out_data_182,
  output [7:0]  io_pipe_phv_out_data_183,
  output [7:0]  io_pipe_phv_out_data_184,
  output [7:0]  io_pipe_phv_out_data_185,
  output [7:0]  io_pipe_phv_out_data_186,
  output [7:0]  io_pipe_phv_out_data_187,
  output [7:0]  io_pipe_phv_out_data_188,
  output [7:0]  io_pipe_phv_out_data_189,
  output [7:0]  io_pipe_phv_out_data_190,
  output [7:0]  io_pipe_phv_out_data_191,
  output [7:0]  io_pipe_phv_out_data_192,
  output [7:0]  io_pipe_phv_out_data_193,
  output [7:0]  io_pipe_phv_out_data_194,
  output [7:0]  io_pipe_phv_out_data_195,
  output [7:0]  io_pipe_phv_out_data_196,
  output [7:0]  io_pipe_phv_out_data_197,
  output [7:0]  io_pipe_phv_out_data_198,
  output [7:0]  io_pipe_phv_out_data_199,
  output [7:0]  io_pipe_phv_out_data_200,
  output [7:0]  io_pipe_phv_out_data_201,
  output [7:0]  io_pipe_phv_out_data_202,
  output [7:0]  io_pipe_phv_out_data_203,
  output [7:0]  io_pipe_phv_out_data_204,
  output [7:0]  io_pipe_phv_out_data_205,
  output [7:0]  io_pipe_phv_out_data_206,
  output [7:0]  io_pipe_phv_out_data_207,
  output [7:0]  io_pipe_phv_out_data_208,
  output [7:0]  io_pipe_phv_out_data_209,
  output [7:0]  io_pipe_phv_out_data_210,
  output [7:0]  io_pipe_phv_out_data_211,
  output [7:0]  io_pipe_phv_out_data_212,
  output [7:0]  io_pipe_phv_out_data_213,
  output [7:0]  io_pipe_phv_out_data_214,
  output [7:0]  io_pipe_phv_out_data_215,
  output [7:0]  io_pipe_phv_out_data_216,
  output [7:0]  io_pipe_phv_out_data_217,
  output [7:0]  io_pipe_phv_out_data_218,
  output [7:0]  io_pipe_phv_out_data_219,
  output [7:0]  io_pipe_phv_out_data_220,
  output [7:0]  io_pipe_phv_out_data_221,
  output [7:0]  io_pipe_phv_out_data_222,
  output [7:0]  io_pipe_phv_out_data_223,
  output [7:0]  io_pipe_phv_out_data_224,
  output [7:0]  io_pipe_phv_out_data_225,
  output [7:0]  io_pipe_phv_out_data_226,
  output [7:0]  io_pipe_phv_out_data_227,
  output [7:0]  io_pipe_phv_out_data_228,
  output [7:0]  io_pipe_phv_out_data_229,
  output [7:0]  io_pipe_phv_out_data_230,
  output [7:0]  io_pipe_phv_out_data_231,
  output [7:0]  io_pipe_phv_out_data_232,
  output [7:0]  io_pipe_phv_out_data_233,
  output [7:0]  io_pipe_phv_out_data_234,
  output [7:0]  io_pipe_phv_out_data_235,
  output [7:0]  io_pipe_phv_out_data_236,
  output [7:0]  io_pipe_phv_out_data_237,
  output [7:0]  io_pipe_phv_out_data_238,
  output [7:0]  io_pipe_phv_out_data_239,
  output [7:0]  io_pipe_phv_out_data_240,
  output [7:0]  io_pipe_phv_out_data_241,
  output [7:0]  io_pipe_phv_out_data_242,
  output [7:0]  io_pipe_phv_out_data_243,
  output [7:0]  io_pipe_phv_out_data_244,
  output [7:0]  io_pipe_phv_out_data_245,
  output [7:0]  io_pipe_phv_out_data_246,
  output [7:0]  io_pipe_phv_out_data_247,
  output [7:0]  io_pipe_phv_out_data_248,
  output [7:0]  io_pipe_phv_out_data_249,
  output [7:0]  io_pipe_phv_out_data_250,
  output [7:0]  io_pipe_phv_out_data_251,
  output [7:0]  io_pipe_phv_out_data_252,
  output [7:0]  io_pipe_phv_out_data_253,
  output [7:0]  io_pipe_phv_out_data_254,
  output [7:0]  io_pipe_phv_out_data_255,
  output [15:0] io_pipe_phv_out_header_0,
  output [15:0] io_pipe_phv_out_header_1,
  output [15:0] io_pipe_phv_out_header_2,
  output [15:0] io_pipe_phv_out_header_3,
  output [15:0] io_pipe_phv_out_header_4,
  output [15:0] io_pipe_phv_out_header_5,
  output [15:0] io_pipe_phv_out_header_6,
  output [15:0] io_pipe_phv_out_header_7,
  output [15:0] io_pipe_phv_out_header_8,
  output [15:0] io_pipe_phv_out_header_9,
  output [15:0] io_pipe_phv_out_header_10,
  output [15:0] io_pipe_phv_out_header_11,
  output [15:0] io_pipe_phv_out_header_12,
  output [15:0] io_pipe_phv_out_header_13,
  output [15:0] io_pipe_phv_out_header_14,
  output [15:0] io_pipe_phv_out_header_15,
  output [7:0]  io_pipe_phv_out_parse_current_state,
  output [7:0]  io_pipe_phv_out_parse_current_offset,
  output [15:0] io_pipe_phv_out_parse_transition_field,
  output [2:0]  io_pipe_phv_out_next_processor_id,
  output        io_pipe_phv_out_next_config_id,
  output        io_pipe_phv_out_is_valid_processor,
  input         io_mod_en,
  input         io_mod_last_mau_id_mod,
  input  [1:0]  io_mod_last_mau_id,
  input  [1:0]  io_mod_cs,
  input         io_mod_module_mod_state_id_mod,
  input  [7:0]  io_mod_module_mod_state_id,
  input         io_mod_module_mod_sram_w_cs,
  input         io_mod_module_mod_sram_w_en,
  input  [7:0]  io_mod_module_mod_sram_w_addr,
  input  [63:0] io_mod_module_mod_sram_w_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  mau_0_clock; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_0; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_1; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_2; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_3; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_4; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_5; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_6; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_7; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_8; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_9; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_10; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_11; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_12; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_13; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_14; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_15; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_16; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_17; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_18; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_19; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_20; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_21; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_22; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_23; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_24; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_25; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_26; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_27; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_28; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_29; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_30; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_31; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_32; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_33; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_34; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_35; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_36; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_37; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_38; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_39; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_40; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_41; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_42; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_43; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_44; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_45; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_46; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_47; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_48; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_49; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_50; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_51; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_52; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_53; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_54; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_55; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_56; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_57; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_58; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_59; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_60; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_61; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_62; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_63; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_64; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_65; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_66; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_67; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_68; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_69; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_70; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_71; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_72; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_73; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_74; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_75; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_76; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_77; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_78; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_79; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_80; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_81; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_82; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_83; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_84; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_85; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_86; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_87; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_88; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_89; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_90; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_91; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_92; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_93; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_94; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_95; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_96; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_97; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_98; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_99; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_100; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_101; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_102; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_103; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_104; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_105; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_106; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_107; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_108; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_109; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_110; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_111; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_112; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_113; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_114; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_115; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_116; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_117; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_118; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_119; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_120; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_121; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_122; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_123; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_124; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_125; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_126; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_127; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_128; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_129; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_130; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_131; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_132; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_133; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_134; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_135; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_136; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_137; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_138; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_139; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_140; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_141; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_142; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_143; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_144; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_145; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_146; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_147; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_148; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_149; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_150; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_151; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_152; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_153; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_154; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_155; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_156; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_157; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_158; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_159; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_160; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_161; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_162; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_163; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_164; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_165; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_166; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_167; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_168; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_169; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_170; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_171; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_172; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_173; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_174; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_175; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_176; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_177; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_178; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_179; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_180; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_181; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_182; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_183; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_184; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_185; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_186; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_187; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_188; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_189; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_190; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_191; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_192; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_193; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_194; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_195; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_196; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_197; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_198; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_199; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_200; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_201; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_202; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_203; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_204; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_205; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_206; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_207; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_208; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_209; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_210; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_211; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_212; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_213; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_214; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_215; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_216; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_217; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_218; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_219; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_220; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_221; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_222; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_223; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_224; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_225; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_226; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_227; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_228; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_229; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_230; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_231; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_232; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_233; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_234; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_235; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_236; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_237; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_238; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_239; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_240; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_241; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_242; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_243; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_244; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_245; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_246; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_247; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_248; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_249; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_250; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_251; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_252; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_253; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_254; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_255; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_0; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_1; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_2; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_3; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_4; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_5; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_6; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_7; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_8; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_9; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_10; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_11; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_12; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_13; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_14; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_15; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_parse_current_state; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_parse_current_offset; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_in_parse_transition_field; // @[parser.scala 21:25]
  wire [2:0] mau_0_io_pipe_phv_in_next_processor_id; // @[parser.scala 21:25]
  wire  mau_0_io_pipe_phv_in_next_config_id; // @[parser.scala 21:25]
  wire  mau_0_io_pipe_phv_in_is_valid_processor; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_0; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_1; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_2; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_3; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_4; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_5; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_6; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_7; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_8; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_9; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_10; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_11; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_12; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_13; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_14; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_15; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_16; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_17; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_18; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_19; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_20; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_21; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_22; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_23; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_24; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_25; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_26; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_27; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_28; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_29; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_30; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_31; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_32; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_33; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_34; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_35; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_36; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_37; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_38; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_39; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_40; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_41; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_42; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_43; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_44; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_45; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_46; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_47; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_48; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_49; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_50; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_51; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_52; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_53; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_54; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_55; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_56; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_57; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_58; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_59; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_60; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_61; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_62; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_63; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_64; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_65; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_66; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_67; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_68; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_69; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_70; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_71; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_72; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_73; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_74; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_75; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_76; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_77; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_78; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_79; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_80; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_81; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_82; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_83; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_84; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_85; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_86; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_87; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_88; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_89; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_90; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_91; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_92; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_93; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_94; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_95; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_96; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_97; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_98; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_99; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_100; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_101; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_102; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_103; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_104; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_105; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_106; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_107; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_108; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_109; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_110; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_111; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_112; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_113; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_114; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_115; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_116; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_117; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_118; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_119; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_120; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_121; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_122; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_123; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_124; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_125; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_126; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_127; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_128; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_129; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_130; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_131; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_132; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_133; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_134; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_135; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_136; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_137; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_138; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_139; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_140; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_141; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_142; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_143; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_144; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_145; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_146; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_147; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_148; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_149; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_150; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_151; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_152; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_153; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_154; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_155; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_156; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_157; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_158; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_159; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_160; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_161; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_162; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_163; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_164; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_165; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_166; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_167; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_168; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_169; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_170; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_171; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_172; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_173; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_174; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_175; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_176; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_177; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_178; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_179; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_180; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_181; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_182; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_183; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_184; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_185; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_186; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_187; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_188; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_189; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_190; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_191; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_192; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_193; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_194; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_195; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_196; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_197; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_198; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_199; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_200; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_201; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_202; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_203; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_204; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_205; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_206; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_207; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_208; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_209; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_210; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_211; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_212; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_213; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_214; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_215; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_216; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_217; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_218; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_219; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_220; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_221; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_222; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_223; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_224; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_225; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_226; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_227; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_228; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_229; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_230; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_231; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_232; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_233; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_234; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_235; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_236; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_237; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_238; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_239; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_240; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_241; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_242; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_243; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_244; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_245; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_246; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_247; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_248; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_249; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_250; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_251; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_252; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_253; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_254; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_255; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_0; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_1; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_2; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_3; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_4; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_5; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_6; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_7; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_8; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_9; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_10; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_11; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_12; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_13; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_14; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_15; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_parse_current_state; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_parse_current_offset; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_out_parse_transition_field; // @[parser.scala 21:25]
  wire [2:0] mau_0_io_pipe_phv_out_next_processor_id; // @[parser.scala 21:25]
  wire  mau_0_io_pipe_phv_out_next_config_id; // @[parser.scala 21:25]
  wire  mau_0_io_pipe_phv_out_is_valid_processor; // @[parser.scala 21:25]
  wire  mau_0_io_mod_state_id_mod; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_mod_state_id; // @[parser.scala 21:25]
  wire  mau_0_io_mod_sram_w_cs; // @[parser.scala 21:25]
  wire  mau_0_io_mod_sram_w_en; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_mod_sram_w_addr; // @[parser.scala 21:25]
  wire [63:0] mau_0_io_mod_sram_w_data; // @[parser.scala 21:25]
  wire  mau_1_clock; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_0; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_1; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_2; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_3; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_4; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_5; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_6; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_7; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_8; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_9; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_10; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_11; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_12; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_13; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_14; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_15; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_16; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_17; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_18; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_19; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_20; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_21; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_22; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_23; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_24; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_25; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_26; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_27; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_28; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_29; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_30; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_31; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_32; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_33; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_34; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_35; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_36; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_37; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_38; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_39; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_40; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_41; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_42; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_43; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_44; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_45; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_46; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_47; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_48; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_49; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_50; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_51; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_52; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_53; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_54; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_55; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_56; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_57; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_58; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_59; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_60; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_61; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_62; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_63; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_64; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_65; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_66; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_67; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_68; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_69; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_70; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_71; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_72; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_73; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_74; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_75; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_76; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_77; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_78; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_79; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_80; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_81; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_82; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_83; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_84; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_85; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_86; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_87; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_88; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_89; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_90; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_91; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_92; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_93; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_94; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_95; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_96; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_97; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_98; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_99; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_100; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_101; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_102; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_103; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_104; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_105; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_106; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_107; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_108; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_109; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_110; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_111; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_112; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_113; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_114; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_115; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_116; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_117; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_118; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_119; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_120; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_121; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_122; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_123; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_124; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_125; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_126; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_127; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_128; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_129; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_130; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_131; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_132; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_133; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_134; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_135; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_136; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_137; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_138; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_139; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_140; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_141; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_142; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_143; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_144; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_145; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_146; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_147; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_148; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_149; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_150; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_151; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_152; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_153; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_154; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_155; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_156; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_157; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_158; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_159; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_160; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_161; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_162; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_163; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_164; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_165; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_166; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_167; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_168; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_169; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_170; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_171; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_172; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_173; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_174; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_175; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_176; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_177; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_178; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_179; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_180; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_181; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_182; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_183; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_184; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_185; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_186; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_187; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_188; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_189; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_190; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_191; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_192; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_193; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_194; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_195; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_196; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_197; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_198; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_199; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_200; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_201; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_202; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_203; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_204; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_205; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_206; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_207; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_208; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_209; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_210; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_211; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_212; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_213; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_214; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_215; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_216; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_217; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_218; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_219; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_220; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_221; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_222; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_223; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_224; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_225; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_226; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_227; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_228; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_229; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_230; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_231; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_232; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_233; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_234; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_235; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_236; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_237; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_238; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_239; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_240; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_241; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_242; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_243; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_244; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_245; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_246; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_247; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_248; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_249; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_250; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_251; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_252; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_253; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_254; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_255; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_0; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_1; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_2; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_3; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_4; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_5; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_6; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_7; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_8; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_9; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_10; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_11; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_12; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_13; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_14; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_15; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_parse_current_state; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_parse_current_offset; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_in_parse_transition_field; // @[parser.scala 21:25]
  wire [2:0] mau_1_io_pipe_phv_in_next_processor_id; // @[parser.scala 21:25]
  wire  mau_1_io_pipe_phv_in_next_config_id; // @[parser.scala 21:25]
  wire  mau_1_io_pipe_phv_in_is_valid_processor; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_0; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_1; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_2; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_3; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_4; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_5; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_6; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_7; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_8; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_9; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_10; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_11; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_12; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_13; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_14; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_15; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_16; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_17; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_18; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_19; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_20; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_21; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_22; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_23; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_24; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_25; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_26; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_27; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_28; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_29; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_30; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_31; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_32; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_33; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_34; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_35; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_36; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_37; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_38; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_39; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_40; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_41; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_42; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_43; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_44; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_45; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_46; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_47; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_48; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_49; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_50; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_51; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_52; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_53; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_54; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_55; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_56; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_57; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_58; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_59; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_60; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_61; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_62; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_63; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_64; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_65; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_66; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_67; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_68; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_69; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_70; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_71; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_72; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_73; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_74; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_75; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_76; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_77; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_78; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_79; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_80; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_81; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_82; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_83; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_84; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_85; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_86; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_87; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_88; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_89; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_90; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_91; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_92; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_93; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_94; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_95; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_96; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_97; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_98; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_99; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_100; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_101; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_102; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_103; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_104; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_105; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_106; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_107; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_108; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_109; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_110; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_111; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_112; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_113; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_114; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_115; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_116; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_117; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_118; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_119; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_120; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_121; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_122; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_123; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_124; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_125; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_126; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_127; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_128; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_129; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_130; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_131; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_132; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_133; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_134; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_135; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_136; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_137; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_138; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_139; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_140; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_141; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_142; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_143; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_144; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_145; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_146; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_147; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_148; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_149; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_150; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_151; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_152; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_153; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_154; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_155; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_156; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_157; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_158; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_159; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_160; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_161; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_162; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_163; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_164; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_165; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_166; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_167; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_168; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_169; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_170; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_171; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_172; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_173; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_174; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_175; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_176; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_177; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_178; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_179; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_180; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_181; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_182; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_183; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_184; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_185; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_186; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_187; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_188; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_189; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_190; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_191; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_192; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_193; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_194; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_195; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_196; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_197; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_198; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_199; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_200; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_201; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_202; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_203; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_204; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_205; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_206; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_207; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_208; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_209; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_210; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_211; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_212; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_213; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_214; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_215; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_216; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_217; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_218; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_219; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_220; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_221; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_222; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_223; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_224; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_225; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_226; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_227; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_228; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_229; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_230; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_231; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_232; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_233; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_234; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_235; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_236; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_237; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_238; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_239; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_240; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_241; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_242; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_243; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_244; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_245; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_246; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_247; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_248; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_249; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_250; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_251; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_252; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_253; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_254; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_255; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_0; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_1; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_2; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_3; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_4; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_5; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_6; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_7; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_8; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_9; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_10; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_11; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_12; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_13; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_14; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_15; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_parse_current_state; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_parse_current_offset; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_out_parse_transition_field; // @[parser.scala 21:25]
  wire [2:0] mau_1_io_pipe_phv_out_next_processor_id; // @[parser.scala 21:25]
  wire  mau_1_io_pipe_phv_out_next_config_id; // @[parser.scala 21:25]
  wire  mau_1_io_pipe_phv_out_is_valid_processor; // @[parser.scala 21:25]
  wire  mau_1_io_mod_state_id_mod; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_mod_state_id; // @[parser.scala 21:25]
  wire  mau_1_io_mod_sram_w_cs; // @[parser.scala 21:25]
  wire  mau_1_io_mod_sram_w_en; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_mod_sram_w_addr; // @[parser.scala 21:25]
  wire [63:0] mau_1_io_mod_sram_w_data; // @[parser.scala 21:25]
  wire  mau_2_clock; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_0; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_1; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_2; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_3; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_4; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_5; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_6; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_7; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_8; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_9; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_10; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_11; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_12; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_13; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_14; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_15; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_16; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_17; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_18; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_19; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_20; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_21; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_22; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_23; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_24; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_25; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_26; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_27; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_28; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_29; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_30; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_31; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_32; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_33; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_34; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_35; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_36; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_37; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_38; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_39; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_40; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_41; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_42; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_43; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_44; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_45; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_46; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_47; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_48; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_49; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_50; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_51; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_52; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_53; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_54; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_55; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_56; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_57; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_58; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_59; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_60; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_61; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_62; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_63; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_64; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_65; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_66; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_67; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_68; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_69; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_70; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_71; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_72; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_73; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_74; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_75; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_76; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_77; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_78; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_79; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_80; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_81; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_82; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_83; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_84; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_85; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_86; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_87; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_88; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_89; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_90; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_91; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_92; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_93; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_94; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_95; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_96; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_97; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_98; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_99; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_100; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_101; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_102; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_103; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_104; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_105; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_106; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_107; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_108; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_109; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_110; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_111; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_112; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_113; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_114; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_115; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_116; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_117; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_118; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_119; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_120; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_121; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_122; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_123; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_124; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_125; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_126; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_127; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_128; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_129; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_130; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_131; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_132; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_133; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_134; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_135; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_136; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_137; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_138; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_139; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_140; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_141; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_142; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_143; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_144; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_145; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_146; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_147; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_148; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_149; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_150; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_151; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_152; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_153; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_154; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_155; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_156; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_157; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_158; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_159; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_160; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_161; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_162; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_163; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_164; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_165; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_166; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_167; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_168; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_169; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_170; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_171; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_172; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_173; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_174; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_175; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_176; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_177; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_178; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_179; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_180; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_181; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_182; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_183; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_184; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_185; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_186; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_187; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_188; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_189; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_190; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_191; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_192; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_193; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_194; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_195; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_196; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_197; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_198; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_199; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_200; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_201; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_202; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_203; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_204; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_205; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_206; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_207; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_208; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_209; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_210; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_211; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_212; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_213; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_214; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_215; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_216; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_217; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_218; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_219; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_220; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_221; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_222; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_223; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_224; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_225; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_226; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_227; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_228; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_229; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_230; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_231; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_232; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_233; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_234; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_235; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_236; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_237; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_238; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_239; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_240; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_241; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_242; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_243; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_244; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_245; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_246; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_247; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_248; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_249; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_250; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_251; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_252; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_253; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_254; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_255; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_0; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_1; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_2; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_3; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_4; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_5; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_6; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_7; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_8; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_9; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_10; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_11; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_12; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_13; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_14; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_15; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_parse_current_state; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_parse_current_offset; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_in_parse_transition_field; // @[parser.scala 21:25]
  wire [2:0] mau_2_io_pipe_phv_in_next_processor_id; // @[parser.scala 21:25]
  wire  mau_2_io_pipe_phv_in_next_config_id; // @[parser.scala 21:25]
  wire  mau_2_io_pipe_phv_in_is_valid_processor; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_0; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_1; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_2; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_3; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_4; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_5; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_6; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_7; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_8; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_9; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_10; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_11; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_12; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_13; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_14; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_15; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_16; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_17; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_18; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_19; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_20; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_21; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_22; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_23; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_24; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_25; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_26; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_27; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_28; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_29; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_30; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_31; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_32; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_33; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_34; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_35; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_36; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_37; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_38; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_39; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_40; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_41; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_42; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_43; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_44; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_45; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_46; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_47; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_48; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_49; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_50; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_51; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_52; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_53; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_54; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_55; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_56; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_57; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_58; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_59; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_60; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_61; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_62; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_63; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_64; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_65; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_66; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_67; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_68; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_69; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_70; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_71; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_72; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_73; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_74; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_75; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_76; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_77; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_78; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_79; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_80; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_81; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_82; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_83; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_84; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_85; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_86; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_87; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_88; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_89; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_90; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_91; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_92; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_93; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_94; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_95; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_96; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_97; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_98; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_99; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_100; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_101; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_102; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_103; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_104; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_105; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_106; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_107; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_108; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_109; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_110; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_111; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_112; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_113; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_114; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_115; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_116; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_117; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_118; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_119; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_120; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_121; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_122; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_123; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_124; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_125; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_126; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_127; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_128; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_129; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_130; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_131; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_132; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_133; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_134; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_135; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_136; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_137; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_138; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_139; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_140; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_141; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_142; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_143; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_144; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_145; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_146; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_147; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_148; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_149; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_150; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_151; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_152; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_153; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_154; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_155; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_156; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_157; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_158; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_159; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_160; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_161; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_162; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_163; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_164; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_165; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_166; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_167; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_168; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_169; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_170; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_171; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_172; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_173; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_174; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_175; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_176; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_177; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_178; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_179; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_180; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_181; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_182; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_183; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_184; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_185; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_186; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_187; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_188; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_189; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_190; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_191; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_192; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_193; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_194; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_195; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_196; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_197; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_198; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_199; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_200; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_201; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_202; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_203; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_204; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_205; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_206; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_207; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_208; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_209; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_210; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_211; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_212; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_213; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_214; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_215; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_216; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_217; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_218; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_219; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_220; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_221; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_222; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_223; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_224; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_225; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_226; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_227; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_228; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_229; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_230; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_231; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_232; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_233; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_234; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_235; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_236; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_237; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_238; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_239; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_240; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_241; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_242; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_243; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_244; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_245; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_246; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_247; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_248; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_249; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_250; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_251; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_252; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_253; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_254; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_255; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_0; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_1; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_2; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_3; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_4; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_5; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_6; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_7; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_8; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_9; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_10; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_11; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_12; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_13; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_14; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_15; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_parse_current_state; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_parse_current_offset; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_out_parse_transition_field; // @[parser.scala 21:25]
  wire [2:0] mau_2_io_pipe_phv_out_next_processor_id; // @[parser.scala 21:25]
  wire  mau_2_io_pipe_phv_out_next_config_id; // @[parser.scala 21:25]
  wire  mau_2_io_pipe_phv_out_is_valid_processor; // @[parser.scala 21:25]
  wire  mau_2_io_mod_state_id_mod; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_mod_state_id; // @[parser.scala 21:25]
  wire  mau_2_io_mod_sram_w_cs; // @[parser.scala 21:25]
  wire  mau_2_io_mod_sram_w_en; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_mod_sram_w_addr; // @[parser.scala 21:25]
  wire [63:0] mau_2_io_mod_sram_w_data; // @[parser.scala 21:25]
  wire  mau_3_clock; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_0; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_1; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_2; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_3; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_4; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_5; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_6; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_7; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_8; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_9; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_10; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_11; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_12; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_13; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_14; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_15; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_16; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_17; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_18; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_19; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_20; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_21; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_22; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_23; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_24; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_25; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_26; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_27; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_28; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_29; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_30; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_31; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_32; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_33; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_34; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_35; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_36; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_37; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_38; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_39; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_40; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_41; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_42; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_43; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_44; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_45; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_46; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_47; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_48; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_49; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_50; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_51; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_52; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_53; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_54; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_55; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_56; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_57; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_58; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_59; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_60; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_61; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_62; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_63; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_64; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_65; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_66; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_67; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_68; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_69; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_70; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_71; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_72; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_73; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_74; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_75; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_76; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_77; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_78; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_79; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_80; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_81; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_82; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_83; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_84; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_85; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_86; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_87; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_88; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_89; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_90; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_91; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_92; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_93; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_94; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_95; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_96; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_97; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_98; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_99; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_100; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_101; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_102; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_103; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_104; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_105; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_106; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_107; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_108; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_109; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_110; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_111; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_112; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_113; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_114; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_115; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_116; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_117; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_118; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_119; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_120; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_121; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_122; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_123; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_124; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_125; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_126; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_127; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_128; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_129; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_130; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_131; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_132; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_133; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_134; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_135; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_136; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_137; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_138; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_139; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_140; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_141; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_142; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_143; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_144; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_145; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_146; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_147; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_148; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_149; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_150; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_151; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_152; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_153; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_154; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_155; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_156; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_157; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_158; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_159; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_160; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_161; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_162; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_163; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_164; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_165; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_166; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_167; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_168; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_169; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_170; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_171; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_172; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_173; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_174; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_175; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_176; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_177; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_178; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_179; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_180; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_181; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_182; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_183; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_184; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_185; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_186; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_187; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_188; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_189; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_190; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_191; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_192; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_193; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_194; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_195; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_196; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_197; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_198; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_199; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_200; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_201; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_202; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_203; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_204; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_205; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_206; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_207; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_208; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_209; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_210; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_211; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_212; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_213; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_214; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_215; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_216; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_217; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_218; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_219; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_220; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_221; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_222; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_223; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_224; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_225; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_226; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_227; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_228; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_229; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_230; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_231; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_232; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_233; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_234; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_235; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_236; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_237; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_238; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_239; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_240; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_241; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_242; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_243; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_244; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_245; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_246; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_247; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_248; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_249; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_250; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_251; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_252; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_253; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_254; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_255; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_0; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_1; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_2; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_3; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_4; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_5; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_6; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_7; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_8; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_9; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_10; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_11; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_12; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_13; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_14; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_15; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_parse_current_state; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_parse_current_offset; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_in_parse_transition_field; // @[parser.scala 21:25]
  wire [2:0] mau_3_io_pipe_phv_in_next_processor_id; // @[parser.scala 21:25]
  wire  mau_3_io_pipe_phv_in_next_config_id; // @[parser.scala 21:25]
  wire  mau_3_io_pipe_phv_in_is_valid_processor; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_0; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_1; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_2; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_3; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_4; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_5; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_6; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_7; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_8; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_9; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_10; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_11; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_12; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_13; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_14; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_15; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_16; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_17; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_18; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_19; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_20; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_21; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_22; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_23; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_24; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_25; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_26; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_27; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_28; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_29; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_30; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_31; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_32; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_33; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_34; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_35; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_36; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_37; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_38; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_39; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_40; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_41; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_42; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_43; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_44; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_45; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_46; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_47; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_48; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_49; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_50; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_51; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_52; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_53; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_54; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_55; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_56; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_57; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_58; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_59; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_60; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_61; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_62; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_63; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_64; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_65; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_66; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_67; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_68; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_69; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_70; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_71; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_72; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_73; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_74; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_75; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_76; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_77; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_78; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_79; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_80; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_81; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_82; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_83; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_84; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_85; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_86; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_87; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_88; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_89; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_90; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_91; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_92; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_93; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_94; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_95; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_96; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_97; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_98; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_99; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_100; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_101; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_102; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_103; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_104; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_105; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_106; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_107; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_108; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_109; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_110; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_111; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_112; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_113; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_114; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_115; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_116; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_117; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_118; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_119; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_120; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_121; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_122; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_123; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_124; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_125; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_126; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_127; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_128; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_129; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_130; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_131; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_132; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_133; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_134; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_135; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_136; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_137; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_138; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_139; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_140; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_141; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_142; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_143; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_144; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_145; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_146; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_147; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_148; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_149; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_150; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_151; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_152; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_153; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_154; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_155; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_156; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_157; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_158; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_159; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_160; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_161; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_162; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_163; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_164; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_165; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_166; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_167; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_168; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_169; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_170; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_171; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_172; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_173; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_174; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_175; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_176; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_177; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_178; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_179; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_180; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_181; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_182; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_183; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_184; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_185; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_186; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_187; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_188; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_189; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_190; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_191; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_192; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_193; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_194; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_195; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_196; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_197; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_198; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_199; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_200; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_201; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_202; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_203; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_204; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_205; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_206; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_207; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_208; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_209; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_210; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_211; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_212; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_213; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_214; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_215; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_216; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_217; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_218; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_219; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_220; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_221; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_222; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_223; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_224; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_225; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_226; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_227; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_228; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_229; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_230; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_231; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_232; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_233; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_234; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_235; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_236; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_237; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_238; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_239; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_240; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_241; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_242; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_243; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_244; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_245; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_246; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_247; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_248; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_249; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_250; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_251; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_252; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_253; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_254; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_255; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_0; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_1; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_2; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_3; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_4; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_5; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_6; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_7; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_8; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_9; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_10; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_11; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_12; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_13; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_14; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_15; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_parse_current_state; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_parse_current_offset; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_out_parse_transition_field; // @[parser.scala 21:25]
  wire [2:0] mau_3_io_pipe_phv_out_next_processor_id; // @[parser.scala 21:25]
  wire  mau_3_io_pipe_phv_out_next_config_id; // @[parser.scala 21:25]
  wire  mau_3_io_pipe_phv_out_is_valid_processor; // @[parser.scala 21:25]
  wire  mau_3_io_mod_state_id_mod; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_mod_state_id; // @[parser.scala 21:25]
  wire  mau_3_io_mod_sram_w_cs; // @[parser.scala 21:25]
  wire  mau_3_io_mod_sram_w_en; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_mod_sram_w_addr; // @[parser.scala 21:25]
  wire [63:0] mau_3_io_mod_sram_w_data; // @[parser.scala 21:25]
  reg [2:0] last_mau_id; // @[parser.scala 14:26]
  wire  _GEN_0 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_is_valid_processor : io_pipe_phv_in_is_valid_processor; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire  _GEN_1 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_next_config_id : io_pipe_phv_in_next_config_id; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [2:0] _GEN_2 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_next_processor_id : io_pipe_phv_in_next_processor_id; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [15:0] _GEN_3 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_parse_transition_field :
    io_pipe_phv_in_parse_transition_field; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_4 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_parse_current_offset :
    io_pipe_phv_in_parse_current_offset; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_5 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_parse_current_state :
    io_pipe_phv_in_parse_current_state; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [15:0] _GEN_6 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_header_0 : io_pipe_phv_in_header_0; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [15:0] _GEN_7 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_header_1 : io_pipe_phv_in_header_1; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [15:0] _GEN_8 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_header_2 : io_pipe_phv_in_header_2; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [15:0] _GEN_9 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_header_3 : io_pipe_phv_in_header_3; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [15:0] _GEN_10 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_header_4 : io_pipe_phv_in_header_4; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [15:0] _GEN_11 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_header_5 : io_pipe_phv_in_header_5; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [15:0] _GEN_12 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_header_6 : io_pipe_phv_in_header_6; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [15:0] _GEN_13 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_header_7 : io_pipe_phv_in_header_7; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [15:0] _GEN_14 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_header_8 : io_pipe_phv_in_header_8; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [15:0] _GEN_15 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_header_9 : io_pipe_phv_in_header_9; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [15:0] _GEN_16 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_header_10 : io_pipe_phv_in_header_10; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [15:0] _GEN_17 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_header_11 : io_pipe_phv_in_header_11; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [15:0] _GEN_18 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_header_12 : io_pipe_phv_in_header_12; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [15:0] _GEN_19 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_header_13 : io_pipe_phv_in_header_13; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [15:0] _GEN_20 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_header_14 : io_pipe_phv_in_header_14; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [15:0] _GEN_21 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_header_15 : io_pipe_phv_in_header_15; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_22 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_0 : io_pipe_phv_in_data_0; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_23 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_1 : io_pipe_phv_in_data_1; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_24 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_2 : io_pipe_phv_in_data_2; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_25 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_3 : io_pipe_phv_in_data_3; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_26 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_4 : io_pipe_phv_in_data_4; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_27 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_5 : io_pipe_phv_in_data_5; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_28 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_6 : io_pipe_phv_in_data_6; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_29 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_7 : io_pipe_phv_in_data_7; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_30 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_8 : io_pipe_phv_in_data_8; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_31 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_9 : io_pipe_phv_in_data_9; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_32 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_10 : io_pipe_phv_in_data_10; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_33 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_11 : io_pipe_phv_in_data_11; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_34 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_12 : io_pipe_phv_in_data_12; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_35 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_13 : io_pipe_phv_in_data_13; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_36 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_14 : io_pipe_phv_in_data_14; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_37 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_15 : io_pipe_phv_in_data_15; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_38 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_16 : io_pipe_phv_in_data_16; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_39 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_17 : io_pipe_phv_in_data_17; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_40 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_18 : io_pipe_phv_in_data_18; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_41 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_19 : io_pipe_phv_in_data_19; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_42 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_20 : io_pipe_phv_in_data_20; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_43 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_21 : io_pipe_phv_in_data_21; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_44 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_22 : io_pipe_phv_in_data_22; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_45 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_23 : io_pipe_phv_in_data_23; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_46 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_24 : io_pipe_phv_in_data_24; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_47 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_25 : io_pipe_phv_in_data_25; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_48 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_26 : io_pipe_phv_in_data_26; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_49 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_27 : io_pipe_phv_in_data_27; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_50 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_28 : io_pipe_phv_in_data_28; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_51 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_29 : io_pipe_phv_in_data_29; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_52 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_30 : io_pipe_phv_in_data_30; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_53 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_31 : io_pipe_phv_in_data_31; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_54 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_32 : io_pipe_phv_in_data_32; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_55 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_33 : io_pipe_phv_in_data_33; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_56 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_34 : io_pipe_phv_in_data_34; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_57 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_35 : io_pipe_phv_in_data_35; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_58 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_36 : io_pipe_phv_in_data_36; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_59 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_37 : io_pipe_phv_in_data_37; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_60 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_38 : io_pipe_phv_in_data_38; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_61 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_39 : io_pipe_phv_in_data_39; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_62 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_40 : io_pipe_phv_in_data_40; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_63 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_41 : io_pipe_phv_in_data_41; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_64 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_42 : io_pipe_phv_in_data_42; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_65 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_43 : io_pipe_phv_in_data_43; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_66 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_44 : io_pipe_phv_in_data_44; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_67 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_45 : io_pipe_phv_in_data_45; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_68 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_46 : io_pipe_phv_in_data_46; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_69 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_47 : io_pipe_phv_in_data_47; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_70 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_48 : io_pipe_phv_in_data_48; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_71 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_49 : io_pipe_phv_in_data_49; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_72 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_50 : io_pipe_phv_in_data_50; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_73 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_51 : io_pipe_phv_in_data_51; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_74 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_52 : io_pipe_phv_in_data_52; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_75 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_53 : io_pipe_phv_in_data_53; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_76 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_54 : io_pipe_phv_in_data_54; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_77 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_55 : io_pipe_phv_in_data_55; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_78 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_56 : io_pipe_phv_in_data_56; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_79 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_57 : io_pipe_phv_in_data_57; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_80 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_58 : io_pipe_phv_in_data_58; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_81 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_59 : io_pipe_phv_in_data_59; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_82 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_60 : io_pipe_phv_in_data_60; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_83 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_61 : io_pipe_phv_in_data_61; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_84 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_62 : io_pipe_phv_in_data_62; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_85 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_63 : io_pipe_phv_in_data_63; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_86 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_64 : io_pipe_phv_in_data_64; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_87 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_65 : io_pipe_phv_in_data_65; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_88 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_66 : io_pipe_phv_in_data_66; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_89 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_67 : io_pipe_phv_in_data_67; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_90 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_68 : io_pipe_phv_in_data_68; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_91 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_69 : io_pipe_phv_in_data_69; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_92 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_70 : io_pipe_phv_in_data_70; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_93 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_71 : io_pipe_phv_in_data_71; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_94 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_72 : io_pipe_phv_in_data_72; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_95 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_73 : io_pipe_phv_in_data_73; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_96 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_74 : io_pipe_phv_in_data_74; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_97 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_75 : io_pipe_phv_in_data_75; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_98 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_76 : io_pipe_phv_in_data_76; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_99 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_77 : io_pipe_phv_in_data_77; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_100 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_78 : io_pipe_phv_in_data_78; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_101 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_79 : io_pipe_phv_in_data_79; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_102 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_80 : io_pipe_phv_in_data_80; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_103 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_81 : io_pipe_phv_in_data_81; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_104 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_82 : io_pipe_phv_in_data_82; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_105 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_83 : io_pipe_phv_in_data_83; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_106 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_84 : io_pipe_phv_in_data_84; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_107 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_85 : io_pipe_phv_in_data_85; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_108 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_86 : io_pipe_phv_in_data_86; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_109 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_87 : io_pipe_phv_in_data_87; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_110 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_88 : io_pipe_phv_in_data_88; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_111 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_89 : io_pipe_phv_in_data_89; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_112 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_90 : io_pipe_phv_in_data_90; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_113 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_91 : io_pipe_phv_in_data_91; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_114 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_92 : io_pipe_phv_in_data_92; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_115 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_93 : io_pipe_phv_in_data_93; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_116 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_94 : io_pipe_phv_in_data_94; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_117 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_95 : io_pipe_phv_in_data_95; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_118 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_96 : io_pipe_phv_in_data_96; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_119 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_97 : io_pipe_phv_in_data_97; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_120 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_98 : io_pipe_phv_in_data_98; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_121 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_99 : io_pipe_phv_in_data_99; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_122 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_100 : io_pipe_phv_in_data_100; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_123 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_101 : io_pipe_phv_in_data_101; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_124 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_102 : io_pipe_phv_in_data_102; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_125 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_103 : io_pipe_phv_in_data_103; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_126 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_104 : io_pipe_phv_in_data_104; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_127 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_105 : io_pipe_phv_in_data_105; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_128 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_106 : io_pipe_phv_in_data_106; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_129 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_107 : io_pipe_phv_in_data_107; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_130 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_108 : io_pipe_phv_in_data_108; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_131 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_109 : io_pipe_phv_in_data_109; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_132 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_110 : io_pipe_phv_in_data_110; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_133 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_111 : io_pipe_phv_in_data_111; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_134 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_112 : io_pipe_phv_in_data_112; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_135 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_113 : io_pipe_phv_in_data_113; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_136 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_114 : io_pipe_phv_in_data_114; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_137 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_115 : io_pipe_phv_in_data_115; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_138 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_116 : io_pipe_phv_in_data_116; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_139 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_117 : io_pipe_phv_in_data_117; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_140 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_118 : io_pipe_phv_in_data_118; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_141 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_119 : io_pipe_phv_in_data_119; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_142 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_120 : io_pipe_phv_in_data_120; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_143 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_121 : io_pipe_phv_in_data_121; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_144 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_122 : io_pipe_phv_in_data_122; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_145 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_123 : io_pipe_phv_in_data_123; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_146 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_124 : io_pipe_phv_in_data_124; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_147 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_125 : io_pipe_phv_in_data_125; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_148 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_126 : io_pipe_phv_in_data_126; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_149 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_127 : io_pipe_phv_in_data_127; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_150 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_128 : io_pipe_phv_in_data_128; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_151 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_129 : io_pipe_phv_in_data_129; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_152 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_130 : io_pipe_phv_in_data_130; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_153 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_131 : io_pipe_phv_in_data_131; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_154 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_132 : io_pipe_phv_in_data_132; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_155 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_133 : io_pipe_phv_in_data_133; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_156 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_134 : io_pipe_phv_in_data_134; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_157 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_135 : io_pipe_phv_in_data_135; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_158 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_136 : io_pipe_phv_in_data_136; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_159 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_137 : io_pipe_phv_in_data_137; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_160 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_138 : io_pipe_phv_in_data_138; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_161 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_139 : io_pipe_phv_in_data_139; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_162 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_140 : io_pipe_phv_in_data_140; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_163 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_141 : io_pipe_phv_in_data_141; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_164 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_142 : io_pipe_phv_in_data_142; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_165 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_143 : io_pipe_phv_in_data_143; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_166 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_144 : io_pipe_phv_in_data_144; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_167 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_145 : io_pipe_phv_in_data_145; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_168 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_146 : io_pipe_phv_in_data_146; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_169 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_147 : io_pipe_phv_in_data_147; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_170 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_148 : io_pipe_phv_in_data_148; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_171 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_149 : io_pipe_phv_in_data_149; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_172 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_150 : io_pipe_phv_in_data_150; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_173 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_151 : io_pipe_phv_in_data_151; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_174 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_152 : io_pipe_phv_in_data_152; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_175 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_153 : io_pipe_phv_in_data_153; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_176 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_154 : io_pipe_phv_in_data_154; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_177 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_155 : io_pipe_phv_in_data_155; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_178 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_156 : io_pipe_phv_in_data_156; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_179 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_157 : io_pipe_phv_in_data_157; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_180 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_158 : io_pipe_phv_in_data_158; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_181 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_159 : io_pipe_phv_in_data_159; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_182 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_160 : io_pipe_phv_in_data_160; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_183 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_161 : io_pipe_phv_in_data_161; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_184 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_162 : io_pipe_phv_in_data_162; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_185 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_163 : io_pipe_phv_in_data_163; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_186 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_164 : io_pipe_phv_in_data_164; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_187 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_165 : io_pipe_phv_in_data_165; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_188 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_166 : io_pipe_phv_in_data_166; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_189 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_167 : io_pipe_phv_in_data_167; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_190 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_168 : io_pipe_phv_in_data_168; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_191 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_169 : io_pipe_phv_in_data_169; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_192 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_170 : io_pipe_phv_in_data_170; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_193 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_171 : io_pipe_phv_in_data_171; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_194 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_172 : io_pipe_phv_in_data_172; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_195 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_173 : io_pipe_phv_in_data_173; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_196 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_174 : io_pipe_phv_in_data_174; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_197 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_175 : io_pipe_phv_in_data_175; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_198 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_176 : io_pipe_phv_in_data_176; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_199 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_177 : io_pipe_phv_in_data_177; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_200 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_178 : io_pipe_phv_in_data_178; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_201 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_179 : io_pipe_phv_in_data_179; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_202 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_180 : io_pipe_phv_in_data_180; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_203 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_181 : io_pipe_phv_in_data_181; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_204 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_182 : io_pipe_phv_in_data_182; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_205 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_183 : io_pipe_phv_in_data_183; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_206 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_184 : io_pipe_phv_in_data_184; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_207 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_185 : io_pipe_phv_in_data_185; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_208 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_186 : io_pipe_phv_in_data_186; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_209 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_187 : io_pipe_phv_in_data_187; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_210 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_188 : io_pipe_phv_in_data_188; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_211 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_189 : io_pipe_phv_in_data_189; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_212 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_190 : io_pipe_phv_in_data_190; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_213 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_191 : io_pipe_phv_in_data_191; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_214 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_192 : io_pipe_phv_in_data_192; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_215 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_193 : io_pipe_phv_in_data_193; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_216 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_194 : io_pipe_phv_in_data_194; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_217 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_195 : io_pipe_phv_in_data_195; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_218 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_196 : io_pipe_phv_in_data_196; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_219 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_197 : io_pipe_phv_in_data_197; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_220 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_198 : io_pipe_phv_in_data_198; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_221 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_199 : io_pipe_phv_in_data_199; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_222 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_200 : io_pipe_phv_in_data_200; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_223 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_201 : io_pipe_phv_in_data_201; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_224 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_202 : io_pipe_phv_in_data_202; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_225 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_203 : io_pipe_phv_in_data_203; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_226 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_204 : io_pipe_phv_in_data_204; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_227 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_205 : io_pipe_phv_in_data_205; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_228 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_206 : io_pipe_phv_in_data_206; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_229 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_207 : io_pipe_phv_in_data_207; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_230 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_208 : io_pipe_phv_in_data_208; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_231 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_209 : io_pipe_phv_in_data_209; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_232 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_210 : io_pipe_phv_in_data_210; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_233 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_211 : io_pipe_phv_in_data_211; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_234 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_212 : io_pipe_phv_in_data_212; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_235 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_213 : io_pipe_phv_in_data_213; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_236 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_214 : io_pipe_phv_in_data_214; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_237 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_215 : io_pipe_phv_in_data_215; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_238 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_216 : io_pipe_phv_in_data_216; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_239 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_217 : io_pipe_phv_in_data_217; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_240 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_218 : io_pipe_phv_in_data_218; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_241 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_219 : io_pipe_phv_in_data_219; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_242 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_220 : io_pipe_phv_in_data_220; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_243 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_221 : io_pipe_phv_in_data_221; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_244 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_222 : io_pipe_phv_in_data_222; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_245 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_223 : io_pipe_phv_in_data_223; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_246 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_224 : io_pipe_phv_in_data_224; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_247 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_225 : io_pipe_phv_in_data_225; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_248 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_226 : io_pipe_phv_in_data_226; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_249 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_227 : io_pipe_phv_in_data_227; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_250 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_228 : io_pipe_phv_in_data_228; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_251 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_229 : io_pipe_phv_in_data_229; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_252 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_230 : io_pipe_phv_in_data_230; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_253 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_231 : io_pipe_phv_in_data_231; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_254 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_232 : io_pipe_phv_in_data_232; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_255 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_233 : io_pipe_phv_in_data_233; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_256 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_234 : io_pipe_phv_in_data_234; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_257 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_235 : io_pipe_phv_in_data_235; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_258 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_236 : io_pipe_phv_in_data_236; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_259 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_237 : io_pipe_phv_in_data_237; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_260 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_238 : io_pipe_phv_in_data_238; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_261 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_239 : io_pipe_phv_in_data_239; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_262 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_240 : io_pipe_phv_in_data_240; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_263 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_241 : io_pipe_phv_in_data_241; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_264 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_242 : io_pipe_phv_in_data_242; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_265 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_243 : io_pipe_phv_in_data_243; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_266 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_244 : io_pipe_phv_in_data_244; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_267 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_245 : io_pipe_phv_in_data_245; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_268 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_246 : io_pipe_phv_in_data_246; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_269 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_247 : io_pipe_phv_in_data_247; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_270 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_248 : io_pipe_phv_in_data_248; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_271 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_249 : io_pipe_phv_in_data_249; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_272 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_250 : io_pipe_phv_in_data_250; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_273 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_251 : io_pipe_phv_in_data_251; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_274 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_252 : io_pipe_phv_in_data_252; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_275 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_253 : io_pipe_phv_in_data_253; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_276 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_254 : io_pipe_phv_in_data_254; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_277 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_255 : io_pipe_phv_in_data_255; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire  _GEN_278 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_is_valid_processor : _GEN_0; // @[parser.scala 33:62 parser.scala 34:35]
  wire  _GEN_279 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_next_config_id : _GEN_1; // @[parser.scala 33:62 parser.scala 34:35]
  wire [2:0] _GEN_280 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_next_processor_id : _GEN_2; // @[parser.scala 33:62 parser.scala 34:35]
  wire [15:0] _GEN_281 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_parse_transition_field : _GEN_3; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_282 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_parse_current_offset : _GEN_4; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_283 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_parse_current_state : _GEN_5; // @[parser.scala 33:62 parser.scala 34:35]
  wire [15:0] _GEN_284 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_header_0 : _GEN_6; // @[parser.scala 33:62 parser.scala 34:35]
  wire [15:0] _GEN_285 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_header_1 : _GEN_7; // @[parser.scala 33:62 parser.scala 34:35]
  wire [15:0] _GEN_286 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_header_2 : _GEN_8; // @[parser.scala 33:62 parser.scala 34:35]
  wire [15:0] _GEN_287 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_header_3 : _GEN_9; // @[parser.scala 33:62 parser.scala 34:35]
  wire [15:0] _GEN_288 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_header_4 : _GEN_10; // @[parser.scala 33:62 parser.scala 34:35]
  wire [15:0] _GEN_289 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_header_5 : _GEN_11; // @[parser.scala 33:62 parser.scala 34:35]
  wire [15:0] _GEN_290 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_header_6 : _GEN_12; // @[parser.scala 33:62 parser.scala 34:35]
  wire [15:0] _GEN_291 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_header_7 : _GEN_13; // @[parser.scala 33:62 parser.scala 34:35]
  wire [15:0] _GEN_292 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_header_8 : _GEN_14; // @[parser.scala 33:62 parser.scala 34:35]
  wire [15:0] _GEN_293 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_header_9 : _GEN_15; // @[parser.scala 33:62 parser.scala 34:35]
  wire [15:0] _GEN_294 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_header_10 : _GEN_16; // @[parser.scala 33:62 parser.scala 34:35]
  wire [15:0] _GEN_295 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_header_11 : _GEN_17; // @[parser.scala 33:62 parser.scala 34:35]
  wire [15:0] _GEN_296 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_header_12 : _GEN_18; // @[parser.scala 33:62 parser.scala 34:35]
  wire [15:0] _GEN_297 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_header_13 : _GEN_19; // @[parser.scala 33:62 parser.scala 34:35]
  wire [15:0] _GEN_298 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_header_14 : _GEN_20; // @[parser.scala 33:62 parser.scala 34:35]
  wire [15:0] _GEN_299 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_header_15 : _GEN_21; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_300 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_0 : _GEN_22; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_301 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_1 : _GEN_23; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_302 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_2 : _GEN_24; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_303 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_3 : _GEN_25; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_304 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_4 : _GEN_26; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_305 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_5 : _GEN_27; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_306 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_6 : _GEN_28; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_307 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_7 : _GEN_29; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_308 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_8 : _GEN_30; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_309 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_9 : _GEN_31; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_310 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_10 : _GEN_32; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_311 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_11 : _GEN_33; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_312 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_12 : _GEN_34; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_313 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_13 : _GEN_35; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_314 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_14 : _GEN_36; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_315 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_15 : _GEN_37; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_316 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_16 : _GEN_38; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_317 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_17 : _GEN_39; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_318 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_18 : _GEN_40; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_319 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_19 : _GEN_41; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_320 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_20 : _GEN_42; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_321 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_21 : _GEN_43; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_322 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_22 : _GEN_44; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_323 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_23 : _GEN_45; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_324 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_24 : _GEN_46; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_325 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_25 : _GEN_47; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_326 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_26 : _GEN_48; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_327 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_27 : _GEN_49; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_328 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_28 : _GEN_50; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_329 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_29 : _GEN_51; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_330 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_30 : _GEN_52; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_331 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_31 : _GEN_53; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_332 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_32 : _GEN_54; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_333 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_33 : _GEN_55; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_334 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_34 : _GEN_56; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_335 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_35 : _GEN_57; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_336 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_36 : _GEN_58; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_337 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_37 : _GEN_59; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_338 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_38 : _GEN_60; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_339 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_39 : _GEN_61; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_340 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_40 : _GEN_62; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_341 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_41 : _GEN_63; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_342 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_42 : _GEN_64; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_343 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_43 : _GEN_65; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_344 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_44 : _GEN_66; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_345 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_45 : _GEN_67; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_346 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_46 : _GEN_68; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_347 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_47 : _GEN_69; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_348 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_48 : _GEN_70; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_349 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_49 : _GEN_71; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_350 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_50 : _GEN_72; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_351 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_51 : _GEN_73; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_352 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_52 : _GEN_74; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_353 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_53 : _GEN_75; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_354 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_54 : _GEN_76; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_355 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_55 : _GEN_77; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_356 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_56 : _GEN_78; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_357 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_57 : _GEN_79; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_358 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_58 : _GEN_80; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_359 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_59 : _GEN_81; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_360 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_60 : _GEN_82; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_361 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_61 : _GEN_83; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_362 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_62 : _GEN_84; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_363 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_63 : _GEN_85; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_364 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_64 : _GEN_86; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_365 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_65 : _GEN_87; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_366 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_66 : _GEN_88; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_367 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_67 : _GEN_89; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_368 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_68 : _GEN_90; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_369 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_69 : _GEN_91; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_370 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_70 : _GEN_92; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_371 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_71 : _GEN_93; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_372 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_72 : _GEN_94; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_373 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_73 : _GEN_95; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_374 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_74 : _GEN_96; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_375 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_75 : _GEN_97; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_376 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_76 : _GEN_98; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_377 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_77 : _GEN_99; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_378 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_78 : _GEN_100; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_379 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_79 : _GEN_101; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_380 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_80 : _GEN_102; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_381 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_81 : _GEN_103; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_382 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_82 : _GEN_104; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_383 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_83 : _GEN_105; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_384 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_84 : _GEN_106; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_385 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_85 : _GEN_107; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_386 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_86 : _GEN_108; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_387 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_87 : _GEN_109; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_388 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_88 : _GEN_110; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_389 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_89 : _GEN_111; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_390 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_90 : _GEN_112; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_391 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_91 : _GEN_113; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_392 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_92 : _GEN_114; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_393 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_93 : _GEN_115; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_394 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_94 : _GEN_116; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_395 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_95 : _GEN_117; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_396 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_96 : _GEN_118; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_397 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_97 : _GEN_119; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_398 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_98 : _GEN_120; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_399 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_99 : _GEN_121; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_400 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_100 : _GEN_122; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_401 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_101 : _GEN_123; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_402 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_102 : _GEN_124; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_403 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_103 : _GEN_125; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_404 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_104 : _GEN_126; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_405 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_105 : _GEN_127; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_406 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_106 : _GEN_128; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_407 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_107 : _GEN_129; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_408 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_108 : _GEN_130; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_409 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_109 : _GEN_131; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_410 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_110 : _GEN_132; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_411 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_111 : _GEN_133; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_412 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_112 : _GEN_134; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_413 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_113 : _GEN_135; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_414 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_114 : _GEN_136; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_415 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_115 : _GEN_137; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_416 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_116 : _GEN_138; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_417 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_117 : _GEN_139; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_418 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_118 : _GEN_140; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_419 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_119 : _GEN_141; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_420 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_120 : _GEN_142; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_421 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_121 : _GEN_143; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_422 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_122 : _GEN_144; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_423 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_123 : _GEN_145; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_424 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_124 : _GEN_146; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_425 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_125 : _GEN_147; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_426 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_126 : _GEN_148; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_427 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_127 : _GEN_149; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_428 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_128 : _GEN_150; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_429 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_129 : _GEN_151; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_430 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_130 : _GEN_152; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_431 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_131 : _GEN_153; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_432 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_132 : _GEN_154; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_433 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_133 : _GEN_155; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_434 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_134 : _GEN_156; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_435 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_135 : _GEN_157; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_436 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_136 : _GEN_158; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_437 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_137 : _GEN_159; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_438 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_138 : _GEN_160; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_439 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_139 : _GEN_161; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_440 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_140 : _GEN_162; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_441 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_141 : _GEN_163; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_442 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_142 : _GEN_164; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_443 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_143 : _GEN_165; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_444 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_144 : _GEN_166; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_445 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_145 : _GEN_167; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_446 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_146 : _GEN_168; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_447 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_147 : _GEN_169; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_448 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_148 : _GEN_170; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_449 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_149 : _GEN_171; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_450 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_150 : _GEN_172; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_451 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_151 : _GEN_173; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_452 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_152 : _GEN_174; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_453 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_153 : _GEN_175; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_454 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_154 : _GEN_176; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_455 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_155 : _GEN_177; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_456 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_156 : _GEN_178; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_457 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_157 : _GEN_179; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_458 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_158 : _GEN_180; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_459 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_159 : _GEN_181; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_460 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_160 : _GEN_182; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_461 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_161 : _GEN_183; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_462 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_162 : _GEN_184; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_463 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_163 : _GEN_185; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_464 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_164 : _GEN_186; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_465 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_165 : _GEN_187; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_466 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_166 : _GEN_188; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_467 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_167 : _GEN_189; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_468 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_168 : _GEN_190; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_469 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_169 : _GEN_191; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_470 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_170 : _GEN_192; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_471 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_171 : _GEN_193; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_472 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_172 : _GEN_194; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_473 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_173 : _GEN_195; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_474 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_174 : _GEN_196; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_475 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_175 : _GEN_197; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_476 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_176 : _GEN_198; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_477 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_177 : _GEN_199; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_478 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_178 : _GEN_200; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_479 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_179 : _GEN_201; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_480 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_180 : _GEN_202; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_481 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_181 : _GEN_203; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_482 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_182 : _GEN_204; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_483 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_183 : _GEN_205; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_484 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_184 : _GEN_206; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_485 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_185 : _GEN_207; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_486 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_186 : _GEN_208; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_487 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_187 : _GEN_209; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_488 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_188 : _GEN_210; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_489 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_189 : _GEN_211; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_490 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_190 : _GEN_212; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_491 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_191 : _GEN_213; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_492 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_192 : _GEN_214; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_493 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_193 : _GEN_215; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_494 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_194 : _GEN_216; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_495 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_195 : _GEN_217; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_496 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_196 : _GEN_218; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_497 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_197 : _GEN_219; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_498 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_198 : _GEN_220; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_499 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_199 : _GEN_221; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_500 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_200 : _GEN_222; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_501 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_201 : _GEN_223; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_502 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_202 : _GEN_224; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_503 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_203 : _GEN_225; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_504 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_204 : _GEN_226; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_505 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_205 : _GEN_227; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_506 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_206 : _GEN_228; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_507 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_207 : _GEN_229; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_508 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_208 : _GEN_230; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_509 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_209 : _GEN_231; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_510 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_210 : _GEN_232; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_511 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_211 : _GEN_233; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_512 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_212 : _GEN_234; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_513 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_213 : _GEN_235; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_514 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_214 : _GEN_236; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_515 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_215 : _GEN_237; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_516 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_216 : _GEN_238; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_517 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_217 : _GEN_239; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_518 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_218 : _GEN_240; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_519 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_219 : _GEN_241; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_520 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_220 : _GEN_242; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_521 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_221 : _GEN_243; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_522 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_222 : _GEN_244; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_523 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_223 : _GEN_245; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_524 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_224 : _GEN_246; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_525 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_225 : _GEN_247; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_526 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_226 : _GEN_248; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_527 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_227 : _GEN_249; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_528 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_228 : _GEN_250; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_529 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_229 : _GEN_251; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_530 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_230 : _GEN_252; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_531 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_231 : _GEN_253; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_532 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_232 : _GEN_254; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_533 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_233 : _GEN_255; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_534 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_234 : _GEN_256; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_535 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_235 : _GEN_257; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_536 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_236 : _GEN_258; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_537 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_237 : _GEN_259; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_538 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_238 : _GEN_260; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_539 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_239 : _GEN_261; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_540 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_240 : _GEN_262; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_541 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_241 : _GEN_263; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_542 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_242 : _GEN_264; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_543 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_243 : _GEN_265; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_544 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_244 : _GEN_266; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_545 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_245 : _GEN_267; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_546 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_246 : _GEN_268; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_547 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_247 : _GEN_269; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_548 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_248 : _GEN_270; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_549 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_249 : _GEN_271; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_550 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_250 : _GEN_272; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_551 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_251 : _GEN_273; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_552 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_252 : _GEN_274; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_553 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_253 : _GEN_275; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_554 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_254 : _GEN_276; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_555 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_255 : _GEN_277; // @[parser.scala 33:62 parser.scala 34:35]
  wire  mod_j = io_mod_cs == 2'h0; // @[parser.scala 46:35]
  wire  mod_j_1 = io_mod_cs == 2'h1; // @[parser.scala 46:35]
  wire  mod_j_2 = io_mod_cs == 2'h2; // @[parser.scala 46:35]
  wire  mod_j_3 = io_mod_cs == 2'h3; // @[parser.scala 46:35]
  ParseModule mau_0 ( // @[parser.scala 21:25]
    .clock(mau_0_clock),
    .io_pipe_phv_in_data_0(mau_0_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(mau_0_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(mau_0_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(mau_0_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(mau_0_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(mau_0_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(mau_0_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(mau_0_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(mau_0_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(mau_0_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(mau_0_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(mau_0_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(mau_0_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(mau_0_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(mau_0_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(mau_0_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(mau_0_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(mau_0_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(mau_0_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(mau_0_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(mau_0_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(mau_0_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(mau_0_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(mau_0_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(mau_0_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(mau_0_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(mau_0_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(mau_0_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(mau_0_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(mau_0_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(mau_0_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(mau_0_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(mau_0_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(mau_0_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(mau_0_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(mau_0_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(mau_0_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(mau_0_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(mau_0_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(mau_0_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(mau_0_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(mau_0_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(mau_0_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(mau_0_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(mau_0_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(mau_0_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(mau_0_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(mau_0_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(mau_0_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(mau_0_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(mau_0_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(mau_0_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(mau_0_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(mau_0_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(mau_0_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(mau_0_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(mau_0_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(mau_0_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(mau_0_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(mau_0_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(mau_0_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(mau_0_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(mau_0_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(mau_0_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(mau_0_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(mau_0_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(mau_0_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(mau_0_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(mau_0_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(mau_0_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(mau_0_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(mau_0_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(mau_0_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(mau_0_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(mau_0_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(mau_0_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(mau_0_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(mau_0_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(mau_0_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(mau_0_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(mau_0_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(mau_0_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(mau_0_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(mau_0_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(mau_0_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(mau_0_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(mau_0_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(mau_0_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(mau_0_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(mau_0_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(mau_0_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(mau_0_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(mau_0_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(mau_0_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(mau_0_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(mau_0_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(mau_0_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(mau_0_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(mau_0_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(mau_0_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(mau_0_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(mau_0_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(mau_0_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(mau_0_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(mau_0_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(mau_0_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(mau_0_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(mau_0_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(mau_0_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(mau_0_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(mau_0_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(mau_0_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(mau_0_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(mau_0_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(mau_0_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(mau_0_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(mau_0_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(mau_0_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(mau_0_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(mau_0_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(mau_0_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(mau_0_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(mau_0_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(mau_0_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(mau_0_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(mau_0_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(mau_0_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(mau_0_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(mau_0_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(mau_0_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(mau_0_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(mau_0_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(mau_0_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(mau_0_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(mau_0_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(mau_0_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(mau_0_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(mau_0_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(mau_0_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(mau_0_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(mau_0_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(mau_0_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(mau_0_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(mau_0_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(mau_0_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(mau_0_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(mau_0_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(mau_0_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(mau_0_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(mau_0_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(mau_0_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(mau_0_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(mau_0_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(mau_0_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(mau_0_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(mau_0_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(mau_0_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(mau_0_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(mau_0_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(mau_0_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(mau_0_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(mau_0_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(mau_0_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(mau_0_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(mau_0_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(mau_0_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(mau_0_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(mau_0_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(mau_0_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(mau_0_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(mau_0_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(mau_0_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(mau_0_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(mau_0_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(mau_0_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(mau_0_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(mau_0_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(mau_0_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(mau_0_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(mau_0_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(mau_0_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(mau_0_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(mau_0_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(mau_0_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(mau_0_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(mau_0_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(mau_0_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(mau_0_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(mau_0_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(mau_0_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(mau_0_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(mau_0_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(mau_0_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(mau_0_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(mau_0_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(mau_0_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(mau_0_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(mau_0_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(mau_0_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(mau_0_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(mau_0_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(mau_0_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(mau_0_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(mau_0_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(mau_0_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(mau_0_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(mau_0_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(mau_0_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(mau_0_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(mau_0_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(mau_0_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(mau_0_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(mau_0_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(mau_0_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(mau_0_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(mau_0_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(mau_0_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(mau_0_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(mau_0_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(mau_0_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(mau_0_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(mau_0_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(mau_0_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(mau_0_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(mau_0_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(mau_0_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(mau_0_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(mau_0_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(mau_0_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(mau_0_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(mau_0_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(mau_0_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(mau_0_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(mau_0_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(mau_0_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(mau_0_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(mau_0_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(mau_0_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(mau_0_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(mau_0_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(mau_0_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(mau_0_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(mau_0_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(mau_0_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(mau_0_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(mau_0_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(mau_0_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(mau_0_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(mau_0_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(mau_0_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(mau_0_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(mau_0_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(mau_0_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(mau_0_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(mau_0_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(mau_0_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_header_0(mau_0_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(mau_0_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(mau_0_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(mau_0_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(mau_0_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(mau_0_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(mau_0_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(mau_0_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(mau_0_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(mau_0_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(mau_0_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(mau_0_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(mau_0_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(mau_0_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(mau_0_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(mau_0_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(mau_0_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(mau_0_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(mau_0_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(mau_0_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(mau_0_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(mau_0_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(mau_0_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(mau_0_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(mau_0_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(mau_0_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(mau_0_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(mau_0_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(mau_0_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(mau_0_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(mau_0_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(mau_0_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(mau_0_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(mau_0_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(mau_0_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(mau_0_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(mau_0_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(mau_0_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(mau_0_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(mau_0_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(mau_0_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(mau_0_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(mau_0_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(mau_0_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(mau_0_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(mau_0_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(mau_0_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(mau_0_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(mau_0_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(mau_0_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(mau_0_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(mau_0_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(mau_0_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(mau_0_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(mau_0_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(mau_0_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(mau_0_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(mau_0_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(mau_0_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(mau_0_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(mau_0_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(mau_0_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(mau_0_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(mau_0_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(mau_0_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(mau_0_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(mau_0_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(mau_0_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(mau_0_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(mau_0_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(mau_0_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(mau_0_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(mau_0_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(mau_0_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(mau_0_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(mau_0_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(mau_0_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(mau_0_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(mau_0_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(mau_0_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(mau_0_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(mau_0_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(mau_0_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(mau_0_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(mau_0_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(mau_0_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(mau_0_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(mau_0_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(mau_0_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(mau_0_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(mau_0_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(mau_0_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(mau_0_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(mau_0_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(mau_0_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(mau_0_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(mau_0_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(mau_0_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(mau_0_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(mau_0_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(mau_0_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(mau_0_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(mau_0_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(mau_0_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(mau_0_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(mau_0_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(mau_0_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(mau_0_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(mau_0_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(mau_0_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(mau_0_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(mau_0_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(mau_0_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(mau_0_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(mau_0_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(mau_0_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(mau_0_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(mau_0_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(mau_0_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(mau_0_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(mau_0_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(mau_0_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(mau_0_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(mau_0_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(mau_0_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(mau_0_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(mau_0_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(mau_0_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(mau_0_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(mau_0_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(mau_0_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(mau_0_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(mau_0_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(mau_0_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(mau_0_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(mau_0_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(mau_0_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(mau_0_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(mau_0_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(mau_0_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(mau_0_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(mau_0_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(mau_0_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(mau_0_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(mau_0_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(mau_0_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(mau_0_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(mau_0_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(mau_0_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(mau_0_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(mau_0_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(mau_0_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(mau_0_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(mau_0_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(mau_0_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(mau_0_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(mau_0_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(mau_0_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(mau_0_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(mau_0_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(mau_0_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(mau_0_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(mau_0_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(mau_0_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(mau_0_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(mau_0_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(mau_0_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(mau_0_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(mau_0_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(mau_0_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(mau_0_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(mau_0_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(mau_0_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(mau_0_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(mau_0_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(mau_0_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(mau_0_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(mau_0_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(mau_0_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(mau_0_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(mau_0_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(mau_0_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(mau_0_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(mau_0_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(mau_0_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(mau_0_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(mau_0_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(mau_0_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(mau_0_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(mau_0_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(mau_0_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(mau_0_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(mau_0_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(mau_0_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(mau_0_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(mau_0_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(mau_0_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(mau_0_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(mau_0_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(mau_0_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(mau_0_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(mau_0_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(mau_0_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(mau_0_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(mau_0_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(mau_0_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(mau_0_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(mau_0_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(mau_0_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(mau_0_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(mau_0_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(mau_0_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(mau_0_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(mau_0_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(mau_0_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(mau_0_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(mau_0_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(mau_0_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(mau_0_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(mau_0_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(mau_0_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(mau_0_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(mau_0_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(mau_0_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(mau_0_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(mau_0_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(mau_0_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(mau_0_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(mau_0_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(mau_0_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(mau_0_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(mau_0_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(mau_0_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(mau_0_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(mau_0_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(mau_0_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(mau_0_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(mau_0_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(mau_0_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(mau_0_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(mau_0_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(mau_0_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(mau_0_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(mau_0_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(mau_0_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(mau_0_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(mau_0_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(mau_0_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(mau_0_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(mau_0_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(mau_0_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(mau_0_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(mau_0_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(mau_0_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(mau_0_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(mau_0_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(mau_0_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(mau_0_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(mau_0_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(mau_0_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(mau_0_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(mau_0_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(mau_0_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(mau_0_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(mau_0_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(mau_0_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(mau_0_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(mau_0_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(mau_0_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(mau_0_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(mau_0_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(mau_0_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(mau_0_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(mau_0_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(mau_0_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(mau_0_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(mau_0_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(mau_0_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_header_0(mau_0_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(mau_0_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(mau_0_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(mau_0_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(mau_0_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(mau_0_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(mau_0_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(mau_0_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(mau_0_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(mau_0_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(mau_0_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(mau_0_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(mau_0_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(mau_0_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(mau_0_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(mau_0_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(mau_0_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(mau_0_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(mau_0_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(mau_0_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(mau_0_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(mau_0_io_pipe_phv_out_is_valid_processor),
    .io_mod_state_id_mod(mau_0_io_mod_state_id_mod),
    .io_mod_state_id(mau_0_io_mod_state_id),
    .io_mod_sram_w_cs(mau_0_io_mod_sram_w_cs),
    .io_mod_sram_w_en(mau_0_io_mod_sram_w_en),
    .io_mod_sram_w_addr(mau_0_io_mod_sram_w_addr),
    .io_mod_sram_w_data(mau_0_io_mod_sram_w_data)
  );
  ParseModule mau_1 ( // @[parser.scala 21:25]
    .clock(mau_1_clock),
    .io_pipe_phv_in_data_0(mau_1_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(mau_1_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(mau_1_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(mau_1_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(mau_1_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(mau_1_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(mau_1_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(mau_1_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(mau_1_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(mau_1_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(mau_1_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(mau_1_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(mau_1_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(mau_1_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(mau_1_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(mau_1_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(mau_1_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(mau_1_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(mau_1_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(mau_1_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(mau_1_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(mau_1_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(mau_1_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(mau_1_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(mau_1_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(mau_1_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(mau_1_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(mau_1_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(mau_1_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(mau_1_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(mau_1_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(mau_1_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(mau_1_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(mau_1_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(mau_1_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(mau_1_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(mau_1_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(mau_1_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(mau_1_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(mau_1_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(mau_1_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(mau_1_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(mau_1_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(mau_1_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(mau_1_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(mau_1_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(mau_1_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(mau_1_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(mau_1_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(mau_1_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(mau_1_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(mau_1_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(mau_1_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(mau_1_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(mau_1_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(mau_1_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(mau_1_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(mau_1_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(mau_1_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(mau_1_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(mau_1_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(mau_1_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(mau_1_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(mau_1_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(mau_1_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(mau_1_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(mau_1_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(mau_1_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(mau_1_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(mau_1_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(mau_1_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(mau_1_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(mau_1_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(mau_1_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(mau_1_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(mau_1_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(mau_1_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(mau_1_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(mau_1_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(mau_1_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(mau_1_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(mau_1_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(mau_1_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(mau_1_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(mau_1_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(mau_1_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(mau_1_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(mau_1_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(mau_1_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(mau_1_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(mau_1_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(mau_1_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(mau_1_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(mau_1_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(mau_1_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(mau_1_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(mau_1_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(mau_1_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(mau_1_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(mau_1_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(mau_1_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(mau_1_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(mau_1_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(mau_1_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(mau_1_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(mau_1_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(mau_1_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(mau_1_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(mau_1_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(mau_1_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(mau_1_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(mau_1_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(mau_1_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(mau_1_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(mau_1_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(mau_1_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(mau_1_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(mau_1_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(mau_1_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(mau_1_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(mau_1_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(mau_1_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(mau_1_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(mau_1_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(mau_1_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(mau_1_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(mau_1_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(mau_1_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(mau_1_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(mau_1_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(mau_1_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(mau_1_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(mau_1_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(mau_1_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(mau_1_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(mau_1_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(mau_1_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(mau_1_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(mau_1_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(mau_1_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(mau_1_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(mau_1_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(mau_1_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(mau_1_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(mau_1_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(mau_1_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(mau_1_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(mau_1_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(mau_1_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(mau_1_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(mau_1_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(mau_1_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(mau_1_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(mau_1_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(mau_1_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(mau_1_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(mau_1_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(mau_1_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(mau_1_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(mau_1_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(mau_1_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(mau_1_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(mau_1_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(mau_1_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(mau_1_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(mau_1_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(mau_1_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(mau_1_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(mau_1_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(mau_1_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(mau_1_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(mau_1_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(mau_1_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(mau_1_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(mau_1_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(mau_1_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(mau_1_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(mau_1_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(mau_1_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(mau_1_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(mau_1_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(mau_1_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(mau_1_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(mau_1_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(mau_1_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(mau_1_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(mau_1_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(mau_1_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(mau_1_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(mau_1_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(mau_1_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(mau_1_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(mau_1_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(mau_1_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(mau_1_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(mau_1_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(mau_1_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(mau_1_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(mau_1_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(mau_1_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(mau_1_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(mau_1_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(mau_1_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(mau_1_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(mau_1_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(mau_1_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(mau_1_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(mau_1_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(mau_1_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(mau_1_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(mau_1_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(mau_1_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(mau_1_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(mau_1_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(mau_1_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(mau_1_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(mau_1_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(mau_1_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(mau_1_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(mau_1_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(mau_1_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(mau_1_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(mau_1_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(mau_1_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(mau_1_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(mau_1_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(mau_1_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(mau_1_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(mau_1_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(mau_1_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(mau_1_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(mau_1_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(mau_1_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(mau_1_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(mau_1_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(mau_1_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(mau_1_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(mau_1_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(mau_1_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(mau_1_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(mau_1_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(mau_1_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(mau_1_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(mau_1_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(mau_1_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(mau_1_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(mau_1_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(mau_1_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(mau_1_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(mau_1_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(mau_1_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(mau_1_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(mau_1_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(mau_1_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(mau_1_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(mau_1_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_header_0(mau_1_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(mau_1_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(mau_1_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(mau_1_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(mau_1_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(mau_1_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(mau_1_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(mau_1_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(mau_1_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(mau_1_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(mau_1_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(mau_1_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(mau_1_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(mau_1_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(mau_1_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(mau_1_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(mau_1_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(mau_1_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(mau_1_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(mau_1_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(mau_1_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(mau_1_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(mau_1_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(mau_1_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(mau_1_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(mau_1_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(mau_1_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(mau_1_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(mau_1_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(mau_1_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(mau_1_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(mau_1_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(mau_1_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(mau_1_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(mau_1_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(mau_1_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(mau_1_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(mau_1_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(mau_1_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(mau_1_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(mau_1_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(mau_1_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(mau_1_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(mau_1_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(mau_1_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(mau_1_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(mau_1_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(mau_1_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(mau_1_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(mau_1_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(mau_1_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(mau_1_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(mau_1_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(mau_1_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(mau_1_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(mau_1_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(mau_1_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(mau_1_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(mau_1_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(mau_1_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(mau_1_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(mau_1_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(mau_1_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(mau_1_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(mau_1_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(mau_1_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(mau_1_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(mau_1_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(mau_1_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(mau_1_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(mau_1_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(mau_1_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(mau_1_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(mau_1_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(mau_1_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(mau_1_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(mau_1_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(mau_1_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(mau_1_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(mau_1_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(mau_1_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(mau_1_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(mau_1_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(mau_1_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(mau_1_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(mau_1_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(mau_1_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(mau_1_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(mau_1_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(mau_1_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(mau_1_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(mau_1_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(mau_1_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(mau_1_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(mau_1_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(mau_1_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(mau_1_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(mau_1_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(mau_1_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(mau_1_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(mau_1_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(mau_1_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(mau_1_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(mau_1_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(mau_1_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(mau_1_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(mau_1_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(mau_1_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(mau_1_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(mau_1_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(mau_1_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(mau_1_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(mau_1_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(mau_1_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(mau_1_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(mau_1_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(mau_1_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(mau_1_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(mau_1_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(mau_1_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(mau_1_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(mau_1_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(mau_1_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(mau_1_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(mau_1_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(mau_1_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(mau_1_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(mau_1_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(mau_1_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(mau_1_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(mau_1_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(mau_1_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(mau_1_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(mau_1_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(mau_1_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(mau_1_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(mau_1_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(mau_1_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(mau_1_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(mau_1_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(mau_1_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(mau_1_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(mau_1_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(mau_1_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(mau_1_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(mau_1_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(mau_1_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(mau_1_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(mau_1_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(mau_1_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(mau_1_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(mau_1_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(mau_1_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(mau_1_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(mau_1_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(mau_1_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(mau_1_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(mau_1_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(mau_1_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(mau_1_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(mau_1_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(mau_1_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(mau_1_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(mau_1_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(mau_1_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(mau_1_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(mau_1_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(mau_1_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(mau_1_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(mau_1_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(mau_1_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(mau_1_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(mau_1_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(mau_1_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(mau_1_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(mau_1_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(mau_1_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(mau_1_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(mau_1_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(mau_1_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(mau_1_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(mau_1_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(mau_1_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(mau_1_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(mau_1_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(mau_1_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(mau_1_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(mau_1_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(mau_1_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(mau_1_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(mau_1_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(mau_1_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(mau_1_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(mau_1_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(mau_1_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(mau_1_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(mau_1_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(mau_1_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(mau_1_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(mau_1_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(mau_1_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(mau_1_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(mau_1_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(mau_1_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(mau_1_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(mau_1_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(mau_1_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(mau_1_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(mau_1_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(mau_1_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(mau_1_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(mau_1_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(mau_1_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(mau_1_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(mau_1_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(mau_1_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(mau_1_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(mau_1_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(mau_1_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(mau_1_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(mau_1_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(mau_1_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(mau_1_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(mau_1_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(mau_1_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(mau_1_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(mau_1_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(mau_1_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(mau_1_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(mau_1_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(mau_1_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(mau_1_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(mau_1_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(mau_1_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(mau_1_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(mau_1_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(mau_1_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(mau_1_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(mau_1_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(mau_1_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(mau_1_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(mau_1_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(mau_1_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(mau_1_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(mau_1_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(mau_1_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(mau_1_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(mau_1_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(mau_1_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(mau_1_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(mau_1_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(mau_1_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(mau_1_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(mau_1_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(mau_1_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(mau_1_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(mau_1_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(mau_1_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(mau_1_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(mau_1_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(mau_1_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(mau_1_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(mau_1_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(mau_1_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(mau_1_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(mau_1_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(mau_1_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(mau_1_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(mau_1_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(mau_1_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(mau_1_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(mau_1_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(mau_1_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(mau_1_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(mau_1_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(mau_1_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(mau_1_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(mau_1_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_header_0(mau_1_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(mau_1_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(mau_1_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(mau_1_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(mau_1_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(mau_1_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(mau_1_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(mau_1_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(mau_1_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(mau_1_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(mau_1_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(mau_1_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(mau_1_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(mau_1_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(mau_1_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(mau_1_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(mau_1_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(mau_1_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(mau_1_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(mau_1_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(mau_1_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(mau_1_io_pipe_phv_out_is_valid_processor),
    .io_mod_state_id_mod(mau_1_io_mod_state_id_mod),
    .io_mod_state_id(mau_1_io_mod_state_id),
    .io_mod_sram_w_cs(mau_1_io_mod_sram_w_cs),
    .io_mod_sram_w_en(mau_1_io_mod_sram_w_en),
    .io_mod_sram_w_addr(mau_1_io_mod_sram_w_addr),
    .io_mod_sram_w_data(mau_1_io_mod_sram_w_data)
  );
  ParseModule mau_2 ( // @[parser.scala 21:25]
    .clock(mau_2_clock),
    .io_pipe_phv_in_data_0(mau_2_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(mau_2_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(mau_2_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(mau_2_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(mau_2_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(mau_2_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(mau_2_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(mau_2_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(mau_2_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(mau_2_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(mau_2_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(mau_2_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(mau_2_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(mau_2_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(mau_2_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(mau_2_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(mau_2_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(mau_2_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(mau_2_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(mau_2_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(mau_2_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(mau_2_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(mau_2_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(mau_2_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(mau_2_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(mau_2_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(mau_2_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(mau_2_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(mau_2_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(mau_2_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(mau_2_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(mau_2_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(mau_2_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(mau_2_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(mau_2_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(mau_2_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(mau_2_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(mau_2_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(mau_2_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(mau_2_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(mau_2_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(mau_2_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(mau_2_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(mau_2_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(mau_2_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(mau_2_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(mau_2_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(mau_2_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(mau_2_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(mau_2_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(mau_2_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(mau_2_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(mau_2_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(mau_2_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(mau_2_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(mau_2_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(mau_2_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(mau_2_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(mau_2_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(mau_2_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(mau_2_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(mau_2_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(mau_2_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(mau_2_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(mau_2_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(mau_2_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(mau_2_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(mau_2_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(mau_2_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(mau_2_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(mau_2_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(mau_2_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(mau_2_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(mau_2_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(mau_2_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(mau_2_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(mau_2_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(mau_2_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(mau_2_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(mau_2_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(mau_2_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(mau_2_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(mau_2_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(mau_2_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(mau_2_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(mau_2_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(mau_2_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(mau_2_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(mau_2_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(mau_2_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(mau_2_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(mau_2_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(mau_2_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(mau_2_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(mau_2_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(mau_2_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(mau_2_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(mau_2_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(mau_2_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(mau_2_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(mau_2_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(mau_2_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(mau_2_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(mau_2_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(mau_2_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(mau_2_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(mau_2_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(mau_2_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(mau_2_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(mau_2_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(mau_2_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(mau_2_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(mau_2_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(mau_2_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(mau_2_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(mau_2_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(mau_2_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(mau_2_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(mau_2_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(mau_2_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(mau_2_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(mau_2_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(mau_2_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(mau_2_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(mau_2_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(mau_2_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(mau_2_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(mau_2_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(mau_2_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(mau_2_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(mau_2_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(mau_2_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(mau_2_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(mau_2_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(mau_2_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(mau_2_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(mau_2_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(mau_2_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(mau_2_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(mau_2_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(mau_2_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(mau_2_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(mau_2_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(mau_2_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(mau_2_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(mau_2_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(mau_2_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(mau_2_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(mau_2_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(mau_2_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(mau_2_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(mau_2_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(mau_2_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(mau_2_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(mau_2_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(mau_2_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(mau_2_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(mau_2_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(mau_2_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(mau_2_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(mau_2_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(mau_2_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(mau_2_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(mau_2_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(mau_2_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(mau_2_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(mau_2_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(mau_2_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(mau_2_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(mau_2_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(mau_2_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(mau_2_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(mau_2_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(mau_2_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(mau_2_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(mau_2_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(mau_2_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(mau_2_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(mau_2_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(mau_2_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(mau_2_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(mau_2_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(mau_2_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(mau_2_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(mau_2_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(mau_2_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(mau_2_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(mau_2_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(mau_2_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(mau_2_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(mau_2_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(mau_2_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(mau_2_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(mau_2_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(mau_2_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(mau_2_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(mau_2_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(mau_2_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(mau_2_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(mau_2_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(mau_2_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(mau_2_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(mau_2_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(mau_2_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(mau_2_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(mau_2_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(mau_2_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(mau_2_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(mau_2_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(mau_2_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(mau_2_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(mau_2_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(mau_2_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(mau_2_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(mau_2_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(mau_2_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(mau_2_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(mau_2_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(mau_2_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(mau_2_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(mau_2_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(mau_2_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(mau_2_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(mau_2_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(mau_2_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(mau_2_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(mau_2_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(mau_2_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(mau_2_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(mau_2_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(mau_2_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(mau_2_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(mau_2_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(mau_2_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(mau_2_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(mau_2_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(mau_2_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(mau_2_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(mau_2_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(mau_2_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(mau_2_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(mau_2_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(mau_2_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(mau_2_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(mau_2_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(mau_2_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(mau_2_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(mau_2_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(mau_2_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(mau_2_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(mau_2_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(mau_2_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(mau_2_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(mau_2_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(mau_2_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(mau_2_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_header_0(mau_2_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(mau_2_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(mau_2_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(mau_2_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(mau_2_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(mau_2_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(mau_2_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(mau_2_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(mau_2_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(mau_2_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(mau_2_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(mau_2_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(mau_2_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(mau_2_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(mau_2_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(mau_2_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(mau_2_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(mau_2_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(mau_2_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(mau_2_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(mau_2_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(mau_2_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(mau_2_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(mau_2_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(mau_2_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(mau_2_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(mau_2_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(mau_2_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(mau_2_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(mau_2_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(mau_2_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(mau_2_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(mau_2_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(mau_2_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(mau_2_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(mau_2_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(mau_2_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(mau_2_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(mau_2_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(mau_2_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(mau_2_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(mau_2_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(mau_2_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(mau_2_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(mau_2_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(mau_2_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(mau_2_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(mau_2_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(mau_2_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(mau_2_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(mau_2_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(mau_2_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(mau_2_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(mau_2_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(mau_2_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(mau_2_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(mau_2_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(mau_2_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(mau_2_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(mau_2_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(mau_2_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(mau_2_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(mau_2_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(mau_2_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(mau_2_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(mau_2_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(mau_2_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(mau_2_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(mau_2_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(mau_2_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(mau_2_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(mau_2_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(mau_2_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(mau_2_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(mau_2_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(mau_2_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(mau_2_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(mau_2_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(mau_2_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(mau_2_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(mau_2_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(mau_2_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(mau_2_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(mau_2_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(mau_2_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(mau_2_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(mau_2_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(mau_2_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(mau_2_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(mau_2_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(mau_2_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(mau_2_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(mau_2_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(mau_2_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(mau_2_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(mau_2_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(mau_2_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(mau_2_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(mau_2_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(mau_2_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(mau_2_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(mau_2_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(mau_2_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(mau_2_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(mau_2_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(mau_2_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(mau_2_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(mau_2_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(mau_2_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(mau_2_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(mau_2_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(mau_2_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(mau_2_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(mau_2_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(mau_2_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(mau_2_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(mau_2_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(mau_2_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(mau_2_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(mau_2_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(mau_2_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(mau_2_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(mau_2_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(mau_2_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(mau_2_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(mau_2_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(mau_2_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(mau_2_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(mau_2_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(mau_2_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(mau_2_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(mau_2_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(mau_2_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(mau_2_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(mau_2_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(mau_2_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(mau_2_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(mau_2_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(mau_2_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(mau_2_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(mau_2_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(mau_2_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(mau_2_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(mau_2_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(mau_2_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(mau_2_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(mau_2_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(mau_2_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(mau_2_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(mau_2_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(mau_2_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(mau_2_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(mau_2_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(mau_2_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(mau_2_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(mau_2_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(mau_2_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(mau_2_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(mau_2_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(mau_2_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(mau_2_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(mau_2_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(mau_2_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(mau_2_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(mau_2_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(mau_2_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(mau_2_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(mau_2_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(mau_2_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(mau_2_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(mau_2_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(mau_2_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(mau_2_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(mau_2_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(mau_2_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(mau_2_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(mau_2_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(mau_2_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(mau_2_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(mau_2_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(mau_2_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(mau_2_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(mau_2_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(mau_2_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(mau_2_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(mau_2_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(mau_2_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(mau_2_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(mau_2_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(mau_2_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(mau_2_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(mau_2_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(mau_2_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(mau_2_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(mau_2_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(mau_2_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(mau_2_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(mau_2_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(mau_2_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(mau_2_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(mau_2_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(mau_2_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(mau_2_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(mau_2_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(mau_2_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(mau_2_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(mau_2_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(mau_2_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(mau_2_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(mau_2_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(mau_2_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(mau_2_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(mau_2_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(mau_2_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(mau_2_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(mau_2_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(mau_2_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(mau_2_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(mau_2_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(mau_2_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(mau_2_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(mau_2_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(mau_2_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(mau_2_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(mau_2_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(mau_2_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(mau_2_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(mau_2_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(mau_2_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(mau_2_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(mau_2_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(mau_2_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(mau_2_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(mau_2_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(mau_2_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(mau_2_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(mau_2_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(mau_2_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(mau_2_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(mau_2_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(mau_2_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(mau_2_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(mau_2_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(mau_2_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(mau_2_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(mau_2_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(mau_2_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(mau_2_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(mau_2_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(mau_2_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(mau_2_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(mau_2_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(mau_2_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(mau_2_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(mau_2_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(mau_2_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(mau_2_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(mau_2_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(mau_2_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(mau_2_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(mau_2_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(mau_2_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(mau_2_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(mau_2_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(mau_2_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(mau_2_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(mau_2_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(mau_2_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(mau_2_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(mau_2_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(mau_2_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(mau_2_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(mau_2_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(mau_2_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(mau_2_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(mau_2_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(mau_2_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(mau_2_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_header_0(mau_2_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(mau_2_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(mau_2_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(mau_2_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(mau_2_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(mau_2_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(mau_2_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(mau_2_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(mau_2_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(mau_2_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(mau_2_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(mau_2_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(mau_2_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(mau_2_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(mau_2_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(mau_2_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(mau_2_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(mau_2_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(mau_2_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(mau_2_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(mau_2_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(mau_2_io_pipe_phv_out_is_valid_processor),
    .io_mod_state_id_mod(mau_2_io_mod_state_id_mod),
    .io_mod_state_id(mau_2_io_mod_state_id),
    .io_mod_sram_w_cs(mau_2_io_mod_sram_w_cs),
    .io_mod_sram_w_en(mau_2_io_mod_sram_w_en),
    .io_mod_sram_w_addr(mau_2_io_mod_sram_w_addr),
    .io_mod_sram_w_data(mau_2_io_mod_sram_w_data)
  );
  ParseModule mau_3 ( // @[parser.scala 21:25]
    .clock(mau_3_clock),
    .io_pipe_phv_in_data_0(mau_3_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(mau_3_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(mau_3_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(mau_3_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(mau_3_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(mau_3_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(mau_3_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(mau_3_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(mau_3_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(mau_3_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(mau_3_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(mau_3_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(mau_3_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(mau_3_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(mau_3_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(mau_3_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(mau_3_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(mau_3_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(mau_3_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(mau_3_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(mau_3_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(mau_3_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(mau_3_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(mau_3_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(mau_3_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(mau_3_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(mau_3_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(mau_3_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(mau_3_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(mau_3_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(mau_3_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(mau_3_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(mau_3_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(mau_3_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(mau_3_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(mau_3_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(mau_3_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(mau_3_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(mau_3_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(mau_3_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(mau_3_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(mau_3_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(mau_3_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(mau_3_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(mau_3_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(mau_3_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(mau_3_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(mau_3_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(mau_3_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(mau_3_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(mau_3_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(mau_3_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(mau_3_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(mau_3_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(mau_3_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(mau_3_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(mau_3_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(mau_3_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(mau_3_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(mau_3_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(mau_3_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(mau_3_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(mau_3_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(mau_3_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(mau_3_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(mau_3_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(mau_3_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(mau_3_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(mau_3_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(mau_3_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(mau_3_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(mau_3_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(mau_3_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(mau_3_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(mau_3_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(mau_3_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(mau_3_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(mau_3_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(mau_3_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(mau_3_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(mau_3_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(mau_3_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(mau_3_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(mau_3_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(mau_3_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(mau_3_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(mau_3_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(mau_3_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(mau_3_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(mau_3_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(mau_3_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(mau_3_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(mau_3_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(mau_3_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(mau_3_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(mau_3_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(mau_3_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(mau_3_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(mau_3_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(mau_3_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(mau_3_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(mau_3_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(mau_3_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(mau_3_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(mau_3_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(mau_3_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(mau_3_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(mau_3_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(mau_3_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(mau_3_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(mau_3_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(mau_3_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(mau_3_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(mau_3_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(mau_3_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(mau_3_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(mau_3_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(mau_3_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(mau_3_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(mau_3_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(mau_3_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(mau_3_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(mau_3_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(mau_3_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(mau_3_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(mau_3_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(mau_3_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(mau_3_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(mau_3_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(mau_3_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(mau_3_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(mau_3_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(mau_3_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(mau_3_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(mau_3_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(mau_3_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(mau_3_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(mau_3_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(mau_3_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(mau_3_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(mau_3_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(mau_3_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(mau_3_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(mau_3_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(mau_3_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(mau_3_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(mau_3_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(mau_3_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(mau_3_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(mau_3_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(mau_3_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(mau_3_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(mau_3_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(mau_3_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(mau_3_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(mau_3_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(mau_3_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(mau_3_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(mau_3_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(mau_3_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(mau_3_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(mau_3_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(mau_3_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(mau_3_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(mau_3_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(mau_3_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(mau_3_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(mau_3_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(mau_3_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(mau_3_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(mau_3_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(mau_3_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(mau_3_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(mau_3_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(mau_3_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(mau_3_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(mau_3_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(mau_3_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(mau_3_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(mau_3_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(mau_3_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(mau_3_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(mau_3_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(mau_3_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(mau_3_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(mau_3_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(mau_3_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(mau_3_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(mau_3_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(mau_3_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(mau_3_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(mau_3_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(mau_3_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(mau_3_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(mau_3_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(mau_3_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(mau_3_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(mau_3_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(mau_3_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(mau_3_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(mau_3_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(mau_3_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(mau_3_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(mau_3_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(mau_3_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(mau_3_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(mau_3_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(mau_3_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(mau_3_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(mau_3_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(mau_3_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(mau_3_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(mau_3_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(mau_3_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(mau_3_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(mau_3_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(mau_3_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(mau_3_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(mau_3_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(mau_3_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(mau_3_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(mau_3_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(mau_3_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(mau_3_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(mau_3_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(mau_3_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(mau_3_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(mau_3_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(mau_3_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(mau_3_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(mau_3_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(mau_3_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(mau_3_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(mau_3_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(mau_3_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(mau_3_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(mau_3_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(mau_3_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(mau_3_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(mau_3_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(mau_3_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(mau_3_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(mau_3_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(mau_3_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(mau_3_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(mau_3_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(mau_3_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(mau_3_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(mau_3_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(mau_3_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(mau_3_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(mau_3_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(mau_3_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(mau_3_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(mau_3_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(mau_3_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_header_0(mau_3_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(mau_3_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(mau_3_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(mau_3_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(mau_3_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(mau_3_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(mau_3_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(mau_3_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(mau_3_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(mau_3_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(mau_3_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(mau_3_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(mau_3_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(mau_3_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(mau_3_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(mau_3_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(mau_3_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(mau_3_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(mau_3_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(mau_3_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(mau_3_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(mau_3_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(mau_3_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(mau_3_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(mau_3_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(mau_3_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(mau_3_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(mau_3_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(mau_3_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(mau_3_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(mau_3_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(mau_3_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(mau_3_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(mau_3_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(mau_3_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(mau_3_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(mau_3_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(mau_3_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(mau_3_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(mau_3_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(mau_3_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(mau_3_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(mau_3_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(mau_3_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(mau_3_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(mau_3_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(mau_3_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(mau_3_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(mau_3_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(mau_3_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(mau_3_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(mau_3_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(mau_3_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(mau_3_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(mau_3_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(mau_3_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(mau_3_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(mau_3_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(mau_3_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(mau_3_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(mau_3_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(mau_3_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(mau_3_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(mau_3_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(mau_3_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(mau_3_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(mau_3_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(mau_3_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(mau_3_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(mau_3_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(mau_3_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(mau_3_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(mau_3_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(mau_3_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(mau_3_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(mau_3_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(mau_3_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(mau_3_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(mau_3_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(mau_3_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(mau_3_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(mau_3_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(mau_3_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(mau_3_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(mau_3_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(mau_3_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(mau_3_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(mau_3_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(mau_3_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(mau_3_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(mau_3_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(mau_3_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(mau_3_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(mau_3_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(mau_3_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(mau_3_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(mau_3_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(mau_3_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(mau_3_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(mau_3_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(mau_3_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(mau_3_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(mau_3_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(mau_3_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(mau_3_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(mau_3_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(mau_3_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(mau_3_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(mau_3_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(mau_3_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(mau_3_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(mau_3_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(mau_3_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(mau_3_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(mau_3_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(mau_3_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(mau_3_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(mau_3_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(mau_3_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(mau_3_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(mau_3_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(mau_3_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(mau_3_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(mau_3_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(mau_3_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(mau_3_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(mau_3_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(mau_3_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(mau_3_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(mau_3_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(mau_3_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(mau_3_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(mau_3_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(mau_3_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(mau_3_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(mau_3_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(mau_3_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(mau_3_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(mau_3_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(mau_3_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(mau_3_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(mau_3_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(mau_3_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(mau_3_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(mau_3_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(mau_3_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(mau_3_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(mau_3_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(mau_3_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(mau_3_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(mau_3_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(mau_3_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(mau_3_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(mau_3_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(mau_3_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(mau_3_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(mau_3_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(mau_3_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(mau_3_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(mau_3_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(mau_3_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(mau_3_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(mau_3_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(mau_3_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(mau_3_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(mau_3_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(mau_3_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(mau_3_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(mau_3_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(mau_3_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(mau_3_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(mau_3_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(mau_3_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(mau_3_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(mau_3_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(mau_3_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(mau_3_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(mau_3_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(mau_3_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(mau_3_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(mau_3_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(mau_3_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(mau_3_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(mau_3_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(mau_3_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(mau_3_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(mau_3_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(mau_3_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(mau_3_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(mau_3_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(mau_3_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(mau_3_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(mau_3_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(mau_3_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(mau_3_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(mau_3_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(mau_3_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(mau_3_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(mau_3_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(mau_3_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(mau_3_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(mau_3_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(mau_3_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(mau_3_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(mau_3_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(mau_3_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(mau_3_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(mau_3_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(mau_3_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(mau_3_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(mau_3_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(mau_3_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(mau_3_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(mau_3_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(mau_3_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(mau_3_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(mau_3_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(mau_3_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(mau_3_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(mau_3_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(mau_3_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(mau_3_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(mau_3_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(mau_3_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(mau_3_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(mau_3_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(mau_3_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(mau_3_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(mau_3_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(mau_3_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(mau_3_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(mau_3_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(mau_3_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(mau_3_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(mau_3_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(mau_3_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(mau_3_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(mau_3_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(mau_3_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(mau_3_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(mau_3_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(mau_3_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(mau_3_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(mau_3_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(mau_3_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(mau_3_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(mau_3_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(mau_3_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(mau_3_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(mau_3_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(mau_3_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(mau_3_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(mau_3_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(mau_3_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(mau_3_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(mau_3_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(mau_3_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(mau_3_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(mau_3_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(mau_3_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(mau_3_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(mau_3_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(mau_3_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(mau_3_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(mau_3_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(mau_3_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(mau_3_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(mau_3_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(mau_3_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(mau_3_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(mau_3_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(mau_3_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(mau_3_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(mau_3_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(mau_3_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(mau_3_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(mau_3_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(mau_3_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_header_0(mau_3_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(mau_3_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(mau_3_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(mau_3_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(mau_3_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(mau_3_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(mau_3_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(mau_3_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(mau_3_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(mau_3_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(mau_3_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(mau_3_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(mau_3_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(mau_3_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(mau_3_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(mau_3_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(mau_3_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(mau_3_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(mau_3_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(mau_3_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(mau_3_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(mau_3_io_pipe_phv_out_is_valid_processor),
    .io_mod_state_id_mod(mau_3_io_mod_state_id_mod),
    .io_mod_state_id(mau_3_io_mod_state_id),
    .io_mod_sram_w_cs(mau_3_io_mod_sram_w_cs),
    .io_mod_sram_w_en(mau_3_io_mod_sram_w_en),
    .io_mod_sram_w_addr(mau_3_io_mod_sram_w_addr),
    .io_mod_sram_w_data(mau_3_io_mod_sram_w_data)
  );
  assign io_pipe_phv_out_data_0 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_0 : _GEN_300; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_1 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_1 : _GEN_301; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_2 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_2 : _GEN_302; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_3 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_3 : _GEN_303; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_4 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_4 : _GEN_304; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_5 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_5 : _GEN_305; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_6 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_6 : _GEN_306; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_7 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_7 : _GEN_307; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_8 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_8 : _GEN_308; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_9 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_9 : _GEN_309; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_10 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_10 : _GEN_310; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_11 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_11 : _GEN_311; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_12 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_12 : _GEN_312; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_13 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_13 : _GEN_313; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_14 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_14 : _GEN_314; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_15 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_15 : _GEN_315; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_16 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_16 : _GEN_316; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_17 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_17 : _GEN_317; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_18 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_18 : _GEN_318; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_19 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_19 : _GEN_319; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_20 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_20 : _GEN_320; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_21 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_21 : _GEN_321; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_22 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_22 : _GEN_322; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_23 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_23 : _GEN_323; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_24 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_24 : _GEN_324; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_25 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_25 : _GEN_325; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_26 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_26 : _GEN_326; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_27 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_27 : _GEN_327; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_28 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_28 : _GEN_328; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_29 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_29 : _GEN_329; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_30 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_30 : _GEN_330; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_31 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_31 : _GEN_331; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_32 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_32 : _GEN_332; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_33 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_33 : _GEN_333; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_34 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_34 : _GEN_334; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_35 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_35 : _GEN_335; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_36 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_36 : _GEN_336; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_37 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_37 : _GEN_337; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_38 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_38 : _GEN_338; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_39 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_39 : _GEN_339; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_40 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_40 : _GEN_340; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_41 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_41 : _GEN_341; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_42 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_42 : _GEN_342; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_43 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_43 : _GEN_343; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_44 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_44 : _GEN_344; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_45 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_45 : _GEN_345; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_46 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_46 : _GEN_346; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_47 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_47 : _GEN_347; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_48 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_48 : _GEN_348; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_49 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_49 : _GEN_349; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_50 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_50 : _GEN_350; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_51 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_51 : _GEN_351; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_52 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_52 : _GEN_352; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_53 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_53 : _GEN_353; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_54 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_54 : _GEN_354; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_55 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_55 : _GEN_355; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_56 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_56 : _GEN_356; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_57 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_57 : _GEN_357; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_58 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_58 : _GEN_358; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_59 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_59 : _GEN_359; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_60 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_60 : _GEN_360; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_61 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_61 : _GEN_361; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_62 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_62 : _GEN_362; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_63 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_63 : _GEN_363; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_64 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_64 : _GEN_364; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_65 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_65 : _GEN_365; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_66 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_66 : _GEN_366; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_67 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_67 : _GEN_367; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_68 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_68 : _GEN_368; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_69 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_69 : _GEN_369; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_70 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_70 : _GEN_370; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_71 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_71 : _GEN_371; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_72 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_72 : _GEN_372; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_73 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_73 : _GEN_373; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_74 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_74 : _GEN_374; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_75 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_75 : _GEN_375; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_76 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_76 : _GEN_376; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_77 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_77 : _GEN_377; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_78 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_78 : _GEN_378; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_79 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_79 : _GEN_379; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_80 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_80 : _GEN_380; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_81 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_81 : _GEN_381; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_82 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_82 : _GEN_382; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_83 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_83 : _GEN_383; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_84 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_84 : _GEN_384; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_85 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_85 : _GEN_385; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_86 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_86 : _GEN_386; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_87 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_87 : _GEN_387; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_88 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_88 : _GEN_388; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_89 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_89 : _GEN_389; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_90 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_90 : _GEN_390; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_91 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_91 : _GEN_391; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_92 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_92 : _GEN_392; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_93 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_93 : _GEN_393; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_94 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_94 : _GEN_394; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_95 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_95 : _GEN_395; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_96 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_96 : _GEN_396; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_97 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_97 : _GEN_397; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_98 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_98 : _GEN_398; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_99 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_99 : _GEN_399; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_100 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_100 : _GEN_400; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_101 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_101 : _GEN_401; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_102 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_102 : _GEN_402; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_103 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_103 : _GEN_403; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_104 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_104 : _GEN_404; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_105 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_105 : _GEN_405; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_106 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_106 : _GEN_406; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_107 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_107 : _GEN_407; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_108 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_108 : _GEN_408; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_109 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_109 : _GEN_409; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_110 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_110 : _GEN_410; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_111 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_111 : _GEN_411; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_112 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_112 : _GEN_412; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_113 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_113 : _GEN_413; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_114 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_114 : _GEN_414; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_115 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_115 : _GEN_415; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_116 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_116 : _GEN_416; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_117 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_117 : _GEN_417; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_118 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_118 : _GEN_418; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_119 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_119 : _GEN_419; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_120 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_120 : _GEN_420; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_121 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_121 : _GEN_421; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_122 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_122 : _GEN_422; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_123 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_123 : _GEN_423; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_124 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_124 : _GEN_424; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_125 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_125 : _GEN_425; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_126 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_126 : _GEN_426; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_127 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_127 : _GEN_427; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_128 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_128 : _GEN_428; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_129 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_129 : _GEN_429; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_130 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_130 : _GEN_430; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_131 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_131 : _GEN_431; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_132 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_132 : _GEN_432; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_133 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_133 : _GEN_433; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_134 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_134 : _GEN_434; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_135 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_135 : _GEN_435; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_136 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_136 : _GEN_436; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_137 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_137 : _GEN_437; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_138 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_138 : _GEN_438; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_139 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_139 : _GEN_439; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_140 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_140 : _GEN_440; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_141 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_141 : _GEN_441; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_142 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_142 : _GEN_442; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_143 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_143 : _GEN_443; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_144 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_144 : _GEN_444; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_145 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_145 : _GEN_445; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_146 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_146 : _GEN_446; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_147 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_147 : _GEN_447; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_148 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_148 : _GEN_448; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_149 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_149 : _GEN_449; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_150 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_150 : _GEN_450; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_151 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_151 : _GEN_451; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_152 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_152 : _GEN_452; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_153 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_153 : _GEN_453; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_154 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_154 : _GEN_454; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_155 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_155 : _GEN_455; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_156 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_156 : _GEN_456; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_157 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_157 : _GEN_457; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_158 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_158 : _GEN_458; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_159 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_159 : _GEN_459; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_160 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_160 : _GEN_460; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_161 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_161 : _GEN_461; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_162 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_162 : _GEN_462; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_163 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_163 : _GEN_463; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_164 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_164 : _GEN_464; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_165 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_165 : _GEN_465; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_166 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_166 : _GEN_466; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_167 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_167 : _GEN_467; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_168 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_168 : _GEN_468; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_169 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_169 : _GEN_469; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_170 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_170 : _GEN_470; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_171 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_171 : _GEN_471; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_172 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_172 : _GEN_472; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_173 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_173 : _GEN_473; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_174 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_174 : _GEN_474; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_175 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_175 : _GEN_475; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_176 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_176 : _GEN_476; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_177 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_177 : _GEN_477; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_178 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_178 : _GEN_478; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_179 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_179 : _GEN_479; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_180 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_180 : _GEN_480; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_181 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_181 : _GEN_481; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_182 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_182 : _GEN_482; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_183 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_183 : _GEN_483; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_184 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_184 : _GEN_484; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_185 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_185 : _GEN_485; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_186 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_186 : _GEN_486; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_187 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_187 : _GEN_487; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_188 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_188 : _GEN_488; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_189 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_189 : _GEN_489; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_190 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_190 : _GEN_490; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_191 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_191 : _GEN_491; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_192 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_192 : _GEN_492; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_193 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_193 : _GEN_493; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_194 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_194 : _GEN_494; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_195 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_195 : _GEN_495; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_196 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_196 : _GEN_496; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_197 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_197 : _GEN_497; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_198 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_198 : _GEN_498; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_199 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_199 : _GEN_499; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_200 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_200 : _GEN_500; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_201 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_201 : _GEN_501; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_202 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_202 : _GEN_502; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_203 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_203 : _GEN_503; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_204 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_204 : _GEN_504; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_205 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_205 : _GEN_505; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_206 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_206 : _GEN_506; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_207 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_207 : _GEN_507; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_208 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_208 : _GEN_508; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_209 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_209 : _GEN_509; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_210 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_210 : _GEN_510; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_211 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_211 : _GEN_511; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_212 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_212 : _GEN_512; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_213 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_213 : _GEN_513; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_214 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_214 : _GEN_514; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_215 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_215 : _GEN_515; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_216 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_216 : _GEN_516; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_217 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_217 : _GEN_517; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_218 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_218 : _GEN_518; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_219 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_219 : _GEN_519; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_220 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_220 : _GEN_520; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_221 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_221 : _GEN_521; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_222 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_222 : _GEN_522; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_223 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_223 : _GEN_523; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_224 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_224 : _GEN_524; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_225 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_225 : _GEN_525; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_226 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_226 : _GEN_526; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_227 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_227 : _GEN_527; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_228 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_228 : _GEN_528; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_229 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_229 : _GEN_529; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_230 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_230 : _GEN_530; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_231 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_231 : _GEN_531; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_232 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_232 : _GEN_532; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_233 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_233 : _GEN_533; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_234 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_234 : _GEN_534; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_235 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_235 : _GEN_535; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_236 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_236 : _GEN_536; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_237 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_237 : _GEN_537; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_238 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_238 : _GEN_538; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_239 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_239 : _GEN_539; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_240 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_240 : _GEN_540; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_241 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_241 : _GEN_541; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_242 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_242 : _GEN_542; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_243 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_243 : _GEN_543; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_244 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_244 : _GEN_544; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_245 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_245 : _GEN_545; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_246 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_246 : _GEN_546; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_247 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_247 : _GEN_547; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_248 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_248 : _GEN_548; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_249 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_249 : _GEN_549; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_250 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_250 : _GEN_550; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_251 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_251 : _GEN_551; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_252 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_252 : _GEN_552; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_253 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_253 : _GEN_553; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_254 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_254 : _GEN_554; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_255 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_255 : _GEN_555; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_header_0 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_header_0 : _GEN_284; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_header_1 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_header_1 : _GEN_285; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_header_2 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_header_2 : _GEN_286; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_header_3 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_header_3 : _GEN_287; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_header_4 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_header_4 : _GEN_288; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_header_5 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_header_5 : _GEN_289; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_header_6 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_header_6 : _GEN_290; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_header_7 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_header_7 : _GEN_291; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_header_8 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_header_8 : _GEN_292; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_header_9 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_header_9 : _GEN_293; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_header_10 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_header_10 : _GEN_294; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_header_11 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_header_11 : _GEN_295; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_header_12 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_header_12 : _GEN_296; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_header_13 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_header_13 : _GEN_297; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_header_14 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_header_14 : _GEN_298; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_header_15 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_header_15 : _GEN_299; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_parse_current_state = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_parse_current_state :
    _GEN_283; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_parse_current_offset = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_parse_current_offset :
    _GEN_282; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_parse_transition_field = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_parse_transition_field :
    _GEN_281; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_next_processor_id = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_next_processor_id : _GEN_280; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_next_config_id = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_next_config_id : _GEN_279; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_is_valid_processor = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_is_valid_processor : _GEN_278; // @[parser.scala 33:62 parser.scala 34:35]
  assign mau_0_clock = clock;
  assign mau_0_io_pipe_phv_in_data_0 = io_pipe_phv_in_data_0; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_1 = io_pipe_phv_in_data_1; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_2 = io_pipe_phv_in_data_2; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_3 = io_pipe_phv_in_data_3; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_4 = io_pipe_phv_in_data_4; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_5 = io_pipe_phv_in_data_5; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_6 = io_pipe_phv_in_data_6; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_7 = io_pipe_phv_in_data_7; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_8 = io_pipe_phv_in_data_8; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_9 = io_pipe_phv_in_data_9; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_10 = io_pipe_phv_in_data_10; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_11 = io_pipe_phv_in_data_11; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_12 = io_pipe_phv_in_data_12; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_13 = io_pipe_phv_in_data_13; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_14 = io_pipe_phv_in_data_14; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_15 = io_pipe_phv_in_data_15; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_16 = io_pipe_phv_in_data_16; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_17 = io_pipe_phv_in_data_17; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_18 = io_pipe_phv_in_data_18; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_19 = io_pipe_phv_in_data_19; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_20 = io_pipe_phv_in_data_20; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_21 = io_pipe_phv_in_data_21; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_22 = io_pipe_phv_in_data_22; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_23 = io_pipe_phv_in_data_23; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_24 = io_pipe_phv_in_data_24; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_25 = io_pipe_phv_in_data_25; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_26 = io_pipe_phv_in_data_26; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_27 = io_pipe_phv_in_data_27; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_28 = io_pipe_phv_in_data_28; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_29 = io_pipe_phv_in_data_29; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_30 = io_pipe_phv_in_data_30; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_31 = io_pipe_phv_in_data_31; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_32 = io_pipe_phv_in_data_32; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_33 = io_pipe_phv_in_data_33; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_34 = io_pipe_phv_in_data_34; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_35 = io_pipe_phv_in_data_35; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_36 = io_pipe_phv_in_data_36; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_37 = io_pipe_phv_in_data_37; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_38 = io_pipe_phv_in_data_38; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_39 = io_pipe_phv_in_data_39; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_40 = io_pipe_phv_in_data_40; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_41 = io_pipe_phv_in_data_41; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_42 = io_pipe_phv_in_data_42; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_43 = io_pipe_phv_in_data_43; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_44 = io_pipe_phv_in_data_44; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_45 = io_pipe_phv_in_data_45; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_46 = io_pipe_phv_in_data_46; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_47 = io_pipe_phv_in_data_47; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_48 = io_pipe_phv_in_data_48; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_49 = io_pipe_phv_in_data_49; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_50 = io_pipe_phv_in_data_50; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_51 = io_pipe_phv_in_data_51; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_52 = io_pipe_phv_in_data_52; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_53 = io_pipe_phv_in_data_53; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_54 = io_pipe_phv_in_data_54; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_55 = io_pipe_phv_in_data_55; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_56 = io_pipe_phv_in_data_56; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_57 = io_pipe_phv_in_data_57; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_58 = io_pipe_phv_in_data_58; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_59 = io_pipe_phv_in_data_59; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_60 = io_pipe_phv_in_data_60; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_61 = io_pipe_phv_in_data_61; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_62 = io_pipe_phv_in_data_62; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_63 = io_pipe_phv_in_data_63; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_64 = io_pipe_phv_in_data_64; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_65 = io_pipe_phv_in_data_65; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_66 = io_pipe_phv_in_data_66; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_67 = io_pipe_phv_in_data_67; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_68 = io_pipe_phv_in_data_68; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_69 = io_pipe_phv_in_data_69; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_70 = io_pipe_phv_in_data_70; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_71 = io_pipe_phv_in_data_71; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_72 = io_pipe_phv_in_data_72; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_73 = io_pipe_phv_in_data_73; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_74 = io_pipe_phv_in_data_74; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_75 = io_pipe_phv_in_data_75; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_76 = io_pipe_phv_in_data_76; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_77 = io_pipe_phv_in_data_77; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_78 = io_pipe_phv_in_data_78; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_79 = io_pipe_phv_in_data_79; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_80 = io_pipe_phv_in_data_80; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_81 = io_pipe_phv_in_data_81; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_82 = io_pipe_phv_in_data_82; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_83 = io_pipe_phv_in_data_83; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_84 = io_pipe_phv_in_data_84; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_85 = io_pipe_phv_in_data_85; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_86 = io_pipe_phv_in_data_86; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_87 = io_pipe_phv_in_data_87; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_88 = io_pipe_phv_in_data_88; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_89 = io_pipe_phv_in_data_89; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_90 = io_pipe_phv_in_data_90; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_91 = io_pipe_phv_in_data_91; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_92 = io_pipe_phv_in_data_92; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_93 = io_pipe_phv_in_data_93; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_94 = io_pipe_phv_in_data_94; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_95 = io_pipe_phv_in_data_95; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_96 = io_pipe_phv_in_data_96; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_97 = io_pipe_phv_in_data_97; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_98 = io_pipe_phv_in_data_98; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_99 = io_pipe_phv_in_data_99; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_100 = io_pipe_phv_in_data_100; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_101 = io_pipe_phv_in_data_101; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_102 = io_pipe_phv_in_data_102; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_103 = io_pipe_phv_in_data_103; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_104 = io_pipe_phv_in_data_104; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_105 = io_pipe_phv_in_data_105; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_106 = io_pipe_phv_in_data_106; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_107 = io_pipe_phv_in_data_107; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_108 = io_pipe_phv_in_data_108; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_109 = io_pipe_phv_in_data_109; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_110 = io_pipe_phv_in_data_110; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_111 = io_pipe_phv_in_data_111; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_112 = io_pipe_phv_in_data_112; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_113 = io_pipe_phv_in_data_113; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_114 = io_pipe_phv_in_data_114; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_115 = io_pipe_phv_in_data_115; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_116 = io_pipe_phv_in_data_116; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_117 = io_pipe_phv_in_data_117; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_118 = io_pipe_phv_in_data_118; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_119 = io_pipe_phv_in_data_119; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_120 = io_pipe_phv_in_data_120; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_121 = io_pipe_phv_in_data_121; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_122 = io_pipe_phv_in_data_122; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_123 = io_pipe_phv_in_data_123; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_124 = io_pipe_phv_in_data_124; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_125 = io_pipe_phv_in_data_125; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_126 = io_pipe_phv_in_data_126; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_127 = io_pipe_phv_in_data_127; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_128 = io_pipe_phv_in_data_128; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_129 = io_pipe_phv_in_data_129; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_130 = io_pipe_phv_in_data_130; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_131 = io_pipe_phv_in_data_131; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_132 = io_pipe_phv_in_data_132; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_133 = io_pipe_phv_in_data_133; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_134 = io_pipe_phv_in_data_134; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_135 = io_pipe_phv_in_data_135; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_136 = io_pipe_phv_in_data_136; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_137 = io_pipe_phv_in_data_137; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_138 = io_pipe_phv_in_data_138; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_139 = io_pipe_phv_in_data_139; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_140 = io_pipe_phv_in_data_140; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_141 = io_pipe_phv_in_data_141; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_142 = io_pipe_phv_in_data_142; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_143 = io_pipe_phv_in_data_143; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_144 = io_pipe_phv_in_data_144; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_145 = io_pipe_phv_in_data_145; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_146 = io_pipe_phv_in_data_146; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_147 = io_pipe_phv_in_data_147; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_148 = io_pipe_phv_in_data_148; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_149 = io_pipe_phv_in_data_149; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_150 = io_pipe_phv_in_data_150; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_151 = io_pipe_phv_in_data_151; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_152 = io_pipe_phv_in_data_152; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_153 = io_pipe_phv_in_data_153; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_154 = io_pipe_phv_in_data_154; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_155 = io_pipe_phv_in_data_155; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_156 = io_pipe_phv_in_data_156; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_157 = io_pipe_phv_in_data_157; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_158 = io_pipe_phv_in_data_158; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_159 = io_pipe_phv_in_data_159; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_160 = io_pipe_phv_in_data_160; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_161 = io_pipe_phv_in_data_161; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_162 = io_pipe_phv_in_data_162; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_163 = io_pipe_phv_in_data_163; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_164 = io_pipe_phv_in_data_164; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_165 = io_pipe_phv_in_data_165; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_166 = io_pipe_phv_in_data_166; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_167 = io_pipe_phv_in_data_167; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_168 = io_pipe_phv_in_data_168; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_169 = io_pipe_phv_in_data_169; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_170 = io_pipe_phv_in_data_170; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_171 = io_pipe_phv_in_data_171; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_172 = io_pipe_phv_in_data_172; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_173 = io_pipe_phv_in_data_173; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_174 = io_pipe_phv_in_data_174; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_175 = io_pipe_phv_in_data_175; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_176 = io_pipe_phv_in_data_176; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_177 = io_pipe_phv_in_data_177; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_178 = io_pipe_phv_in_data_178; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_179 = io_pipe_phv_in_data_179; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_180 = io_pipe_phv_in_data_180; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_181 = io_pipe_phv_in_data_181; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_182 = io_pipe_phv_in_data_182; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_183 = io_pipe_phv_in_data_183; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_184 = io_pipe_phv_in_data_184; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_185 = io_pipe_phv_in_data_185; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_186 = io_pipe_phv_in_data_186; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_187 = io_pipe_phv_in_data_187; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_188 = io_pipe_phv_in_data_188; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_189 = io_pipe_phv_in_data_189; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_190 = io_pipe_phv_in_data_190; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_191 = io_pipe_phv_in_data_191; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_192 = io_pipe_phv_in_data_192; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_193 = io_pipe_phv_in_data_193; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_194 = io_pipe_phv_in_data_194; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_195 = io_pipe_phv_in_data_195; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_196 = io_pipe_phv_in_data_196; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_197 = io_pipe_phv_in_data_197; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_198 = io_pipe_phv_in_data_198; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_199 = io_pipe_phv_in_data_199; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_200 = io_pipe_phv_in_data_200; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_201 = io_pipe_phv_in_data_201; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_202 = io_pipe_phv_in_data_202; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_203 = io_pipe_phv_in_data_203; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_204 = io_pipe_phv_in_data_204; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_205 = io_pipe_phv_in_data_205; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_206 = io_pipe_phv_in_data_206; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_207 = io_pipe_phv_in_data_207; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_208 = io_pipe_phv_in_data_208; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_209 = io_pipe_phv_in_data_209; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_210 = io_pipe_phv_in_data_210; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_211 = io_pipe_phv_in_data_211; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_212 = io_pipe_phv_in_data_212; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_213 = io_pipe_phv_in_data_213; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_214 = io_pipe_phv_in_data_214; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_215 = io_pipe_phv_in_data_215; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_216 = io_pipe_phv_in_data_216; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_217 = io_pipe_phv_in_data_217; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_218 = io_pipe_phv_in_data_218; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_219 = io_pipe_phv_in_data_219; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_220 = io_pipe_phv_in_data_220; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_221 = io_pipe_phv_in_data_221; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_222 = io_pipe_phv_in_data_222; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_223 = io_pipe_phv_in_data_223; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_224 = io_pipe_phv_in_data_224; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_225 = io_pipe_phv_in_data_225; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_226 = io_pipe_phv_in_data_226; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_227 = io_pipe_phv_in_data_227; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_228 = io_pipe_phv_in_data_228; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_229 = io_pipe_phv_in_data_229; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_230 = io_pipe_phv_in_data_230; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_231 = io_pipe_phv_in_data_231; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_232 = io_pipe_phv_in_data_232; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_233 = io_pipe_phv_in_data_233; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_234 = io_pipe_phv_in_data_234; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_235 = io_pipe_phv_in_data_235; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_236 = io_pipe_phv_in_data_236; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_237 = io_pipe_phv_in_data_237; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_238 = io_pipe_phv_in_data_238; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_239 = io_pipe_phv_in_data_239; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_240 = io_pipe_phv_in_data_240; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_241 = io_pipe_phv_in_data_241; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_242 = io_pipe_phv_in_data_242; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_243 = io_pipe_phv_in_data_243; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_244 = io_pipe_phv_in_data_244; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_245 = io_pipe_phv_in_data_245; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_246 = io_pipe_phv_in_data_246; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_247 = io_pipe_phv_in_data_247; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_248 = io_pipe_phv_in_data_248; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_249 = io_pipe_phv_in_data_249; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_250 = io_pipe_phv_in_data_250; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_251 = io_pipe_phv_in_data_251; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_252 = io_pipe_phv_in_data_252; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_253 = io_pipe_phv_in_data_253; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_254 = io_pipe_phv_in_data_254; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_255 = io_pipe_phv_in_data_255; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_header_0 = io_pipe_phv_in_header_0; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_header_1 = io_pipe_phv_in_header_1; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_header_2 = io_pipe_phv_in_header_2; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_header_3 = io_pipe_phv_in_header_3; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_header_4 = io_pipe_phv_in_header_4; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_header_5 = io_pipe_phv_in_header_5; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_header_6 = io_pipe_phv_in_header_6; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_header_7 = io_pipe_phv_in_header_7; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_header_8 = io_pipe_phv_in_header_8; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_header_9 = io_pipe_phv_in_header_9; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_header_10 = io_pipe_phv_in_header_10; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_header_11 = io_pipe_phv_in_header_11; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_header_12 = io_pipe_phv_in_header_12; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_header_13 = io_pipe_phv_in_header_13; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_header_14 = io_pipe_phv_in_header_14; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_header_15 = io_pipe_phv_in_header_15; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_parse_current_state = io_pipe_phv_in_parse_current_state; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_parse_current_offset = io_pipe_phv_in_parse_current_offset; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_parse_transition_field = io_pipe_phv_in_parse_transition_field; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_next_processor_id = io_pipe_phv_in_next_processor_id; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_next_config_id = io_pipe_phv_in_next_config_id; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_is_valid_processor = io_pipe_phv_in_is_valid_processor; // @[parser.scala 30:35]
  assign mau_0_io_mod_state_id_mod = io_mod_en ? io_mod_module_mod_state_id_mod & mod_j : io_mod_module_mod_state_id_mod
    ; // @[parser.scala 41:22 parser.scala 48:40 parser.scala 37:23]
  assign mau_0_io_mod_state_id = io_mod_module_mod_state_id; // @[parser.scala 37:23]
  assign mau_0_io_mod_sram_w_cs = io_mod_module_mod_sram_w_cs; // @[parser.scala 37:23]
  assign mau_0_io_mod_sram_w_en = io_mod_en ? io_mod_module_mod_sram_w_en & mod_j : io_mod_module_mod_sram_w_en; // @[parser.scala 41:22 parser.scala 47:40 parser.scala 37:23]
  assign mau_0_io_mod_sram_w_addr = io_mod_module_mod_sram_w_addr; // @[parser.scala 37:23]
  assign mau_0_io_mod_sram_w_data = io_mod_module_mod_sram_w_data; // @[parser.scala 37:23]
  assign mau_1_clock = clock;
  assign mau_1_io_pipe_phv_in_data_0 = mau_0_io_pipe_phv_out_data_0; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_1 = mau_0_io_pipe_phv_out_data_1; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_2 = mau_0_io_pipe_phv_out_data_2; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_3 = mau_0_io_pipe_phv_out_data_3; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_4 = mau_0_io_pipe_phv_out_data_4; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_5 = mau_0_io_pipe_phv_out_data_5; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_6 = mau_0_io_pipe_phv_out_data_6; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_7 = mau_0_io_pipe_phv_out_data_7; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_8 = mau_0_io_pipe_phv_out_data_8; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_9 = mau_0_io_pipe_phv_out_data_9; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_10 = mau_0_io_pipe_phv_out_data_10; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_11 = mau_0_io_pipe_phv_out_data_11; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_12 = mau_0_io_pipe_phv_out_data_12; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_13 = mau_0_io_pipe_phv_out_data_13; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_14 = mau_0_io_pipe_phv_out_data_14; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_15 = mau_0_io_pipe_phv_out_data_15; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_16 = mau_0_io_pipe_phv_out_data_16; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_17 = mau_0_io_pipe_phv_out_data_17; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_18 = mau_0_io_pipe_phv_out_data_18; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_19 = mau_0_io_pipe_phv_out_data_19; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_20 = mau_0_io_pipe_phv_out_data_20; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_21 = mau_0_io_pipe_phv_out_data_21; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_22 = mau_0_io_pipe_phv_out_data_22; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_23 = mau_0_io_pipe_phv_out_data_23; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_24 = mau_0_io_pipe_phv_out_data_24; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_25 = mau_0_io_pipe_phv_out_data_25; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_26 = mau_0_io_pipe_phv_out_data_26; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_27 = mau_0_io_pipe_phv_out_data_27; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_28 = mau_0_io_pipe_phv_out_data_28; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_29 = mau_0_io_pipe_phv_out_data_29; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_30 = mau_0_io_pipe_phv_out_data_30; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_31 = mau_0_io_pipe_phv_out_data_31; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_32 = mau_0_io_pipe_phv_out_data_32; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_33 = mau_0_io_pipe_phv_out_data_33; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_34 = mau_0_io_pipe_phv_out_data_34; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_35 = mau_0_io_pipe_phv_out_data_35; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_36 = mau_0_io_pipe_phv_out_data_36; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_37 = mau_0_io_pipe_phv_out_data_37; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_38 = mau_0_io_pipe_phv_out_data_38; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_39 = mau_0_io_pipe_phv_out_data_39; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_40 = mau_0_io_pipe_phv_out_data_40; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_41 = mau_0_io_pipe_phv_out_data_41; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_42 = mau_0_io_pipe_phv_out_data_42; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_43 = mau_0_io_pipe_phv_out_data_43; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_44 = mau_0_io_pipe_phv_out_data_44; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_45 = mau_0_io_pipe_phv_out_data_45; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_46 = mau_0_io_pipe_phv_out_data_46; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_47 = mau_0_io_pipe_phv_out_data_47; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_48 = mau_0_io_pipe_phv_out_data_48; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_49 = mau_0_io_pipe_phv_out_data_49; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_50 = mau_0_io_pipe_phv_out_data_50; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_51 = mau_0_io_pipe_phv_out_data_51; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_52 = mau_0_io_pipe_phv_out_data_52; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_53 = mau_0_io_pipe_phv_out_data_53; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_54 = mau_0_io_pipe_phv_out_data_54; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_55 = mau_0_io_pipe_phv_out_data_55; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_56 = mau_0_io_pipe_phv_out_data_56; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_57 = mau_0_io_pipe_phv_out_data_57; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_58 = mau_0_io_pipe_phv_out_data_58; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_59 = mau_0_io_pipe_phv_out_data_59; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_60 = mau_0_io_pipe_phv_out_data_60; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_61 = mau_0_io_pipe_phv_out_data_61; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_62 = mau_0_io_pipe_phv_out_data_62; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_63 = mau_0_io_pipe_phv_out_data_63; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_64 = mau_0_io_pipe_phv_out_data_64; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_65 = mau_0_io_pipe_phv_out_data_65; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_66 = mau_0_io_pipe_phv_out_data_66; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_67 = mau_0_io_pipe_phv_out_data_67; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_68 = mau_0_io_pipe_phv_out_data_68; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_69 = mau_0_io_pipe_phv_out_data_69; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_70 = mau_0_io_pipe_phv_out_data_70; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_71 = mau_0_io_pipe_phv_out_data_71; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_72 = mau_0_io_pipe_phv_out_data_72; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_73 = mau_0_io_pipe_phv_out_data_73; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_74 = mau_0_io_pipe_phv_out_data_74; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_75 = mau_0_io_pipe_phv_out_data_75; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_76 = mau_0_io_pipe_phv_out_data_76; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_77 = mau_0_io_pipe_phv_out_data_77; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_78 = mau_0_io_pipe_phv_out_data_78; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_79 = mau_0_io_pipe_phv_out_data_79; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_80 = mau_0_io_pipe_phv_out_data_80; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_81 = mau_0_io_pipe_phv_out_data_81; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_82 = mau_0_io_pipe_phv_out_data_82; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_83 = mau_0_io_pipe_phv_out_data_83; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_84 = mau_0_io_pipe_phv_out_data_84; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_85 = mau_0_io_pipe_phv_out_data_85; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_86 = mau_0_io_pipe_phv_out_data_86; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_87 = mau_0_io_pipe_phv_out_data_87; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_88 = mau_0_io_pipe_phv_out_data_88; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_89 = mau_0_io_pipe_phv_out_data_89; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_90 = mau_0_io_pipe_phv_out_data_90; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_91 = mau_0_io_pipe_phv_out_data_91; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_92 = mau_0_io_pipe_phv_out_data_92; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_93 = mau_0_io_pipe_phv_out_data_93; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_94 = mau_0_io_pipe_phv_out_data_94; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_95 = mau_0_io_pipe_phv_out_data_95; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_96 = mau_0_io_pipe_phv_out_data_96; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_97 = mau_0_io_pipe_phv_out_data_97; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_98 = mau_0_io_pipe_phv_out_data_98; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_99 = mau_0_io_pipe_phv_out_data_99; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_100 = mau_0_io_pipe_phv_out_data_100; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_101 = mau_0_io_pipe_phv_out_data_101; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_102 = mau_0_io_pipe_phv_out_data_102; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_103 = mau_0_io_pipe_phv_out_data_103; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_104 = mau_0_io_pipe_phv_out_data_104; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_105 = mau_0_io_pipe_phv_out_data_105; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_106 = mau_0_io_pipe_phv_out_data_106; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_107 = mau_0_io_pipe_phv_out_data_107; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_108 = mau_0_io_pipe_phv_out_data_108; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_109 = mau_0_io_pipe_phv_out_data_109; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_110 = mau_0_io_pipe_phv_out_data_110; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_111 = mau_0_io_pipe_phv_out_data_111; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_112 = mau_0_io_pipe_phv_out_data_112; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_113 = mau_0_io_pipe_phv_out_data_113; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_114 = mau_0_io_pipe_phv_out_data_114; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_115 = mau_0_io_pipe_phv_out_data_115; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_116 = mau_0_io_pipe_phv_out_data_116; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_117 = mau_0_io_pipe_phv_out_data_117; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_118 = mau_0_io_pipe_phv_out_data_118; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_119 = mau_0_io_pipe_phv_out_data_119; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_120 = mau_0_io_pipe_phv_out_data_120; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_121 = mau_0_io_pipe_phv_out_data_121; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_122 = mau_0_io_pipe_phv_out_data_122; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_123 = mau_0_io_pipe_phv_out_data_123; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_124 = mau_0_io_pipe_phv_out_data_124; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_125 = mau_0_io_pipe_phv_out_data_125; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_126 = mau_0_io_pipe_phv_out_data_126; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_127 = mau_0_io_pipe_phv_out_data_127; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_128 = mau_0_io_pipe_phv_out_data_128; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_129 = mau_0_io_pipe_phv_out_data_129; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_130 = mau_0_io_pipe_phv_out_data_130; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_131 = mau_0_io_pipe_phv_out_data_131; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_132 = mau_0_io_pipe_phv_out_data_132; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_133 = mau_0_io_pipe_phv_out_data_133; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_134 = mau_0_io_pipe_phv_out_data_134; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_135 = mau_0_io_pipe_phv_out_data_135; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_136 = mau_0_io_pipe_phv_out_data_136; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_137 = mau_0_io_pipe_phv_out_data_137; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_138 = mau_0_io_pipe_phv_out_data_138; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_139 = mau_0_io_pipe_phv_out_data_139; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_140 = mau_0_io_pipe_phv_out_data_140; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_141 = mau_0_io_pipe_phv_out_data_141; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_142 = mau_0_io_pipe_phv_out_data_142; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_143 = mau_0_io_pipe_phv_out_data_143; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_144 = mau_0_io_pipe_phv_out_data_144; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_145 = mau_0_io_pipe_phv_out_data_145; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_146 = mau_0_io_pipe_phv_out_data_146; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_147 = mau_0_io_pipe_phv_out_data_147; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_148 = mau_0_io_pipe_phv_out_data_148; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_149 = mau_0_io_pipe_phv_out_data_149; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_150 = mau_0_io_pipe_phv_out_data_150; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_151 = mau_0_io_pipe_phv_out_data_151; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_152 = mau_0_io_pipe_phv_out_data_152; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_153 = mau_0_io_pipe_phv_out_data_153; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_154 = mau_0_io_pipe_phv_out_data_154; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_155 = mau_0_io_pipe_phv_out_data_155; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_156 = mau_0_io_pipe_phv_out_data_156; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_157 = mau_0_io_pipe_phv_out_data_157; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_158 = mau_0_io_pipe_phv_out_data_158; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_159 = mau_0_io_pipe_phv_out_data_159; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_160 = mau_0_io_pipe_phv_out_data_160; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_161 = mau_0_io_pipe_phv_out_data_161; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_162 = mau_0_io_pipe_phv_out_data_162; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_163 = mau_0_io_pipe_phv_out_data_163; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_164 = mau_0_io_pipe_phv_out_data_164; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_165 = mau_0_io_pipe_phv_out_data_165; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_166 = mau_0_io_pipe_phv_out_data_166; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_167 = mau_0_io_pipe_phv_out_data_167; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_168 = mau_0_io_pipe_phv_out_data_168; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_169 = mau_0_io_pipe_phv_out_data_169; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_170 = mau_0_io_pipe_phv_out_data_170; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_171 = mau_0_io_pipe_phv_out_data_171; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_172 = mau_0_io_pipe_phv_out_data_172; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_173 = mau_0_io_pipe_phv_out_data_173; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_174 = mau_0_io_pipe_phv_out_data_174; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_175 = mau_0_io_pipe_phv_out_data_175; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_176 = mau_0_io_pipe_phv_out_data_176; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_177 = mau_0_io_pipe_phv_out_data_177; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_178 = mau_0_io_pipe_phv_out_data_178; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_179 = mau_0_io_pipe_phv_out_data_179; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_180 = mau_0_io_pipe_phv_out_data_180; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_181 = mau_0_io_pipe_phv_out_data_181; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_182 = mau_0_io_pipe_phv_out_data_182; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_183 = mau_0_io_pipe_phv_out_data_183; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_184 = mau_0_io_pipe_phv_out_data_184; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_185 = mau_0_io_pipe_phv_out_data_185; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_186 = mau_0_io_pipe_phv_out_data_186; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_187 = mau_0_io_pipe_phv_out_data_187; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_188 = mau_0_io_pipe_phv_out_data_188; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_189 = mau_0_io_pipe_phv_out_data_189; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_190 = mau_0_io_pipe_phv_out_data_190; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_191 = mau_0_io_pipe_phv_out_data_191; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_192 = mau_0_io_pipe_phv_out_data_192; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_193 = mau_0_io_pipe_phv_out_data_193; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_194 = mau_0_io_pipe_phv_out_data_194; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_195 = mau_0_io_pipe_phv_out_data_195; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_196 = mau_0_io_pipe_phv_out_data_196; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_197 = mau_0_io_pipe_phv_out_data_197; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_198 = mau_0_io_pipe_phv_out_data_198; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_199 = mau_0_io_pipe_phv_out_data_199; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_200 = mau_0_io_pipe_phv_out_data_200; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_201 = mau_0_io_pipe_phv_out_data_201; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_202 = mau_0_io_pipe_phv_out_data_202; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_203 = mau_0_io_pipe_phv_out_data_203; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_204 = mau_0_io_pipe_phv_out_data_204; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_205 = mau_0_io_pipe_phv_out_data_205; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_206 = mau_0_io_pipe_phv_out_data_206; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_207 = mau_0_io_pipe_phv_out_data_207; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_208 = mau_0_io_pipe_phv_out_data_208; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_209 = mau_0_io_pipe_phv_out_data_209; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_210 = mau_0_io_pipe_phv_out_data_210; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_211 = mau_0_io_pipe_phv_out_data_211; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_212 = mau_0_io_pipe_phv_out_data_212; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_213 = mau_0_io_pipe_phv_out_data_213; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_214 = mau_0_io_pipe_phv_out_data_214; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_215 = mau_0_io_pipe_phv_out_data_215; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_216 = mau_0_io_pipe_phv_out_data_216; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_217 = mau_0_io_pipe_phv_out_data_217; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_218 = mau_0_io_pipe_phv_out_data_218; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_219 = mau_0_io_pipe_phv_out_data_219; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_220 = mau_0_io_pipe_phv_out_data_220; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_221 = mau_0_io_pipe_phv_out_data_221; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_222 = mau_0_io_pipe_phv_out_data_222; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_223 = mau_0_io_pipe_phv_out_data_223; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_224 = mau_0_io_pipe_phv_out_data_224; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_225 = mau_0_io_pipe_phv_out_data_225; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_226 = mau_0_io_pipe_phv_out_data_226; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_227 = mau_0_io_pipe_phv_out_data_227; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_228 = mau_0_io_pipe_phv_out_data_228; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_229 = mau_0_io_pipe_phv_out_data_229; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_230 = mau_0_io_pipe_phv_out_data_230; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_231 = mau_0_io_pipe_phv_out_data_231; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_232 = mau_0_io_pipe_phv_out_data_232; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_233 = mau_0_io_pipe_phv_out_data_233; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_234 = mau_0_io_pipe_phv_out_data_234; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_235 = mau_0_io_pipe_phv_out_data_235; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_236 = mau_0_io_pipe_phv_out_data_236; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_237 = mau_0_io_pipe_phv_out_data_237; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_238 = mau_0_io_pipe_phv_out_data_238; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_239 = mau_0_io_pipe_phv_out_data_239; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_240 = mau_0_io_pipe_phv_out_data_240; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_241 = mau_0_io_pipe_phv_out_data_241; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_242 = mau_0_io_pipe_phv_out_data_242; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_243 = mau_0_io_pipe_phv_out_data_243; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_244 = mau_0_io_pipe_phv_out_data_244; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_245 = mau_0_io_pipe_phv_out_data_245; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_246 = mau_0_io_pipe_phv_out_data_246; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_247 = mau_0_io_pipe_phv_out_data_247; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_248 = mau_0_io_pipe_phv_out_data_248; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_249 = mau_0_io_pipe_phv_out_data_249; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_250 = mau_0_io_pipe_phv_out_data_250; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_251 = mau_0_io_pipe_phv_out_data_251; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_252 = mau_0_io_pipe_phv_out_data_252; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_253 = mau_0_io_pipe_phv_out_data_253; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_254 = mau_0_io_pipe_phv_out_data_254; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_255 = mau_0_io_pipe_phv_out_data_255; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_header_0 = mau_0_io_pipe_phv_out_header_0; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_header_1 = mau_0_io_pipe_phv_out_header_1; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_header_2 = mau_0_io_pipe_phv_out_header_2; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_header_3 = mau_0_io_pipe_phv_out_header_3; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_header_4 = mau_0_io_pipe_phv_out_header_4; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_header_5 = mau_0_io_pipe_phv_out_header_5; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_header_6 = mau_0_io_pipe_phv_out_header_6; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_header_7 = mau_0_io_pipe_phv_out_header_7; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_header_8 = mau_0_io_pipe_phv_out_header_8; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_header_9 = mau_0_io_pipe_phv_out_header_9; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_header_10 = mau_0_io_pipe_phv_out_header_10; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_header_11 = mau_0_io_pipe_phv_out_header_11; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_header_12 = mau_0_io_pipe_phv_out_header_12; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_header_13 = mau_0_io_pipe_phv_out_header_13; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_header_14 = mau_0_io_pipe_phv_out_header_14; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_header_15 = mau_0_io_pipe_phv_out_header_15; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_parse_current_state = mau_0_io_pipe_phv_out_parse_current_state; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_parse_current_offset = mau_0_io_pipe_phv_out_parse_current_offset; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_parse_transition_field = mau_0_io_pipe_phv_out_parse_transition_field; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_next_processor_id = mau_0_io_pipe_phv_out_next_processor_id; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_next_config_id = mau_0_io_pipe_phv_out_next_config_id; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_is_valid_processor = mau_0_io_pipe_phv_out_is_valid_processor; // @[parser.scala 32:35]
  assign mau_1_io_mod_state_id_mod = io_mod_en ? io_mod_module_mod_state_id_mod & mod_j_1 :
    io_mod_module_mod_state_id_mod; // @[parser.scala 41:22 parser.scala 48:40 parser.scala 37:23]
  assign mau_1_io_mod_state_id = io_mod_module_mod_state_id; // @[parser.scala 37:23]
  assign mau_1_io_mod_sram_w_cs = io_mod_module_mod_sram_w_cs; // @[parser.scala 37:23]
  assign mau_1_io_mod_sram_w_en = io_mod_en ? io_mod_module_mod_sram_w_en & mod_j_1 : io_mod_module_mod_sram_w_en; // @[parser.scala 41:22 parser.scala 47:40 parser.scala 37:23]
  assign mau_1_io_mod_sram_w_addr = io_mod_module_mod_sram_w_addr; // @[parser.scala 37:23]
  assign mau_1_io_mod_sram_w_data = io_mod_module_mod_sram_w_data; // @[parser.scala 37:23]
  assign mau_2_clock = clock;
  assign mau_2_io_pipe_phv_in_data_0 = mau_1_io_pipe_phv_out_data_0; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_1 = mau_1_io_pipe_phv_out_data_1; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_2 = mau_1_io_pipe_phv_out_data_2; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_3 = mau_1_io_pipe_phv_out_data_3; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_4 = mau_1_io_pipe_phv_out_data_4; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_5 = mau_1_io_pipe_phv_out_data_5; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_6 = mau_1_io_pipe_phv_out_data_6; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_7 = mau_1_io_pipe_phv_out_data_7; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_8 = mau_1_io_pipe_phv_out_data_8; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_9 = mau_1_io_pipe_phv_out_data_9; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_10 = mau_1_io_pipe_phv_out_data_10; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_11 = mau_1_io_pipe_phv_out_data_11; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_12 = mau_1_io_pipe_phv_out_data_12; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_13 = mau_1_io_pipe_phv_out_data_13; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_14 = mau_1_io_pipe_phv_out_data_14; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_15 = mau_1_io_pipe_phv_out_data_15; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_16 = mau_1_io_pipe_phv_out_data_16; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_17 = mau_1_io_pipe_phv_out_data_17; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_18 = mau_1_io_pipe_phv_out_data_18; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_19 = mau_1_io_pipe_phv_out_data_19; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_20 = mau_1_io_pipe_phv_out_data_20; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_21 = mau_1_io_pipe_phv_out_data_21; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_22 = mau_1_io_pipe_phv_out_data_22; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_23 = mau_1_io_pipe_phv_out_data_23; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_24 = mau_1_io_pipe_phv_out_data_24; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_25 = mau_1_io_pipe_phv_out_data_25; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_26 = mau_1_io_pipe_phv_out_data_26; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_27 = mau_1_io_pipe_phv_out_data_27; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_28 = mau_1_io_pipe_phv_out_data_28; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_29 = mau_1_io_pipe_phv_out_data_29; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_30 = mau_1_io_pipe_phv_out_data_30; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_31 = mau_1_io_pipe_phv_out_data_31; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_32 = mau_1_io_pipe_phv_out_data_32; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_33 = mau_1_io_pipe_phv_out_data_33; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_34 = mau_1_io_pipe_phv_out_data_34; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_35 = mau_1_io_pipe_phv_out_data_35; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_36 = mau_1_io_pipe_phv_out_data_36; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_37 = mau_1_io_pipe_phv_out_data_37; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_38 = mau_1_io_pipe_phv_out_data_38; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_39 = mau_1_io_pipe_phv_out_data_39; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_40 = mau_1_io_pipe_phv_out_data_40; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_41 = mau_1_io_pipe_phv_out_data_41; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_42 = mau_1_io_pipe_phv_out_data_42; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_43 = mau_1_io_pipe_phv_out_data_43; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_44 = mau_1_io_pipe_phv_out_data_44; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_45 = mau_1_io_pipe_phv_out_data_45; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_46 = mau_1_io_pipe_phv_out_data_46; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_47 = mau_1_io_pipe_phv_out_data_47; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_48 = mau_1_io_pipe_phv_out_data_48; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_49 = mau_1_io_pipe_phv_out_data_49; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_50 = mau_1_io_pipe_phv_out_data_50; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_51 = mau_1_io_pipe_phv_out_data_51; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_52 = mau_1_io_pipe_phv_out_data_52; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_53 = mau_1_io_pipe_phv_out_data_53; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_54 = mau_1_io_pipe_phv_out_data_54; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_55 = mau_1_io_pipe_phv_out_data_55; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_56 = mau_1_io_pipe_phv_out_data_56; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_57 = mau_1_io_pipe_phv_out_data_57; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_58 = mau_1_io_pipe_phv_out_data_58; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_59 = mau_1_io_pipe_phv_out_data_59; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_60 = mau_1_io_pipe_phv_out_data_60; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_61 = mau_1_io_pipe_phv_out_data_61; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_62 = mau_1_io_pipe_phv_out_data_62; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_63 = mau_1_io_pipe_phv_out_data_63; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_64 = mau_1_io_pipe_phv_out_data_64; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_65 = mau_1_io_pipe_phv_out_data_65; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_66 = mau_1_io_pipe_phv_out_data_66; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_67 = mau_1_io_pipe_phv_out_data_67; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_68 = mau_1_io_pipe_phv_out_data_68; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_69 = mau_1_io_pipe_phv_out_data_69; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_70 = mau_1_io_pipe_phv_out_data_70; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_71 = mau_1_io_pipe_phv_out_data_71; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_72 = mau_1_io_pipe_phv_out_data_72; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_73 = mau_1_io_pipe_phv_out_data_73; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_74 = mau_1_io_pipe_phv_out_data_74; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_75 = mau_1_io_pipe_phv_out_data_75; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_76 = mau_1_io_pipe_phv_out_data_76; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_77 = mau_1_io_pipe_phv_out_data_77; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_78 = mau_1_io_pipe_phv_out_data_78; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_79 = mau_1_io_pipe_phv_out_data_79; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_80 = mau_1_io_pipe_phv_out_data_80; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_81 = mau_1_io_pipe_phv_out_data_81; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_82 = mau_1_io_pipe_phv_out_data_82; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_83 = mau_1_io_pipe_phv_out_data_83; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_84 = mau_1_io_pipe_phv_out_data_84; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_85 = mau_1_io_pipe_phv_out_data_85; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_86 = mau_1_io_pipe_phv_out_data_86; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_87 = mau_1_io_pipe_phv_out_data_87; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_88 = mau_1_io_pipe_phv_out_data_88; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_89 = mau_1_io_pipe_phv_out_data_89; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_90 = mau_1_io_pipe_phv_out_data_90; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_91 = mau_1_io_pipe_phv_out_data_91; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_92 = mau_1_io_pipe_phv_out_data_92; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_93 = mau_1_io_pipe_phv_out_data_93; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_94 = mau_1_io_pipe_phv_out_data_94; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_95 = mau_1_io_pipe_phv_out_data_95; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_96 = mau_1_io_pipe_phv_out_data_96; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_97 = mau_1_io_pipe_phv_out_data_97; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_98 = mau_1_io_pipe_phv_out_data_98; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_99 = mau_1_io_pipe_phv_out_data_99; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_100 = mau_1_io_pipe_phv_out_data_100; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_101 = mau_1_io_pipe_phv_out_data_101; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_102 = mau_1_io_pipe_phv_out_data_102; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_103 = mau_1_io_pipe_phv_out_data_103; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_104 = mau_1_io_pipe_phv_out_data_104; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_105 = mau_1_io_pipe_phv_out_data_105; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_106 = mau_1_io_pipe_phv_out_data_106; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_107 = mau_1_io_pipe_phv_out_data_107; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_108 = mau_1_io_pipe_phv_out_data_108; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_109 = mau_1_io_pipe_phv_out_data_109; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_110 = mau_1_io_pipe_phv_out_data_110; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_111 = mau_1_io_pipe_phv_out_data_111; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_112 = mau_1_io_pipe_phv_out_data_112; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_113 = mau_1_io_pipe_phv_out_data_113; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_114 = mau_1_io_pipe_phv_out_data_114; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_115 = mau_1_io_pipe_phv_out_data_115; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_116 = mau_1_io_pipe_phv_out_data_116; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_117 = mau_1_io_pipe_phv_out_data_117; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_118 = mau_1_io_pipe_phv_out_data_118; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_119 = mau_1_io_pipe_phv_out_data_119; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_120 = mau_1_io_pipe_phv_out_data_120; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_121 = mau_1_io_pipe_phv_out_data_121; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_122 = mau_1_io_pipe_phv_out_data_122; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_123 = mau_1_io_pipe_phv_out_data_123; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_124 = mau_1_io_pipe_phv_out_data_124; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_125 = mau_1_io_pipe_phv_out_data_125; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_126 = mau_1_io_pipe_phv_out_data_126; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_127 = mau_1_io_pipe_phv_out_data_127; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_128 = mau_1_io_pipe_phv_out_data_128; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_129 = mau_1_io_pipe_phv_out_data_129; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_130 = mau_1_io_pipe_phv_out_data_130; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_131 = mau_1_io_pipe_phv_out_data_131; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_132 = mau_1_io_pipe_phv_out_data_132; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_133 = mau_1_io_pipe_phv_out_data_133; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_134 = mau_1_io_pipe_phv_out_data_134; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_135 = mau_1_io_pipe_phv_out_data_135; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_136 = mau_1_io_pipe_phv_out_data_136; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_137 = mau_1_io_pipe_phv_out_data_137; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_138 = mau_1_io_pipe_phv_out_data_138; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_139 = mau_1_io_pipe_phv_out_data_139; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_140 = mau_1_io_pipe_phv_out_data_140; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_141 = mau_1_io_pipe_phv_out_data_141; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_142 = mau_1_io_pipe_phv_out_data_142; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_143 = mau_1_io_pipe_phv_out_data_143; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_144 = mau_1_io_pipe_phv_out_data_144; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_145 = mau_1_io_pipe_phv_out_data_145; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_146 = mau_1_io_pipe_phv_out_data_146; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_147 = mau_1_io_pipe_phv_out_data_147; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_148 = mau_1_io_pipe_phv_out_data_148; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_149 = mau_1_io_pipe_phv_out_data_149; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_150 = mau_1_io_pipe_phv_out_data_150; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_151 = mau_1_io_pipe_phv_out_data_151; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_152 = mau_1_io_pipe_phv_out_data_152; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_153 = mau_1_io_pipe_phv_out_data_153; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_154 = mau_1_io_pipe_phv_out_data_154; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_155 = mau_1_io_pipe_phv_out_data_155; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_156 = mau_1_io_pipe_phv_out_data_156; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_157 = mau_1_io_pipe_phv_out_data_157; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_158 = mau_1_io_pipe_phv_out_data_158; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_159 = mau_1_io_pipe_phv_out_data_159; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_160 = mau_1_io_pipe_phv_out_data_160; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_161 = mau_1_io_pipe_phv_out_data_161; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_162 = mau_1_io_pipe_phv_out_data_162; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_163 = mau_1_io_pipe_phv_out_data_163; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_164 = mau_1_io_pipe_phv_out_data_164; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_165 = mau_1_io_pipe_phv_out_data_165; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_166 = mau_1_io_pipe_phv_out_data_166; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_167 = mau_1_io_pipe_phv_out_data_167; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_168 = mau_1_io_pipe_phv_out_data_168; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_169 = mau_1_io_pipe_phv_out_data_169; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_170 = mau_1_io_pipe_phv_out_data_170; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_171 = mau_1_io_pipe_phv_out_data_171; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_172 = mau_1_io_pipe_phv_out_data_172; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_173 = mau_1_io_pipe_phv_out_data_173; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_174 = mau_1_io_pipe_phv_out_data_174; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_175 = mau_1_io_pipe_phv_out_data_175; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_176 = mau_1_io_pipe_phv_out_data_176; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_177 = mau_1_io_pipe_phv_out_data_177; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_178 = mau_1_io_pipe_phv_out_data_178; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_179 = mau_1_io_pipe_phv_out_data_179; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_180 = mau_1_io_pipe_phv_out_data_180; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_181 = mau_1_io_pipe_phv_out_data_181; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_182 = mau_1_io_pipe_phv_out_data_182; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_183 = mau_1_io_pipe_phv_out_data_183; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_184 = mau_1_io_pipe_phv_out_data_184; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_185 = mau_1_io_pipe_phv_out_data_185; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_186 = mau_1_io_pipe_phv_out_data_186; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_187 = mau_1_io_pipe_phv_out_data_187; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_188 = mau_1_io_pipe_phv_out_data_188; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_189 = mau_1_io_pipe_phv_out_data_189; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_190 = mau_1_io_pipe_phv_out_data_190; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_191 = mau_1_io_pipe_phv_out_data_191; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_192 = mau_1_io_pipe_phv_out_data_192; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_193 = mau_1_io_pipe_phv_out_data_193; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_194 = mau_1_io_pipe_phv_out_data_194; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_195 = mau_1_io_pipe_phv_out_data_195; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_196 = mau_1_io_pipe_phv_out_data_196; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_197 = mau_1_io_pipe_phv_out_data_197; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_198 = mau_1_io_pipe_phv_out_data_198; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_199 = mau_1_io_pipe_phv_out_data_199; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_200 = mau_1_io_pipe_phv_out_data_200; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_201 = mau_1_io_pipe_phv_out_data_201; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_202 = mau_1_io_pipe_phv_out_data_202; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_203 = mau_1_io_pipe_phv_out_data_203; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_204 = mau_1_io_pipe_phv_out_data_204; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_205 = mau_1_io_pipe_phv_out_data_205; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_206 = mau_1_io_pipe_phv_out_data_206; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_207 = mau_1_io_pipe_phv_out_data_207; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_208 = mau_1_io_pipe_phv_out_data_208; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_209 = mau_1_io_pipe_phv_out_data_209; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_210 = mau_1_io_pipe_phv_out_data_210; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_211 = mau_1_io_pipe_phv_out_data_211; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_212 = mau_1_io_pipe_phv_out_data_212; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_213 = mau_1_io_pipe_phv_out_data_213; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_214 = mau_1_io_pipe_phv_out_data_214; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_215 = mau_1_io_pipe_phv_out_data_215; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_216 = mau_1_io_pipe_phv_out_data_216; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_217 = mau_1_io_pipe_phv_out_data_217; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_218 = mau_1_io_pipe_phv_out_data_218; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_219 = mau_1_io_pipe_phv_out_data_219; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_220 = mau_1_io_pipe_phv_out_data_220; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_221 = mau_1_io_pipe_phv_out_data_221; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_222 = mau_1_io_pipe_phv_out_data_222; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_223 = mau_1_io_pipe_phv_out_data_223; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_224 = mau_1_io_pipe_phv_out_data_224; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_225 = mau_1_io_pipe_phv_out_data_225; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_226 = mau_1_io_pipe_phv_out_data_226; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_227 = mau_1_io_pipe_phv_out_data_227; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_228 = mau_1_io_pipe_phv_out_data_228; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_229 = mau_1_io_pipe_phv_out_data_229; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_230 = mau_1_io_pipe_phv_out_data_230; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_231 = mau_1_io_pipe_phv_out_data_231; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_232 = mau_1_io_pipe_phv_out_data_232; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_233 = mau_1_io_pipe_phv_out_data_233; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_234 = mau_1_io_pipe_phv_out_data_234; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_235 = mau_1_io_pipe_phv_out_data_235; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_236 = mau_1_io_pipe_phv_out_data_236; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_237 = mau_1_io_pipe_phv_out_data_237; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_238 = mau_1_io_pipe_phv_out_data_238; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_239 = mau_1_io_pipe_phv_out_data_239; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_240 = mau_1_io_pipe_phv_out_data_240; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_241 = mau_1_io_pipe_phv_out_data_241; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_242 = mau_1_io_pipe_phv_out_data_242; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_243 = mau_1_io_pipe_phv_out_data_243; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_244 = mau_1_io_pipe_phv_out_data_244; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_245 = mau_1_io_pipe_phv_out_data_245; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_246 = mau_1_io_pipe_phv_out_data_246; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_247 = mau_1_io_pipe_phv_out_data_247; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_248 = mau_1_io_pipe_phv_out_data_248; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_249 = mau_1_io_pipe_phv_out_data_249; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_250 = mau_1_io_pipe_phv_out_data_250; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_251 = mau_1_io_pipe_phv_out_data_251; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_252 = mau_1_io_pipe_phv_out_data_252; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_253 = mau_1_io_pipe_phv_out_data_253; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_254 = mau_1_io_pipe_phv_out_data_254; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_255 = mau_1_io_pipe_phv_out_data_255; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_header_0 = mau_1_io_pipe_phv_out_header_0; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_header_1 = mau_1_io_pipe_phv_out_header_1; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_header_2 = mau_1_io_pipe_phv_out_header_2; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_header_3 = mau_1_io_pipe_phv_out_header_3; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_header_4 = mau_1_io_pipe_phv_out_header_4; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_header_5 = mau_1_io_pipe_phv_out_header_5; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_header_6 = mau_1_io_pipe_phv_out_header_6; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_header_7 = mau_1_io_pipe_phv_out_header_7; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_header_8 = mau_1_io_pipe_phv_out_header_8; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_header_9 = mau_1_io_pipe_phv_out_header_9; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_header_10 = mau_1_io_pipe_phv_out_header_10; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_header_11 = mau_1_io_pipe_phv_out_header_11; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_header_12 = mau_1_io_pipe_phv_out_header_12; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_header_13 = mau_1_io_pipe_phv_out_header_13; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_header_14 = mau_1_io_pipe_phv_out_header_14; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_header_15 = mau_1_io_pipe_phv_out_header_15; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_parse_current_state = mau_1_io_pipe_phv_out_parse_current_state; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_parse_current_offset = mau_1_io_pipe_phv_out_parse_current_offset; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_parse_transition_field = mau_1_io_pipe_phv_out_parse_transition_field; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_next_processor_id = mau_1_io_pipe_phv_out_next_processor_id; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_next_config_id = mau_1_io_pipe_phv_out_next_config_id; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_is_valid_processor = mau_1_io_pipe_phv_out_is_valid_processor; // @[parser.scala 32:35]
  assign mau_2_io_mod_state_id_mod = io_mod_en ? io_mod_module_mod_state_id_mod & mod_j_2 :
    io_mod_module_mod_state_id_mod; // @[parser.scala 41:22 parser.scala 48:40 parser.scala 37:23]
  assign mau_2_io_mod_state_id = io_mod_module_mod_state_id; // @[parser.scala 37:23]
  assign mau_2_io_mod_sram_w_cs = io_mod_module_mod_sram_w_cs; // @[parser.scala 37:23]
  assign mau_2_io_mod_sram_w_en = io_mod_en ? io_mod_module_mod_sram_w_en & mod_j_2 : io_mod_module_mod_sram_w_en; // @[parser.scala 41:22 parser.scala 47:40 parser.scala 37:23]
  assign mau_2_io_mod_sram_w_addr = io_mod_module_mod_sram_w_addr; // @[parser.scala 37:23]
  assign mau_2_io_mod_sram_w_data = io_mod_module_mod_sram_w_data; // @[parser.scala 37:23]
  assign mau_3_clock = clock;
  assign mau_3_io_pipe_phv_in_data_0 = mau_2_io_pipe_phv_out_data_0; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_1 = mau_2_io_pipe_phv_out_data_1; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_2 = mau_2_io_pipe_phv_out_data_2; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_3 = mau_2_io_pipe_phv_out_data_3; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_4 = mau_2_io_pipe_phv_out_data_4; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_5 = mau_2_io_pipe_phv_out_data_5; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_6 = mau_2_io_pipe_phv_out_data_6; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_7 = mau_2_io_pipe_phv_out_data_7; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_8 = mau_2_io_pipe_phv_out_data_8; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_9 = mau_2_io_pipe_phv_out_data_9; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_10 = mau_2_io_pipe_phv_out_data_10; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_11 = mau_2_io_pipe_phv_out_data_11; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_12 = mau_2_io_pipe_phv_out_data_12; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_13 = mau_2_io_pipe_phv_out_data_13; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_14 = mau_2_io_pipe_phv_out_data_14; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_15 = mau_2_io_pipe_phv_out_data_15; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_16 = mau_2_io_pipe_phv_out_data_16; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_17 = mau_2_io_pipe_phv_out_data_17; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_18 = mau_2_io_pipe_phv_out_data_18; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_19 = mau_2_io_pipe_phv_out_data_19; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_20 = mau_2_io_pipe_phv_out_data_20; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_21 = mau_2_io_pipe_phv_out_data_21; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_22 = mau_2_io_pipe_phv_out_data_22; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_23 = mau_2_io_pipe_phv_out_data_23; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_24 = mau_2_io_pipe_phv_out_data_24; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_25 = mau_2_io_pipe_phv_out_data_25; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_26 = mau_2_io_pipe_phv_out_data_26; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_27 = mau_2_io_pipe_phv_out_data_27; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_28 = mau_2_io_pipe_phv_out_data_28; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_29 = mau_2_io_pipe_phv_out_data_29; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_30 = mau_2_io_pipe_phv_out_data_30; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_31 = mau_2_io_pipe_phv_out_data_31; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_32 = mau_2_io_pipe_phv_out_data_32; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_33 = mau_2_io_pipe_phv_out_data_33; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_34 = mau_2_io_pipe_phv_out_data_34; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_35 = mau_2_io_pipe_phv_out_data_35; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_36 = mau_2_io_pipe_phv_out_data_36; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_37 = mau_2_io_pipe_phv_out_data_37; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_38 = mau_2_io_pipe_phv_out_data_38; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_39 = mau_2_io_pipe_phv_out_data_39; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_40 = mau_2_io_pipe_phv_out_data_40; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_41 = mau_2_io_pipe_phv_out_data_41; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_42 = mau_2_io_pipe_phv_out_data_42; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_43 = mau_2_io_pipe_phv_out_data_43; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_44 = mau_2_io_pipe_phv_out_data_44; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_45 = mau_2_io_pipe_phv_out_data_45; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_46 = mau_2_io_pipe_phv_out_data_46; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_47 = mau_2_io_pipe_phv_out_data_47; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_48 = mau_2_io_pipe_phv_out_data_48; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_49 = mau_2_io_pipe_phv_out_data_49; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_50 = mau_2_io_pipe_phv_out_data_50; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_51 = mau_2_io_pipe_phv_out_data_51; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_52 = mau_2_io_pipe_phv_out_data_52; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_53 = mau_2_io_pipe_phv_out_data_53; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_54 = mau_2_io_pipe_phv_out_data_54; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_55 = mau_2_io_pipe_phv_out_data_55; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_56 = mau_2_io_pipe_phv_out_data_56; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_57 = mau_2_io_pipe_phv_out_data_57; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_58 = mau_2_io_pipe_phv_out_data_58; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_59 = mau_2_io_pipe_phv_out_data_59; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_60 = mau_2_io_pipe_phv_out_data_60; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_61 = mau_2_io_pipe_phv_out_data_61; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_62 = mau_2_io_pipe_phv_out_data_62; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_63 = mau_2_io_pipe_phv_out_data_63; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_64 = mau_2_io_pipe_phv_out_data_64; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_65 = mau_2_io_pipe_phv_out_data_65; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_66 = mau_2_io_pipe_phv_out_data_66; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_67 = mau_2_io_pipe_phv_out_data_67; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_68 = mau_2_io_pipe_phv_out_data_68; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_69 = mau_2_io_pipe_phv_out_data_69; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_70 = mau_2_io_pipe_phv_out_data_70; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_71 = mau_2_io_pipe_phv_out_data_71; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_72 = mau_2_io_pipe_phv_out_data_72; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_73 = mau_2_io_pipe_phv_out_data_73; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_74 = mau_2_io_pipe_phv_out_data_74; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_75 = mau_2_io_pipe_phv_out_data_75; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_76 = mau_2_io_pipe_phv_out_data_76; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_77 = mau_2_io_pipe_phv_out_data_77; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_78 = mau_2_io_pipe_phv_out_data_78; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_79 = mau_2_io_pipe_phv_out_data_79; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_80 = mau_2_io_pipe_phv_out_data_80; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_81 = mau_2_io_pipe_phv_out_data_81; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_82 = mau_2_io_pipe_phv_out_data_82; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_83 = mau_2_io_pipe_phv_out_data_83; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_84 = mau_2_io_pipe_phv_out_data_84; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_85 = mau_2_io_pipe_phv_out_data_85; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_86 = mau_2_io_pipe_phv_out_data_86; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_87 = mau_2_io_pipe_phv_out_data_87; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_88 = mau_2_io_pipe_phv_out_data_88; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_89 = mau_2_io_pipe_phv_out_data_89; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_90 = mau_2_io_pipe_phv_out_data_90; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_91 = mau_2_io_pipe_phv_out_data_91; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_92 = mau_2_io_pipe_phv_out_data_92; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_93 = mau_2_io_pipe_phv_out_data_93; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_94 = mau_2_io_pipe_phv_out_data_94; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_95 = mau_2_io_pipe_phv_out_data_95; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_96 = mau_2_io_pipe_phv_out_data_96; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_97 = mau_2_io_pipe_phv_out_data_97; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_98 = mau_2_io_pipe_phv_out_data_98; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_99 = mau_2_io_pipe_phv_out_data_99; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_100 = mau_2_io_pipe_phv_out_data_100; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_101 = mau_2_io_pipe_phv_out_data_101; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_102 = mau_2_io_pipe_phv_out_data_102; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_103 = mau_2_io_pipe_phv_out_data_103; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_104 = mau_2_io_pipe_phv_out_data_104; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_105 = mau_2_io_pipe_phv_out_data_105; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_106 = mau_2_io_pipe_phv_out_data_106; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_107 = mau_2_io_pipe_phv_out_data_107; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_108 = mau_2_io_pipe_phv_out_data_108; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_109 = mau_2_io_pipe_phv_out_data_109; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_110 = mau_2_io_pipe_phv_out_data_110; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_111 = mau_2_io_pipe_phv_out_data_111; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_112 = mau_2_io_pipe_phv_out_data_112; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_113 = mau_2_io_pipe_phv_out_data_113; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_114 = mau_2_io_pipe_phv_out_data_114; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_115 = mau_2_io_pipe_phv_out_data_115; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_116 = mau_2_io_pipe_phv_out_data_116; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_117 = mau_2_io_pipe_phv_out_data_117; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_118 = mau_2_io_pipe_phv_out_data_118; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_119 = mau_2_io_pipe_phv_out_data_119; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_120 = mau_2_io_pipe_phv_out_data_120; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_121 = mau_2_io_pipe_phv_out_data_121; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_122 = mau_2_io_pipe_phv_out_data_122; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_123 = mau_2_io_pipe_phv_out_data_123; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_124 = mau_2_io_pipe_phv_out_data_124; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_125 = mau_2_io_pipe_phv_out_data_125; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_126 = mau_2_io_pipe_phv_out_data_126; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_127 = mau_2_io_pipe_phv_out_data_127; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_128 = mau_2_io_pipe_phv_out_data_128; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_129 = mau_2_io_pipe_phv_out_data_129; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_130 = mau_2_io_pipe_phv_out_data_130; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_131 = mau_2_io_pipe_phv_out_data_131; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_132 = mau_2_io_pipe_phv_out_data_132; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_133 = mau_2_io_pipe_phv_out_data_133; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_134 = mau_2_io_pipe_phv_out_data_134; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_135 = mau_2_io_pipe_phv_out_data_135; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_136 = mau_2_io_pipe_phv_out_data_136; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_137 = mau_2_io_pipe_phv_out_data_137; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_138 = mau_2_io_pipe_phv_out_data_138; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_139 = mau_2_io_pipe_phv_out_data_139; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_140 = mau_2_io_pipe_phv_out_data_140; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_141 = mau_2_io_pipe_phv_out_data_141; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_142 = mau_2_io_pipe_phv_out_data_142; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_143 = mau_2_io_pipe_phv_out_data_143; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_144 = mau_2_io_pipe_phv_out_data_144; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_145 = mau_2_io_pipe_phv_out_data_145; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_146 = mau_2_io_pipe_phv_out_data_146; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_147 = mau_2_io_pipe_phv_out_data_147; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_148 = mau_2_io_pipe_phv_out_data_148; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_149 = mau_2_io_pipe_phv_out_data_149; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_150 = mau_2_io_pipe_phv_out_data_150; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_151 = mau_2_io_pipe_phv_out_data_151; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_152 = mau_2_io_pipe_phv_out_data_152; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_153 = mau_2_io_pipe_phv_out_data_153; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_154 = mau_2_io_pipe_phv_out_data_154; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_155 = mau_2_io_pipe_phv_out_data_155; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_156 = mau_2_io_pipe_phv_out_data_156; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_157 = mau_2_io_pipe_phv_out_data_157; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_158 = mau_2_io_pipe_phv_out_data_158; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_159 = mau_2_io_pipe_phv_out_data_159; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_160 = mau_2_io_pipe_phv_out_data_160; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_161 = mau_2_io_pipe_phv_out_data_161; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_162 = mau_2_io_pipe_phv_out_data_162; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_163 = mau_2_io_pipe_phv_out_data_163; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_164 = mau_2_io_pipe_phv_out_data_164; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_165 = mau_2_io_pipe_phv_out_data_165; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_166 = mau_2_io_pipe_phv_out_data_166; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_167 = mau_2_io_pipe_phv_out_data_167; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_168 = mau_2_io_pipe_phv_out_data_168; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_169 = mau_2_io_pipe_phv_out_data_169; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_170 = mau_2_io_pipe_phv_out_data_170; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_171 = mau_2_io_pipe_phv_out_data_171; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_172 = mau_2_io_pipe_phv_out_data_172; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_173 = mau_2_io_pipe_phv_out_data_173; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_174 = mau_2_io_pipe_phv_out_data_174; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_175 = mau_2_io_pipe_phv_out_data_175; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_176 = mau_2_io_pipe_phv_out_data_176; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_177 = mau_2_io_pipe_phv_out_data_177; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_178 = mau_2_io_pipe_phv_out_data_178; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_179 = mau_2_io_pipe_phv_out_data_179; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_180 = mau_2_io_pipe_phv_out_data_180; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_181 = mau_2_io_pipe_phv_out_data_181; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_182 = mau_2_io_pipe_phv_out_data_182; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_183 = mau_2_io_pipe_phv_out_data_183; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_184 = mau_2_io_pipe_phv_out_data_184; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_185 = mau_2_io_pipe_phv_out_data_185; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_186 = mau_2_io_pipe_phv_out_data_186; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_187 = mau_2_io_pipe_phv_out_data_187; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_188 = mau_2_io_pipe_phv_out_data_188; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_189 = mau_2_io_pipe_phv_out_data_189; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_190 = mau_2_io_pipe_phv_out_data_190; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_191 = mau_2_io_pipe_phv_out_data_191; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_192 = mau_2_io_pipe_phv_out_data_192; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_193 = mau_2_io_pipe_phv_out_data_193; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_194 = mau_2_io_pipe_phv_out_data_194; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_195 = mau_2_io_pipe_phv_out_data_195; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_196 = mau_2_io_pipe_phv_out_data_196; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_197 = mau_2_io_pipe_phv_out_data_197; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_198 = mau_2_io_pipe_phv_out_data_198; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_199 = mau_2_io_pipe_phv_out_data_199; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_200 = mau_2_io_pipe_phv_out_data_200; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_201 = mau_2_io_pipe_phv_out_data_201; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_202 = mau_2_io_pipe_phv_out_data_202; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_203 = mau_2_io_pipe_phv_out_data_203; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_204 = mau_2_io_pipe_phv_out_data_204; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_205 = mau_2_io_pipe_phv_out_data_205; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_206 = mau_2_io_pipe_phv_out_data_206; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_207 = mau_2_io_pipe_phv_out_data_207; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_208 = mau_2_io_pipe_phv_out_data_208; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_209 = mau_2_io_pipe_phv_out_data_209; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_210 = mau_2_io_pipe_phv_out_data_210; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_211 = mau_2_io_pipe_phv_out_data_211; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_212 = mau_2_io_pipe_phv_out_data_212; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_213 = mau_2_io_pipe_phv_out_data_213; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_214 = mau_2_io_pipe_phv_out_data_214; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_215 = mau_2_io_pipe_phv_out_data_215; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_216 = mau_2_io_pipe_phv_out_data_216; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_217 = mau_2_io_pipe_phv_out_data_217; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_218 = mau_2_io_pipe_phv_out_data_218; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_219 = mau_2_io_pipe_phv_out_data_219; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_220 = mau_2_io_pipe_phv_out_data_220; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_221 = mau_2_io_pipe_phv_out_data_221; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_222 = mau_2_io_pipe_phv_out_data_222; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_223 = mau_2_io_pipe_phv_out_data_223; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_224 = mau_2_io_pipe_phv_out_data_224; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_225 = mau_2_io_pipe_phv_out_data_225; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_226 = mau_2_io_pipe_phv_out_data_226; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_227 = mau_2_io_pipe_phv_out_data_227; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_228 = mau_2_io_pipe_phv_out_data_228; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_229 = mau_2_io_pipe_phv_out_data_229; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_230 = mau_2_io_pipe_phv_out_data_230; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_231 = mau_2_io_pipe_phv_out_data_231; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_232 = mau_2_io_pipe_phv_out_data_232; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_233 = mau_2_io_pipe_phv_out_data_233; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_234 = mau_2_io_pipe_phv_out_data_234; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_235 = mau_2_io_pipe_phv_out_data_235; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_236 = mau_2_io_pipe_phv_out_data_236; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_237 = mau_2_io_pipe_phv_out_data_237; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_238 = mau_2_io_pipe_phv_out_data_238; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_239 = mau_2_io_pipe_phv_out_data_239; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_240 = mau_2_io_pipe_phv_out_data_240; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_241 = mau_2_io_pipe_phv_out_data_241; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_242 = mau_2_io_pipe_phv_out_data_242; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_243 = mau_2_io_pipe_phv_out_data_243; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_244 = mau_2_io_pipe_phv_out_data_244; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_245 = mau_2_io_pipe_phv_out_data_245; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_246 = mau_2_io_pipe_phv_out_data_246; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_247 = mau_2_io_pipe_phv_out_data_247; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_248 = mau_2_io_pipe_phv_out_data_248; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_249 = mau_2_io_pipe_phv_out_data_249; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_250 = mau_2_io_pipe_phv_out_data_250; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_251 = mau_2_io_pipe_phv_out_data_251; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_252 = mau_2_io_pipe_phv_out_data_252; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_253 = mau_2_io_pipe_phv_out_data_253; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_254 = mau_2_io_pipe_phv_out_data_254; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_255 = mau_2_io_pipe_phv_out_data_255; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_header_0 = mau_2_io_pipe_phv_out_header_0; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_header_1 = mau_2_io_pipe_phv_out_header_1; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_header_2 = mau_2_io_pipe_phv_out_header_2; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_header_3 = mau_2_io_pipe_phv_out_header_3; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_header_4 = mau_2_io_pipe_phv_out_header_4; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_header_5 = mau_2_io_pipe_phv_out_header_5; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_header_6 = mau_2_io_pipe_phv_out_header_6; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_header_7 = mau_2_io_pipe_phv_out_header_7; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_header_8 = mau_2_io_pipe_phv_out_header_8; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_header_9 = mau_2_io_pipe_phv_out_header_9; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_header_10 = mau_2_io_pipe_phv_out_header_10; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_header_11 = mau_2_io_pipe_phv_out_header_11; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_header_12 = mau_2_io_pipe_phv_out_header_12; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_header_13 = mau_2_io_pipe_phv_out_header_13; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_header_14 = mau_2_io_pipe_phv_out_header_14; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_header_15 = mau_2_io_pipe_phv_out_header_15; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_parse_current_state = mau_2_io_pipe_phv_out_parse_current_state; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_parse_current_offset = mau_2_io_pipe_phv_out_parse_current_offset; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_parse_transition_field = mau_2_io_pipe_phv_out_parse_transition_field; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_next_processor_id = mau_2_io_pipe_phv_out_next_processor_id; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_next_config_id = mau_2_io_pipe_phv_out_next_config_id; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_is_valid_processor = mau_2_io_pipe_phv_out_is_valid_processor; // @[parser.scala 32:35]
  assign mau_3_io_mod_state_id_mod = io_mod_en ? io_mod_module_mod_state_id_mod & mod_j_3 :
    io_mod_module_mod_state_id_mod; // @[parser.scala 41:22 parser.scala 48:40 parser.scala 37:23]
  assign mau_3_io_mod_state_id = io_mod_module_mod_state_id; // @[parser.scala 37:23]
  assign mau_3_io_mod_sram_w_cs = io_mod_module_mod_sram_w_cs; // @[parser.scala 37:23]
  assign mau_3_io_mod_sram_w_en = io_mod_en ? io_mod_module_mod_sram_w_en & mod_j_3 : io_mod_module_mod_sram_w_en; // @[parser.scala 41:22 parser.scala 47:40 parser.scala 37:23]
  assign mau_3_io_mod_sram_w_addr = io_mod_module_mod_sram_w_addr; // @[parser.scala 37:23]
  assign mau_3_io_mod_sram_w_data = io_mod_module_mod_sram_w_data; // @[parser.scala 37:23]
  always @(posedge clock) begin
    if (io_mod_en) begin // @[parser.scala 41:22]
      if (io_mod_last_mau_id_mod) begin // @[parser.scala 42:39]
        last_mau_id <= {{1'd0}, io_mod_last_mau_id}; // @[parser.scala 43:25]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  last_mau_id = _RAND_0[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
