module IPSA(
  input        clock,
  input  [7:0] io_pipe_phv_in_data_0,
  input  [7:0] io_pipe_phv_in_data_1,
  input  [7:0] io_pipe_phv_in_data_2,
  input  [7:0] io_pipe_phv_in_data_3,
  input  [7:0] io_pipe_phv_in_data_4,
  input  [7:0] io_pipe_phv_in_data_5,
  input  [7:0] io_pipe_phv_in_data_6,
  input  [7:0] io_pipe_phv_in_data_7,
  input  [7:0] io_pipe_phv_in_data_8,
  input  [7:0] io_pipe_phv_in_data_9,
  input  [7:0] io_pipe_phv_in_data_10,
  input  [7:0] io_pipe_phv_in_data_11,
  input  [7:0] io_pipe_phv_in_data_12,
  input  [7:0] io_pipe_phv_in_data_13,
  input  [7:0] io_pipe_phv_in_data_14,
  input  [7:0] io_pipe_phv_in_data_15,
  input  [7:0] io_pipe_phv_in_data_16,
  input  [7:0] io_pipe_phv_in_data_17,
  input  [7:0] io_pipe_phv_in_data_18,
  input  [7:0] io_pipe_phv_in_data_19,
  input  [7:0] io_pipe_phv_in_data_20,
  input  [7:0] io_pipe_phv_in_data_21,
  input  [7:0] io_pipe_phv_in_data_22,
  input  [7:0] io_pipe_phv_in_data_23,
  input  [7:0] io_pipe_phv_in_data_24,
  input  [7:0] io_pipe_phv_in_data_25,
  input  [7:0] io_pipe_phv_in_data_26,
  input  [7:0] io_pipe_phv_in_data_27,
  input  [7:0] io_pipe_phv_in_data_28,
  input  [7:0] io_pipe_phv_in_data_29,
  input  [7:0] io_pipe_phv_in_data_30,
  input  [7:0] io_pipe_phv_in_data_31,
  input  [7:0] io_pipe_phv_in_data_32,
  input  [7:0] io_pipe_phv_in_data_33,
  input  [7:0] io_pipe_phv_in_data_34,
  input  [7:0] io_pipe_phv_in_data_35,
  input  [7:0] io_pipe_phv_in_data_36,
  input  [7:0] io_pipe_phv_in_data_37,
  input  [7:0] io_pipe_phv_in_data_38,
  input  [7:0] io_pipe_phv_in_data_39,
  input  [7:0] io_pipe_phv_in_data_40,
  input  [7:0] io_pipe_phv_in_data_41,
  input  [7:0] io_pipe_phv_in_data_42,
  input  [7:0] io_pipe_phv_in_data_43,
  input  [7:0] io_pipe_phv_in_data_44,
  input  [7:0] io_pipe_phv_in_data_45,
  input  [7:0] io_pipe_phv_in_data_46,
  input  [7:0] io_pipe_phv_in_data_47,
  input  [7:0] io_pipe_phv_in_data_48,
  input  [7:0] io_pipe_phv_in_data_49,
  input  [7:0] io_pipe_phv_in_data_50,
  input  [7:0] io_pipe_phv_in_data_51,
  input  [7:0] io_pipe_phv_in_data_52,
  input  [7:0] io_pipe_phv_in_data_53,
  input  [7:0] io_pipe_phv_in_data_54,
  input  [7:0] io_pipe_phv_in_data_55,
  input  [7:0] io_pipe_phv_in_data_56,
  input  [7:0] io_pipe_phv_in_data_57,
  input  [7:0] io_pipe_phv_in_data_58,
  input  [7:0] io_pipe_phv_in_data_59,
  input  [7:0] io_pipe_phv_in_data_60,
  input  [7:0] io_pipe_phv_in_data_61,
  input  [7:0] io_pipe_phv_in_data_62,
  input  [7:0] io_pipe_phv_in_data_63,
  input  [7:0] io_pipe_phv_in_data_64,
  input  [7:0] io_pipe_phv_in_data_65,
  input  [7:0] io_pipe_phv_in_data_66,
  input  [7:0] io_pipe_phv_in_data_67,
  input  [7:0] io_pipe_phv_in_data_68,
  input  [7:0] io_pipe_phv_in_data_69,
  input  [7:0] io_pipe_phv_in_data_70,
  input  [7:0] io_pipe_phv_in_data_71,
  input  [7:0] io_pipe_phv_in_data_72,
  input  [7:0] io_pipe_phv_in_data_73,
  input  [7:0] io_pipe_phv_in_data_74,
  input  [7:0] io_pipe_phv_in_data_75,
  input  [7:0] io_pipe_phv_in_data_76,
  input  [7:0] io_pipe_phv_in_data_77,
  input  [7:0] io_pipe_phv_in_data_78,
  input  [7:0] io_pipe_phv_in_data_79,
  input  [7:0] io_pipe_phv_in_data_80,
  input  [7:0] io_pipe_phv_in_data_81,
  input  [7:0] io_pipe_phv_in_data_82,
  input  [7:0] io_pipe_phv_in_data_83,
  input  [7:0] io_pipe_phv_in_data_84,
  input  [7:0] io_pipe_phv_in_data_85,
  input  [7:0] io_pipe_phv_in_data_86,
  input  [7:0] io_pipe_phv_in_data_87,
  input  [7:0] io_pipe_phv_in_data_88,
  input  [7:0] io_pipe_phv_in_data_89,
  input  [7:0] io_pipe_phv_in_data_90,
  input  [7:0] io_pipe_phv_in_data_91,
  input  [7:0] io_pipe_phv_in_data_92,
  input  [7:0] io_pipe_phv_in_data_93,
  input  [7:0] io_pipe_phv_in_data_94,
  input  [7:0] io_pipe_phv_in_data_95,
  input  [7:0] io_pipe_phv_in_data_96,
  input  [7:0] io_pipe_phv_in_data_97,
  input  [7:0] io_pipe_phv_in_data_98,
  input  [7:0] io_pipe_phv_in_data_99,
  input  [7:0] io_pipe_phv_in_data_100,
  input  [7:0] io_pipe_phv_in_data_101,
  input  [7:0] io_pipe_phv_in_data_102,
  input  [7:0] io_pipe_phv_in_data_103,
  input  [7:0] io_pipe_phv_in_data_104,
  input  [7:0] io_pipe_phv_in_data_105,
  input  [7:0] io_pipe_phv_in_data_106,
  input  [7:0] io_pipe_phv_in_data_107,
  input  [7:0] io_pipe_phv_in_data_108,
  input  [7:0] io_pipe_phv_in_data_109,
  input  [7:0] io_pipe_phv_in_data_110,
  input  [7:0] io_pipe_phv_in_data_111,
  input  [7:0] io_pipe_phv_in_data_112,
  input  [7:0] io_pipe_phv_in_data_113,
  input  [7:0] io_pipe_phv_in_data_114,
  input  [7:0] io_pipe_phv_in_data_115,
  input  [7:0] io_pipe_phv_in_data_116,
  input  [7:0] io_pipe_phv_in_data_117,
  input  [7:0] io_pipe_phv_in_data_118,
  input  [7:0] io_pipe_phv_in_data_119,
  input  [7:0] io_pipe_phv_in_data_120,
  input  [7:0] io_pipe_phv_in_data_121,
  input  [7:0] io_pipe_phv_in_data_122,
  input  [7:0] io_pipe_phv_in_data_123,
  input  [7:0] io_pipe_phv_in_data_124,
  input  [7:0] io_pipe_phv_in_data_125,
  input  [7:0] io_pipe_phv_in_data_126,
  input  [7:0] io_pipe_phv_in_data_127,
  input        io_pipe_phv_in_valid,
  input        io_pipe_phv_in_last,
  output [7:0] io_pipe_phv_out_data_0,
  output [7:0] io_pipe_phv_out_data_1,
  output [7:0] io_pipe_phv_out_data_2,
  output [7:0] io_pipe_phv_out_data_3,
  output [7:0] io_pipe_phv_out_data_4,
  output [7:0] io_pipe_phv_out_data_5,
  output [7:0] io_pipe_phv_out_data_6,
  output [7:0] io_pipe_phv_out_data_7,
  output [7:0] io_pipe_phv_out_data_8,
  output [7:0] io_pipe_phv_out_data_9,
  output [7:0] io_pipe_phv_out_data_10,
  output [7:0] io_pipe_phv_out_data_11,
  output [7:0] io_pipe_phv_out_data_12,
  output [7:0] io_pipe_phv_out_data_13,
  output [7:0] io_pipe_phv_out_data_14,
  output [7:0] io_pipe_phv_out_data_15,
  output [7:0] io_pipe_phv_out_data_16,
  output [7:0] io_pipe_phv_out_data_17,
  output [7:0] io_pipe_phv_out_data_18,
  output [7:0] io_pipe_phv_out_data_19,
  output [7:0] io_pipe_phv_out_data_20,
  output [7:0] io_pipe_phv_out_data_21,
  output [7:0] io_pipe_phv_out_data_22,
  output [7:0] io_pipe_phv_out_data_23,
  output [7:0] io_pipe_phv_out_data_24,
  output [7:0] io_pipe_phv_out_data_25,
  output [7:0] io_pipe_phv_out_data_26,
  output [7:0] io_pipe_phv_out_data_27,
  output [7:0] io_pipe_phv_out_data_28,
  output [7:0] io_pipe_phv_out_data_29,
  output [7:0] io_pipe_phv_out_data_30,
  output [7:0] io_pipe_phv_out_data_31,
  output [7:0] io_pipe_phv_out_data_32,
  output [7:0] io_pipe_phv_out_data_33,
  output [7:0] io_pipe_phv_out_data_34,
  output [7:0] io_pipe_phv_out_data_35,
  output [7:0] io_pipe_phv_out_data_36,
  output [7:0] io_pipe_phv_out_data_37,
  output [7:0] io_pipe_phv_out_data_38,
  output [7:0] io_pipe_phv_out_data_39,
  output [7:0] io_pipe_phv_out_data_40,
  output [7:0] io_pipe_phv_out_data_41,
  output [7:0] io_pipe_phv_out_data_42,
  output [7:0] io_pipe_phv_out_data_43,
  output [7:0] io_pipe_phv_out_data_44,
  output [7:0] io_pipe_phv_out_data_45,
  output [7:0] io_pipe_phv_out_data_46,
  output [7:0] io_pipe_phv_out_data_47,
  output [7:0] io_pipe_phv_out_data_48,
  output [7:0] io_pipe_phv_out_data_49,
  output [7:0] io_pipe_phv_out_data_50,
  output [7:0] io_pipe_phv_out_data_51,
  output [7:0] io_pipe_phv_out_data_52,
  output [7:0] io_pipe_phv_out_data_53,
  output [7:0] io_pipe_phv_out_data_54,
  output [7:0] io_pipe_phv_out_data_55,
  output [7:0] io_pipe_phv_out_data_56,
  output [7:0] io_pipe_phv_out_data_57,
  output [7:0] io_pipe_phv_out_data_58,
  output [7:0] io_pipe_phv_out_data_59,
  output [7:0] io_pipe_phv_out_data_60,
  output [7:0] io_pipe_phv_out_data_61,
  output [7:0] io_pipe_phv_out_data_62,
  output [7:0] io_pipe_phv_out_data_63,
  output [7:0] io_pipe_phv_out_data_64,
  output [7:0] io_pipe_phv_out_data_65,
  output [7:0] io_pipe_phv_out_data_66,
  output [7:0] io_pipe_phv_out_data_67,
  output [7:0] io_pipe_phv_out_data_68,
  output [7:0] io_pipe_phv_out_data_69,
  output [7:0] io_pipe_phv_out_data_70,
  output [7:0] io_pipe_phv_out_data_71,
  output [7:0] io_pipe_phv_out_data_72,
  output [7:0] io_pipe_phv_out_data_73,
  output [7:0] io_pipe_phv_out_data_74,
  output [7:0] io_pipe_phv_out_data_75,
  output [7:0] io_pipe_phv_out_data_76,
  output [7:0] io_pipe_phv_out_data_77,
  output [7:0] io_pipe_phv_out_data_78,
  output [7:0] io_pipe_phv_out_data_79,
  output [7:0] io_pipe_phv_out_data_80,
  output [7:0] io_pipe_phv_out_data_81,
  output [7:0] io_pipe_phv_out_data_82,
  output [7:0] io_pipe_phv_out_data_83,
  output [7:0] io_pipe_phv_out_data_84,
  output [7:0] io_pipe_phv_out_data_85,
  output [7:0] io_pipe_phv_out_data_86,
  output [7:0] io_pipe_phv_out_data_87,
  output [7:0] io_pipe_phv_out_data_88,
  output [7:0] io_pipe_phv_out_data_89,
  output [7:0] io_pipe_phv_out_data_90,
  output [7:0] io_pipe_phv_out_data_91,
  output [7:0] io_pipe_phv_out_data_92,
  output [7:0] io_pipe_phv_out_data_93,
  output [7:0] io_pipe_phv_out_data_94,
  output [7:0] io_pipe_phv_out_data_95,
  output [7:0] io_pipe_phv_out_data_96,
  output [7:0] io_pipe_phv_out_data_97,
  output [7:0] io_pipe_phv_out_data_98,
  output [7:0] io_pipe_phv_out_data_99,
  output [7:0] io_pipe_phv_out_data_100,
  output [7:0] io_pipe_phv_out_data_101,
  output [7:0] io_pipe_phv_out_data_102,
  output [7:0] io_pipe_phv_out_data_103,
  output [7:0] io_pipe_phv_out_data_104,
  output [7:0] io_pipe_phv_out_data_105,
  output [7:0] io_pipe_phv_out_data_106,
  output [7:0] io_pipe_phv_out_data_107,
  output [7:0] io_pipe_phv_out_data_108,
  output [7:0] io_pipe_phv_out_data_109,
  output [7:0] io_pipe_phv_out_data_110,
  output [7:0] io_pipe_phv_out_data_111,
  output [7:0] io_pipe_phv_out_data_112,
  output [7:0] io_pipe_phv_out_data_113,
  output [7:0] io_pipe_phv_out_data_114,
  output [7:0] io_pipe_phv_out_data_115,
  output [7:0] io_pipe_phv_out_data_116,
  output [7:0] io_pipe_phv_out_data_117,
  output [7:0] io_pipe_phv_out_data_118,
  output [7:0] io_pipe_phv_out_data_119,
  output [7:0] io_pipe_phv_out_data_120,
  output [7:0] io_pipe_phv_out_data_121,
  output [7:0] io_pipe_phv_out_data_122,
  output [7:0] io_pipe_phv_out_data_123,
  output [7:0] io_pipe_phv_out_data_124,
  output [7:0] io_pipe_phv_out_data_125,
  output [7:0] io_pipe_phv_out_data_126,
  output [7:0] io_pipe_phv_out_data_127,
  output       io_pipe_phv_out_valid,
  output       io_pipe_phv_out_last
);
  wire  proc_0_clock; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_0; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_1; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_2; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_3; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_4; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_5; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_6; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_7; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_8; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_9; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_10; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_11; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_12; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_13; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_14; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_16; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_17; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_18; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_19; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_20; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_21; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_22; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_23; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_24; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_25; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_26; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_27; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_28; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_29; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_30; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_31; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_32; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_33; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_34; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_35; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_36; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_37; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_38; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_39; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_40; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_41; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_42; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_43; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_44; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_45; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_46; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_47; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_48; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_49; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_50; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_51; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_52; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_53; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_54; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_55; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_56; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_57; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_58; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_59; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_60; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_61; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_62; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_63; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_64; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_65; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_66; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_67; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_68; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_69; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_70; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_71; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_72; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_73; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_74; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_75; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_76; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_77; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_78; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_79; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_80; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_81; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_82; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_83; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_84; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_85; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_86; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_87; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_88; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_89; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_90; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_91; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_92; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_93; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_94; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_95; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_96; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_97; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_98; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_99; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_100; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_101; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_102; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_103; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_104; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_105; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_106; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_107; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_108; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_109; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_110; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_111; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_112; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_113; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_114; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_115; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_116; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_117; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_118; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_119; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_120; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_121; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_122; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_123; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_124; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_125; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_126; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_127; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_128; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_129; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_130; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_131; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_132; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_133; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_134; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_135; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_136; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_137; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_138; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_139; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_140; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_141; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_142; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_143; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_144; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_145; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_146; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_147; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_148; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_149; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_150; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_151; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_152; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_153; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_154; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_155; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_156; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_157; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_158; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_159; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_in_header_0; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_in_header_1; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_in_header_2; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_in_header_3; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_in_header_4; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_in_header_5; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_in_header_6; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_in_header_7; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_in_header_8; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_in_header_9; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_in_header_10; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_in_header_11; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_in_header_12; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_in_header_13; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_in_header_14; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_in_header_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_parse_current_state; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_parse_current_offset; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_in_parse_transition_field; // @[ipsa.scala 56:25]
  wire [3:0] proc_0_io_pipe_phv_in_next_processor_id; // @[ipsa.scala 56:25]
  wire  proc_0_io_pipe_phv_in_next_config_id; // @[ipsa.scala 56:25]
  wire  proc_0_io_pipe_phv_in_is_valid_processor; // @[ipsa.scala 56:25]
  wire  proc_0_io_pipe_phv_in_valid; // @[ipsa.scala 56:25]
  wire  proc_0_io_pipe_phv_in_last; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_0; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_1; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_2; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_3; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_4; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_5; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_6; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_7; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_8; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_9; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_10; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_11; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_12; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_13; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_14; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_16; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_17; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_18; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_19; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_20; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_21; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_22; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_23; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_24; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_25; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_26; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_27; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_28; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_29; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_30; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_31; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_32; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_33; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_34; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_35; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_36; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_37; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_38; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_39; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_40; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_41; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_42; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_43; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_44; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_45; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_46; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_47; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_48; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_49; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_50; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_51; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_52; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_53; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_54; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_55; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_56; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_57; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_58; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_59; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_60; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_61; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_62; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_63; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_64; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_65; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_66; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_67; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_68; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_69; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_70; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_71; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_72; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_73; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_74; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_75; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_76; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_77; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_78; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_79; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_80; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_81; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_82; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_83; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_84; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_85; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_86; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_87; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_88; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_89; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_90; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_91; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_92; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_93; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_94; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_95; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_96; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_97; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_98; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_99; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_100; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_101; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_102; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_103; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_104; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_105; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_106; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_107; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_108; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_109; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_110; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_111; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_112; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_113; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_114; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_115; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_116; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_117; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_118; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_119; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_120; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_121; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_122; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_123; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_124; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_125; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_126; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_127; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_128; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_129; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_130; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_131; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_132; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_133; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_134; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_135; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_136; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_137; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_138; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_139; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_140; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_141; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_142; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_143; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_144; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_145; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_146; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_147; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_148; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_149; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_150; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_151; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_152; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_153; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_154; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_155; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_156; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_157; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_158; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_159; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_out_header_0; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_out_header_1; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_out_header_2; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_out_header_3; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_out_header_4; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_out_header_5; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_out_header_6; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_out_header_7; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_out_header_8; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_out_header_9; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_out_header_10; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_out_header_11; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_out_header_12; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_out_header_13; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_out_header_14; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_out_header_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 56:25]
  wire [3:0] proc_0_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 56:25]
  wire  proc_0_io_pipe_phv_out_next_config_id; // @[ipsa.scala 56:25]
  wire  proc_0_io_pipe_phv_out_valid; // @[ipsa.scala 56:25]
  wire  proc_0_io_pipe_phv_out_last; // @[ipsa.scala 56:25]
  wire  proc_1_clock; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_0; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_1; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_2; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_3; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_4; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_5; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_6; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_7; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_8; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_9; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_10; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_11; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_12; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_13; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_14; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_16; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_17; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_18; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_19; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_20; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_21; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_22; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_23; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_24; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_25; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_26; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_27; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_28; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_29; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_30; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_31; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_32; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_33; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_34; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_35; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_36; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_37; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_38; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_39; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_40; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_41; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_42; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_43; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_44; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_45; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_46; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_47; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_48; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_49; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_50; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_51; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_52; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_53; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_54; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_55; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_56; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_57; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_58; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_59; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_60; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_61; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_62; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_63; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_64; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_65; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_66; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_67; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_68; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_69; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_70; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_71; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_72; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_73; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_74; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_75; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_76; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_77; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_78; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_79; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_80; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_81; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_82; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_83; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_84; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_85; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_86; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_87; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_88; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_89; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_90; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_91; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_92; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_93; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_94; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_95; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_96; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_97; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_98; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_99; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_100; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_101; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_102; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_103; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_104; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_105; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_106; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_107; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_108; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_109; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_110; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_111; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_112; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_113; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_114; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_115; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_116; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_117; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_118; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_119; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_120; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_121; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_122; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_123; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_124; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_125; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_126; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_127; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_128; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_129; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_130; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_131; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_132; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_133; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_134; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_135; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_136; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_137; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_138; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_139; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_140; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_141; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_142; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_143; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_144; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_145; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_146; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_147; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_148; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_149; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_150; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_151; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_152; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_153; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_154; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_155; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_156; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_157; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_158; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_159; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_in_header_0; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_in_header_1; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_in_header_2; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_in_header_3; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_in_header_4; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_in_header_5; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_in_header_6; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_in_header_7; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_in_header_8; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_in_header_9; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_in_header_10; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_in_header_11; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_in_header_12; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_in_header_13; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_in_header_14; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_in_header_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_parse_current_state; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_parse_current_offset; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_in_parse_transition_field; // @[ipsa.scala 56:25]
  wire [3:0] proc_1_io_pipe_phv_in_next_processor_id; // @[ipsa.scala 56:25]
  wire  proc_1_io_pipe_phv_in_next_config_id; // @[ipsa.scala 56:25]
  wire  proc_1_io_pipe_phv_in_is_valid_processor; // @[ipsa.scala 56:25]
  wire  proc_1_io_pipe_phv_in_valid; // @[ipsa.scala 56:25]
  wire  proc_1_io_pipe_phv_in_last; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_0; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_1; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_2; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_3; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_4; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_5; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_6; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_7; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_8; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_9; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_10; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_11; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_12; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_13; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_14; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_16; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_17; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_18; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_19; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_20; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_21; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_22; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_23; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_24; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_25; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_26; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_27; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_28; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_29; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_30; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_31; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_32; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_33; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_34; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_35; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_36; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_37; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_38; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_39; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_40; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_41; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_42; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_43; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_44; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_45; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_46; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_47; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_48; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_49; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_50; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_51; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_52; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_53; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_54; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_55; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_56; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_57; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_58; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_59; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_60; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_61; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_62; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_63; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_64; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_65; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_66; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_67; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_68; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_69; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_70; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_71; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_72; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_73; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_74; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_75; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_76; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_77; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_78; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_79; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_80; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_81; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_82; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_83; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_84; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_85; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_86; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_87; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_88; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_89; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_90; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_91; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_92; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_93; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_94; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_95; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_96; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_97; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_98; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_99; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_100; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_101; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_102; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_103; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_104; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_105; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_106; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_107; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_108; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_109; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_110; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_111; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_112; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_113; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_114; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_115; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_116; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_117; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_118; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_119; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_120; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_121; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_122; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_123; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_124; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_125; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_126; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_127; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_128; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_129; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_130; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_131; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_132; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_133; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_134; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_135; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_136; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_137; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_138; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_139; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_140; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_141; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_142; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_143; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_144; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_145; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_146; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_147; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_148; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_149; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_150; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_151; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_152; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_153; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_154; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_155; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_156; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_157; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_158; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_159; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_out_header_0; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_out_header_1; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_out_header_2; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_out_header_3; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_out_header_4; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_out_header_5; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_out_header_6; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_out_header_7; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_out_header_8; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_out_header_9; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_out_header_10; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_out_header_11; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_out_header_12; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_out_header_13; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_out_header_14; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_out_header_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 56:25]
  wire [3:0] proc_1_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 56:25]
  wire  proc_1_io_pipe_phv_out_next_config_id; // @[ipsa.scala 56:25]
  wire  proc_1_io_pipe_phv_out_valid; // @[ipsa.scala 56:25]
  wire  proc_1_io_pipe_phv_out_last; // @[ipsa.scala 56:25]
  wire  proc_2_clock; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_0; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_1; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_2; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_3; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_4; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_5; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_6; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_7; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_8; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_9; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_10; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_11; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_12; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_13; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_14; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_16; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_17; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_18; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_19; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_20; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_21; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_22; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_23; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_24; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_25; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_26; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_27; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_28; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_29; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_30; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_31; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_32; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_33; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_34; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_35; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_36; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_37; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_38; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_39; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_40; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_41; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_42; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_43; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_44; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_45; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_46; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_47; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_48; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_49; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_50; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_51; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_52; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_53; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_54; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_55; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_56; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_57; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_58; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_59; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_60; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_61; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_62; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_63; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_64; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_65; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_66; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_67; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_68; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_69; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_70; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_71; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_72; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_73; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_74; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_75; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_76; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_77; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_78; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_79; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_80; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_81; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_82; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_83; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_84; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_85; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_86; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_87; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_88; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_89; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_90; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_91; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_92; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_93; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_94; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_95; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_96; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_97; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_98; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_99; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_100; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_101; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_102; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_103; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_104; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_105; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_106; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_107; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_108; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_109; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_110; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_111; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_112; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_113; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_114; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_115; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_116; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_117; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_118; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_119; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_120; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_121; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_122; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_123; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_124; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_125; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_126; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_127; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_128; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_129; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_130; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_131; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_132; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_133; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_134; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_135; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_136; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_137; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_138; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_139; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_140; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_141; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_142; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_143; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_144; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_145; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_146; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_147; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_148; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_149; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_150; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_151; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_152; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_153; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_154; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_155; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_156; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_157; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_158; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_159; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_in_header_0; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_in_header_1; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_in_header_2; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_in_header_3; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_in_header_4; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_in_header_5; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_in_header_6; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_in_header_7; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_in_header_8; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_in_header_9; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_in_header_10; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_in_header_11; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_in_header_12; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_in_header_13; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_in_header_14; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_in_header_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_parse_current_state; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_parse_current_offset; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_in_parse_transition_field; // @[ipsa.scala 56:25]
  wire [3:0] proc_2_io_pipe_phv_in_next_processor_id; // @[ipsa.scala 56:25]
  wire  proc_2_io_pipe_phv_in_next_config_id; // @[ipsa.scala 56:25]
  wire  proc_2_io_pipe_phv_in_is_valid_processor; // @[ipsa.scala 56:25]
  wire  proc_2_io_pipe_phv_in_valid; // @[ipsa.scala 56:25]
  wire  proc_2_io_pipe_phv_in_last; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_0; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_1; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_2; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_3; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_4; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_5; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_6; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_7; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_8; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_9; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_10; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_11; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_12; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_13; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_14; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_16; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_17; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_18; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_19; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_20; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_21; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_22; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_23; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_24; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_25; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_26; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_27; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_28; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_29; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_30; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_31; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_32; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_33; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_34; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_35; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_36; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_37; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_38; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_39; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_40; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_41; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_42; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_43; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_44; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_45; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_46; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_47; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_48; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_49; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_50; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_51; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_52; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_53; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_54; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_55; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_56; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_57; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_58; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_59; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_60; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_61; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_62; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_63; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_64; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_65; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_66; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_67; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_68; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_69; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_70; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_71; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_72; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_73; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_74; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_75; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_76; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_77; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_78; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_79; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_80; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_81; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_82; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_83; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_84; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_85; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_86; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_87; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_88; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_89; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_90; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_91; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_92; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_93; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_94; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_95; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_96; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_97; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_98; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_99; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_100; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_101; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_102; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_103; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_104; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_105; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_106; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_107; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_108; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_109; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_110; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_111; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_112; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_113; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_114; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_115; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_116; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_117; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_118; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_119; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_120; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_121; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_122; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_123; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_124; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_125; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_126; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_127; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_128; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_129; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_130; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_131; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_132; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_133; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_134; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_135; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_136; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_137; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_138; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_139; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_140; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_141; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_142; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_143; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_144; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_145; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_146; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_147; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_148; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_149; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_150; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_151; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_152; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_153; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_154; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_155; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_156; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_157; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_158; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_159; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_out_header_0; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_out_header_1; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_out_header_2; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_out_header_3; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_out_header_4; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_out_header_5; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_out_header_6; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_out_header_7; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_out_header_8; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_out_header_9; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_out_header_10; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_out_header_11; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_out_header_12; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_out_header_13; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_out_header_14; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_out_header_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 56:25]
  wire [3:0] proc_2_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 56:25]
  wire  proc_2_io_pipe_phv_out_next_config_id; // @[ipsa.scala 56:25]
  wire  proc_2_io_pipe_phv_out_valid; // @[ipsa.scala 56:25]
  wire  proc_2_io_pipe_phv_out_last; // @[ipsa.scala 56:25]
  wire  proc_3_clock; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_0; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_1; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_2; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_3; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_4; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_5; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_6; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_7; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_8; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_9; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_10; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_11; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_12; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_13; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_14; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_16; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_17; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_18; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_19; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_20; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_21; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_22; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_23; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_24; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_25; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_26; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_27; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_28; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_29; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_30; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_31; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_32; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_33; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_34; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_35; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_36; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_37; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_38; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_39; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_40; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_41; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_42; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_43; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_44; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_45; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_46; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_47; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_48; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_49; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_50; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_51; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_52; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_53; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_54; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_55; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_56; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_57; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_58; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_59; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_60; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_61; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_62; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_63; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_64; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_65; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_66; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_67; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_68; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_69; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_70; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_71; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_72; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_73; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_74; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_75; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_76; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_77; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_78; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_79; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_80; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_81; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_82; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_83; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_84; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_85; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_86; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_87; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_88; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_89; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_90; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_91; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_92; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_93; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_94; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_95; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_96; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_97; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_98; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_99; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_100; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_101; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_102; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_103; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_104; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_105; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_106; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_107; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_108; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_109; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_110; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_111; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_112; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_113; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_114; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_115; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_116; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_117; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_118; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_119; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_120; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_121; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_122; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_123; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_124; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_125; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_126; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_127; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_128; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_129; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_130; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_131; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_132; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_133; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_134; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_135; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_136; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_137; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_138; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_139; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_140; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_141; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_142; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_143; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_144; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_145; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_146; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_147; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_148; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_149; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_150; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_151; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_152; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_153; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_154; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_155; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_156; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_157; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_158; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_159; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_in_header_0; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_in_header_1; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_in_header_2; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_in_header_3; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_in_header_4; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_in_header_5; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_in_header_6; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_in_header_7; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_in_header_8; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_in_header_9; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_in_header_10; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_in_header_11; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_in_header_12; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_in_header_13; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_in_header_14; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_in_header_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_parse_current_state; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_parse_current_offset; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_in_parse_transition_field; // @[ipsa.scala 56:25]
  wire [3:0] proc_3_io_pipe_phv_in_next_processor_id; // @[ipsa.scala 56:25]
  wire  proc_3_io_pipe_phv_in_next_config_id; // @[ipsa.scala 56:25]
  wire  proc_3_io_pipe_phv_in_is_valid_processor; // @[ipsa.scala 56:25]
  wire  proc_3_io_pipe_phv_in_valid; // @[ipsa.scala 56:25]
  wire  proc_3_io_pipe_phv_in_last; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_0; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_1; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_2; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_3; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_4; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_5; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_6; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_7; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_8; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_9; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_10; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_11; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_12; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_13; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_14; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_16; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_17; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_18; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_19; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_20; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_21; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_22; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_23; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_24; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_25; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_26; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_27; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_28; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_29; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_30; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_31; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_32; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_33; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_34; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_35; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_36; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_37; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_38; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_39; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_40; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_41; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_42; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_43; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_44; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_45; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_46; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_47; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_48; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_49; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_50; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_51; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_52; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_53; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_54; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_55; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_56; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_57; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_58; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_59; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_60; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_61; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_62; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_63; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_64; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_65; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_66; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_67; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_68; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_69; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_70; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_71; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_72; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_73; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_74; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_75; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_76; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_77; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_78; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_79; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_80; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_81; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_82; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_83; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_84; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_85; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_86; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_87; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_88; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_89; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_90; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_91; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_92; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_93; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_94; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_95; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_96; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_97; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_98; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_99; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_100; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_101; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_102; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_103; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_104; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_105; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_106; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_107; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_108; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_109; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_110; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_111; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_112; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_113; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_114; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_115; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_116; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_117; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_118; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_119; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_120; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_121; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_122; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_123; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_124; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_125; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_126; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_127; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_128; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_129; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_130; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_131; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_132; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_133; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_134; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_135; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_136; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_137; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_138; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_139; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_140; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_141; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_142; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_143; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_144; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_145; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_146; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_147; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_148; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_149; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_150; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_151; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_152; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_153; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_154; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_155; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_156; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_157; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_158; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_159; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_out_header_0; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_out_header_1; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_out_header_2; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_out_header_3; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_out_header_4; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_out_header_5; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_out_header_6; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_out_header_7; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_out_header_8; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_out_header_9; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_out_header_10; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_out_header_11; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_out_header_12; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_out_header_13; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_out_header_14; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_out_header_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 56:25]
  wire [3:0] proc_3_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 56:25]
  wire  proc_3_io_pipe_phv_out_next_config_id; // @[ipsa.scala 56:25]
  wire  proc_3_io_pipe_phv_out_valid; // @[ipsa.scala 56:25]
  wire  proc_3_io_pipe_phv_out_last; // @[ipsa.scala 56:25]
  wire  proc_4_clock; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_0; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_1; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_2; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_3; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_4; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_5; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_6; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_7; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_8; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_9; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_10; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_11; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_12; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_13; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_14; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_16; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_17; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_18; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_19; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_20; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_21; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_22; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_23; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_24; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_25; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_26; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_27; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_28; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_29; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_30; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_31; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_32; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_33; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_34; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_35; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_36; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_37; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_38; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_39; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_40; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_41; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_42; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_43; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_44; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_45; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_46; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_47; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_48; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_49; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_50; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_51; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_52; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_53; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_54; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_55; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_56; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_57; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_58; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_59; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_60; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_61; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_62; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_63; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_64; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_65; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_66; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_67; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_68; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_69; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_70; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_71; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_72; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_73; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_74; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_75; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_76; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_77; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_78; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_79; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_80; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_81; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_82; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_83; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_84; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_85; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_86; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_87; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_88; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_89; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_90; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_91; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_92; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_93; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_94; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_95; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_96; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_97; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_98; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_99; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_100; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_101; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_102; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_103; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_104; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_105; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_106; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_107; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_108; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_109; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_110; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_111; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_112; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_113; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_114; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_115; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_116; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_117; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_118; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_119; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_120; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_121; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_122; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_123; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_124; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_125; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_126; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_127; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_128; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_129; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_130; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_131; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_132; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_133; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_134; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_135; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_136; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_137; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_138; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_139; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_140; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_141; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_142; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_143; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_144; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_145; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_146; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_147; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_148; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_149; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_150; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_151; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_152; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_153; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_154; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_155; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_156; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_157; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_158; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_159; // @[ipsa.scala 56:25]
  wire [15:0] proc_4_io_pipe_phv_in_header_0; // @[ipsa.scala 56:25]
  wire [15:0] proc_4_io_pipe_phv_in_header_1; // @[ipsa.scala 56:25]
  wire [15:0] proc_4_io_pipe_phv_in_header_2; // @[ipsa.scala 56:25]
  wire [15:0] proc_4_io_pipe_phv_in_header_3; // @[ipsa.scala 56:25]
  wire [15:0] proc_4_io_pipe_phv_in_header_4; // @[ipsa.scala 56:25]
  wire [15:0] proc_4_io_pipe_phv_in_header_5; // @[ipsa.scala 56:25]
  wire [15:0] proc_4_io_pipe_phv_in_header_6; // @[ipsa.scala 56:25]
  wire [15:0] proc_4_io_pipe_phv_in_header_7; // @[ipsa.scala 56:25]
  wire [15:0] proc_4_io_pipe_phv_in_header_8; // @[ipsa.scala 56:25]
  wire [15:0] proc_4_io_pipe_phv_in_header_9; // @[ipsa.scala 56:25]
  wire [15:0] proc_4_io_pipe_phv_in_header_10; // @[ipsa.scala 56:25]
  wire [15:0] proc_4_io_pipe_phv_in_header_11; // @[ipsa.scala 56:25]
  wire [15:0] proc_4_io_pipe_phv_in_header_12; // @[ipsa.scala 56:25]
  wire [15:0] proc_4_io_pipe_phv_in_header_13; // @[ipsa.scala 56:25]
  wire [15:0] proc_4_io_pipe_phv_in_header_14; // @[ipsa.scala 56:25]
  wire [15:0] proc_4_io_pipe_phv_in_header_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_parse_current_state; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_in_parse_current_offset; // @[ipsa.scala 56:25]
  wire [15:0] proc_4_io_pipe_phv_in_parse_transition_field; // @[ipsa.scala 56:25]
  wire [3:0] proc_4_io_pipe_phv_in_next_processor_id; // @[ipsa.scala 56:25]
  wire  proc_4_io_pipe_phv_in_next_config_id; // @[ipsa.scala 56:25]
  wire  proc_4_io_pipe_phv_in_is_valid_processor; // @[ipsa.scala 56:25]
  wire  proc_4_io_pipe_phv_in_valid; // @[ipsa.scala 56:25]
  wire  proc_4_io_pipe_phv_in_last; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_0; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_1; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_2; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_3; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_4; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_5; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_6; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_7; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_8; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_9; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_10; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_11; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_12; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_13; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_14; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_16; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_17; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_18; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_19; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_20; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_21; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_22; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_23; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_24; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_25; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_26; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_27; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_28; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_29; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_30; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_31; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_32; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_33; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_34; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_35; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_36; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_37; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_38; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_39; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_40; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_41; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_42; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_43; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_44; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_45; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_46; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_47; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_48; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_49; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_50; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_51; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_52; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_53; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_54; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_55; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_56; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_57; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_58; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_59; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_60; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_61; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_62; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_63; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_64; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_65; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_66; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_67; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_68; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_69; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_70; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_71; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_72; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_73; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_74; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_75; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_76; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_77; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_78; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_79; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_80; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_81; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_82; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_83; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_84; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_85; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_86; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_87; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_88; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_89; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_90; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_91; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_92; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_93; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_94; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_95; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_96; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_97; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_98; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_99; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_100; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_101; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_102; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_103; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_104; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_105; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_106; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_107; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_108; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_109; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_110; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_111; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_112; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_113; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_114; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_115; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_116; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_117; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_118; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_119; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_120; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_121; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_122; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_123; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_124; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_125; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_126; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_127; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_128; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_129; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_130; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_131; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_132; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_133; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_134; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_135; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_136; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_137; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_138; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_139; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_140; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_141; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_142; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_143; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_144; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_145; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_146; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_147; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_148; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_149; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_150; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_151; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_152; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_153; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_154; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_155; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_156; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_157; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_158; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_159; // @[ipsa.scala 56:25]
  wire [15:0] proc_4_io_pipe_phv_out_header_0; // @[ipsa.scala 56:25]
  wire [15:0] proc_4_io_pipe_phv_out_header_1; // @[ipsa.scala 56:25]
  wire [15:0] proc_4_io_pipe_phv_out_header_2; // @[ipsa.scala 56:25]
  wire [15:0] proc_4_io_pipe_phv_out_header_3; // @[ipsa.scala 56:25]
  wire [15:0] proc_4_io_pipe_phv_out_header_4; // @[ipsa.scala 56:25]
  wire [15:0] proc_4_io_pipe_phv_out_header_5; // @[ipsa.scala 56:25]
  wire [15:0] proc_4_io_pipe_phv_out_header_6; // @[ipsa.scala 56:25]
  wire [15:0] proc_4_io_pipe_phv_out_header_7; // @[ipsa.scala 56:25]
  wire [15:0] proc_4_io_pipe_phv_out_header_8; // @[ipsa.scala 56:25]
  wire [15:0] proc_4_io_pipe_phv_out_header_9; // @[ipsa.scala 56:25]
  wire [15:0] proc_4_io_pipe_phv_out_header_10; // @[ipsa.scala 56:25]
  wire [15:0] proc_4_io_pipe_phv_out_header_11; // @[ipsa.scala 56:25]
  wire [15:0] proc_4_io_pipe_phv_out_header_12; // @[ipsa.scala 56:25]
  wire [15:0] proc_4_io_pipe_phv_out_header_13; // @[ipsa.scala 56:25]
  wire [15:0] proc_4_io_pipe_phv_out_header_14; // @[ipsa.scala 56:25]
  wire [15:0] proc_4_io_pipe_phv_out_header_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 56:25]
  wire [7:0] proc_4_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 56:25]
  wire [15:0] proc_4_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 56:25]
  wire [3:0] proc_4_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 56:25]
  wire  proc_4_io_pipe_phv_out_next_config_id; // @[ipsa.scala 56:25]
  wire  proc_4_io_pipe_phv_out_valid; // @[ipsa.scala 56:25]
  wire  proc_4_io_pipe_phv_out_last; // @[ipsa.scala 56:25]
  wire  proc_5_clock; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_0; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_1; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_2; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_3; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_4; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_5; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_6; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_7; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_8; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_9; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_10; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_11; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_12; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_13; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_14; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_16; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_17; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_18; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_19; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_20; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_21; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_22; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_23; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_24; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_25; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_26; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_27; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_28; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_29; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_30; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_31; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_32; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_33; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_34; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_35; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_36; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_37; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_38; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_39; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_40; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_41; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_42; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_43; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_44; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_45; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_46; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_47; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_48; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_49; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_50; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_51; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_52; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_53; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_54; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_55; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_56; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_57; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_58; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_59; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_60; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_61; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_62; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_63; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_64; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_65; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_66; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_67; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_68; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_69; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_70; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_71; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_72; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_73; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_74; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_75; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_76; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_77; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_78; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_79; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_80; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_81; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_82; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_83; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_84; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_85; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_86; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_87; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_88; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_89; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_90; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_91; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_92; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_93; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_94; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_95; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_96; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_97; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_98; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_99; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_100; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_101; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_102; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_103; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_104; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_105; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_106; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_107; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_108; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_109; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_110; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_111; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_112; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_113; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_114; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_115; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_116; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_117; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_118; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_119; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_120; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_121; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_122; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_123; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_124; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_125; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_126; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_127; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_128; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_129; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_130; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_131; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_132; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_133; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_134; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_135; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_136; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_137; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_138; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_139; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_140; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_141; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_142; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_143; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_144; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_145; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_146; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_147; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_148; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_149; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_150; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_151; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_152; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_153; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_154; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_155; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_156; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_157; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_158; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_159; // @[ipsa.scala 56:25]
  wire [15:0] proc_5_io_pipe_phv_in_header_0; // @[ipsa.scala 56:25]
  wire [15:0] proc_5_io_pipe_phv_in_header_1; // @[ipsa.scala 56:25]
  wire [15:0] proc_5_io_pipe_phv_in_header_2; // @[ipsa.scala 56:25]
  wire [15:0] proc_5_io_pipe_phv_in_header_3; // @[ipsa.scala 56:25]
  wire [15:0] proc_5_io_pipe_phv_in_header_4; // @[ipsa.scala 56:25]
  wire [15:0] proc_5_io_pipe_phv_in_header_5; // @[ipsa.scala 56:25]
  wire [15:0] proc_5_io_pipe_phv_in_header_6; // @[ipsa.scala 56:25]
  wire [15:0] proc_5_io_pipe_phv_in_header_7; // @[ipsa.scala 56:25]
  wire [15:0] proc_5_io_pipe_phv_in_header_8; // @[ipsa.scala 56:25]
  wire [15:0] proc_5_io_pipe_phv_in_header_9; // @[ipsa.scala 56:25]
  wire [15:0] proc_5_io_pipe_phv_in_header_10; // @[ipsa.scala 56:25]
  wire [15:0] proc_5_io_pipe_phv_in_header_11; // @[ipsa.scala 56:25]
  wire [15:0] proc_5_io_pipe_phv_in_header_12; // @[ipsa.scala 56:25]
  wire [15:0] proc_5_io_pipe_phv_in_header_13; // @[ipsa.scala 56:25]
  wire [15:0] proc_5_io_pipe_phv_in_header_14; // @[ipsa.scala 56:25]
  wire [15:0] proc_5_io_pipe_phv_in_header_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_parse_current_state; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_in_parse_current_offset; // @[ipsa.scala 56:25]
  wire [15:0] proc_5_io_pipe_phv_in_parse_transition_field; // @[ipsa.scala 56:25]
  wire [3:0] proc_5_io_pipe_phv_in_next_processor_id; // @[ipsa.scala 56:25]
  wire  proc_5_io_pipe_phv_in_next_config_id; // @[ipsa.scala 56:25]
  wire  proc_5_io_pipe_phv_in_is_valid_processor; // @[ipsa.scala 56:25]
  wire  proc_5_io_pipe_phv_in_valid; // @[ipsa.scala 56:25]
  wire  proc_5_io_pipe_phv_in_last; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_0; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_1; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_2; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_3; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_4; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_5; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_6; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_7; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_8; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_9; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_10; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_11; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_12; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_13; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_14; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_16; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_17; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_18; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_19; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_20; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_21; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_22; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_23; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_24; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_25; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_26; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_27; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_28; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_29; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_30; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_31; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_32; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_33; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_34; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_35; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_36; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_37; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_38; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_39; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_40; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_41; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_42; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_43; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_44; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_45; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_46; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_47; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_48; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_49; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_50; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_51; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_52; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_53; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_54; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_55; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_56; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_57; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_58; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_59; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_60; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_61; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_62; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_63; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_64; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_65; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_66; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_67; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_68; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_69; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_70; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_71; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_72; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_73; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_74; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_75; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_76; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_77; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_78; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_79; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_80; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_81; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_82; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_83; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_84; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_85; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_86; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_87; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_88; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_89; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_90; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_91; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_92; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_93; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_94; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_95; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_96; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_97; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_98; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_99; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_100; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_101; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_102; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_103; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_104; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_105; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_106; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_107; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_108; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_109; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_110; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_111; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_112; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_113; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_114; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_115; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_116; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_117; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_118; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_119; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_120; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_121; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_122; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_123; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_124; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_125; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_126; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_127; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_128; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_129; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_130; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_131; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_132; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_133; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_134; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_135; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_136; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_137; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_138; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_139; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_140; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_141; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_142; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_143; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_144; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_145; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_146; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_147; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_148; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_149; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_150; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_151; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_152; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_153; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_154; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_155; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_156; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_157; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_158; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_159; // @[ipsa.scala 56:25]
  wire [15:0] proc_5_io_pipe_phv_out_header_0; // @[ipsa.scala 56:25]
  wire [15:0] proc_5_io_pipe_phv_out_header_1; // @[ipsa.scala 56:25]
  wire [15:0] proc_5_io_pipe_phv_out_header_2; // @[ipsa.scala 56:25]
  wire [15:0] proc_5_io_pipe_phv_out_header_3; // @[ipsa.scala 56:25]
  wire [15:0] proc_5_io_pipe_phv_out_header_4; // @[ipsa.scala 56:25]
  wire [15:0] proc_5_io_pipe_phv_out_header_5; // @[ipsa.scala 56:25]
  wire [15:0] proc_5_io_pipe_phv_out_header_6; // @[ipsa.scala 56:25]
  wire [15:0] proc_5_io_pipe_phv_out_header_7; // @[ipsa.scala 56:25]
  wire [15:0] proc_5_io_pipe_phv_out_header_8; // @[ipsa.scala 56:25]
  wire [15:0] proc_5_io_pipe_phv_out_header_9; // @[ipsa.scala 56:25]
  wire [15:0] proc_5_io_pipe_phv_out_header_10; // @[ipsa.scala 56:25]
  wire [15:0] proc_5_io_pipe_phv_out_header_11; // @[ipsa.scala 56:25]
  wire [15:0] proc_5_io_pipe_phv_out_header_12; // @[ipsa.scala 56:25]
  wire [15:0] proc_5_io_pipe_phv_out_header_13; // @[ipsa.scala 56:25]
  wire [15:0] proc_5_io_pipe_phv_out_header_14; // @[ipsa.scala 56:25]
  wire [15:0] proc_5_io_pipe_phv_out_header_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 56:25]
  wire [7:0] proc_5_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 56:25]
  wire [15:0] proc_5_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 56:25]
  wire [3:0] proc_5_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 56:25]
  wire  proc_5_io_pipe_phv_out_next_config_id; // @[ipsa.scala 56:25]
  wire  proc_5_io_pipe_phv_out_valid; // @[ipsa.scala 56:25]
  wire  proc_5_io_pipe_phv_out_last; // @[ipsa.scala 56:25]
  wire  proc_6_clock; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_0; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_1; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_2; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_3; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_4; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_5; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_6; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_7; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_8; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_9; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_10; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_11; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_12; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_13; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_14; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_16; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_17; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_18; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_19; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_20; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_21; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_22; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_23; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_24; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_25; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_26; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_27; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_28; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_29; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_30; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_31; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_32; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_33; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_34; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_35; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_36; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_37; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_38; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_39; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_40; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_41; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_42; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_43; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_44; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_45; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_46; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_47; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_48; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_49; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_50; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_51; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_52; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_53; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_54; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_55; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_56; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_57; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_58; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_59; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_60; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_61; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_62; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_63; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_64; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_65; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_66; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_67; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_68; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_69; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_70; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_71; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_72; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_73; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_74; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_75; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_76; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_77; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_78; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_79; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_80; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_81; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_82; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_83; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_84; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_85; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_86; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_87; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_88; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_89; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_90; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_91; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_92; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_93; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_94; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_95; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_96; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_97; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_98; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_99; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_100; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_101; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_102; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_103; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_104; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_105; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_106; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_107; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_108; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_109; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_110; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_111; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_112; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_113; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_114; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_115; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_116; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_117; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_118; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_119; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_120; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_121; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_122; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_123; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_124; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_125; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_126; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_127; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_128; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_129; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_130; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_131; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_132; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_133; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_134; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_135; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_136; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_137; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_138; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_139; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_140; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_141; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_142; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_143; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_144; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_145; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_146; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_147; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_148; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_149; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_150; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_151; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_152; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_153; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_154; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_155; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_156; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_157; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_158; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_159; // @[ipsa.scala 56:25]
  wire [15:0] proc_6_io_pipe_phv_in_header_0; // @[ipsa.scala 56:25]
  wire [15:0] proc_6_io_pipe_phv_in_header_1; // @[ipsa.scala 56:25]
  wire [15:0] proc_6_io_pipe_phv_in_header_2; // @[ipsa.scala 56:25]
  wire [15:0] proc_6_io_pipe_phv_in_header_3; // @[ipsa.scala 56:25]
  wire [15:0] proc_6_io_pipe_phv_in_header_4; // @[ipsa.scala 56:25]
  wire [15:0] proc_6_io_pipe_phv_in_header_5; // @[ipsa.scala 56:25]
  wire [15:0] proc_6_io_pipe_phv_in_header_6; // @[ipsa.scala 56:25]
  wire [15:0] proc_6_io_pipe_phv_in_header_7; // @[ipsa.scala 56:25]
  wire [15:0] proc_6_io_pipe_phv_in_header_8; // @[ipsa.scala 56:25]
  wire [15:0] proc_6_io_pipe_phv_in_header_9; // @[ipsa.scala 56:25]
  wire [15:0] proc_6_io_pipe_phv_in_header_10; // @[ipsa.scala 56:25]
  wire [15:0] proc_6_io_pipe_phv_in_header_11; // @[ipsa.scala 56:25]
  wire [15:0] proc_6_io_pipe_phv_in_header_12; // @[ipsa.scala 56:25]
  wire [15:0] proc_6_io_pipe_phv_in_header_13; // @[ipsa.scala 56:25]
  wire [15:0] proc_6_io_pipe_phv_in_header_14; // @[ipsa.scala 56:25]
  wire [15:0] proc_6_io_pipe_phv_in_header_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_parse_current_state; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_in_parse_current_offset; // @[ipsa.scala 56:25]
  wire [15:0] proc_6_io_pipe_phv_in_parse_transition_field; // @[ipsa.scala 56:25]
  wire [3:0] proc_6_io_pipe_phv_in_next_processor_id; // @[ipsa.scala 56:25]
  wire  proc_6_io_pipe_phv_in_next_config_id; // @[ipsa.scala 56:25]
  wire  proc_6_io_pipe_phv_in_is_valid_processor; // @[ipsa.scala 56:25]
  wire  proc_6_io_pipe_phv_in_valid; // @[ipsa.scala 56:25]
  wire  proc_6_io_pipe_phv_in_last; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_0; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_1; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_2; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_3; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_4; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_5; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_6; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_7; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_8; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_9; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_10; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_11; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_12; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_13; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_14; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_16; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_17; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_18; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_19; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_20; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_21; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_22; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_23; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_24; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_25; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_26; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_27; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_28; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_29; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_30; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_31; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_32; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_33; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_34; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_35; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_36; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_37; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_38; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_39; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_40; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_41; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_42; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_43; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_44; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_45; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_46; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_47; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_48; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_49; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_50; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_51; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_52; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_53; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_54; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_55; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_56; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_57; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_58; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_59; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_60; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_61; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_62; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_63; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_64; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_65; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_66; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_67; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_68; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_69; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_70; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_71; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_72; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_73; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_74; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_75; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_76; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_77; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_78; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_79; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_80; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_81; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_82; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_83; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_84; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_85; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_86; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_87; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_88; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_89; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_90; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_91; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_92; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_93; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_94; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_95; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_96; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_97; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_98; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_99; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_100; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_101; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_102; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_103; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_104; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_105; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_106; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_107; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_108; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_109; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_110; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_111; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_112; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_113; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_114; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_115; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_116; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_117; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_118; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_119; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_120; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_121; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_122; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_123; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_124; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_125; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_126; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_127; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_128; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_129; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_130; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_131; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_132; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_133; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_134; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_135; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_136; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_137; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_138; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_139; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_140; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_141; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_142; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_143; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_144; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_145; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_146; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_147; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_148; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_149; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_150; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_151; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_152; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_153; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_154; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_155; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_156; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_157; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_158; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_159; // @[ipsa.scala 56:25]
  wire [15:0] proc_6_io_pipe_phv_out_header_0; // @[ipsa.scala 56:25]
  wire [15:0] proc_6_io_pipe_phv_out_header_1; // @[ipsa.scala 56:25]
  wire [15:0] proc_6_io_pipe_phv_out_header_2; // @[ipsa.scala 56:25]
  wire [15:0] proc_6_io_pipe_phv_out_header_3; // @[ipsa.scala 56:25]
  wire [15:0] proc_6_io_pipe_phv_out_header_4; // @[ipsa.scala 56:25]
  wire [15:0] proc_6_io_pipe_phv_out_header_5; // @[ipsa.scala 56:25]
  wire [15:0] proc_6_io_pipe_phv_out_header_6; // @[ipsa.scala 56:25]
  wire [15:0] proc_6_io_pipe_phv_out_header_7; // @[ipsa.scala 56:25]
  wire [15:0] proc_6_io_pipe_phv_out_header_8; // @[ipsa.scala 56:25]
  wire [15:0] proc_6_io_pipe_phv_out_header_9; // @[ipsa.scala 56:25]
  wire [15:0] proc_6_io_pipe_phv_out_header_10; // @[ipsa.scala 56:25]
  wire [15:0] proc_6_io_pipe_phv_out_header_11; // @[ipsa.scala 56:25]
  wire [15:0] proc_6_io_pipe_phv_out_header_12; // @[ipsa.scala 56:25]
  wire [15:0] proc_6_io_pipe_phv_out_header_13; // @[ipsa.scala 56:25]
  wire [15:0] proc_6_io_pipe_phv_out_header_14; // @[ipsa.scala 56:25]
  wire [15:0] proc_6_io_pipe_phv_out_header_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 56:25]
  wire [7:0] proc_6_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 56:25]
  wire [15:0] proc_6_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 56:25]
  wire [3:0] proc_6_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 56:25]
  wire  proc_6_io_pipe_phv_out_next_config_id; // @[ipsa.scala 56:25]
  wire  proc_6_io_pipe_phv_out_valid; // @[ipsa.scala 56:25]
  wire  proc_6_io_pipe_phv_out_last; // @[ipsa.scala 56:25]
  wire  proc_7_clock; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_0; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_1; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_2; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_3; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_4; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_5; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_6; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_7; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_8; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_9; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_10; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_11; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_12; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_13; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_14; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_16; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_17; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_18; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_19; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_20; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_21; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_22; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_23; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_24; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_25; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_26; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_27; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_28; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_29; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_30; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_31; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_32; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_33; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_34; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_35; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_36; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_37; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_38; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_39; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_40; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_41; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_42; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_43; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_44; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_45; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_46; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_47; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_48; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_49; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_50; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_51; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_52; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_53; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_54; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_55; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_56; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_57; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_58; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_59; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_60; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_61; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_62; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_63; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_64; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_65; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_66; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_67; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_68; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_69; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_70; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_71; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_72; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_73; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_74; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_75; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_76; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_77; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_78; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_79; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_80; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_81; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_82; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_83; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_84; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_85; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_86; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_87; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_88; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_89; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_90; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_91; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_92; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_93; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_94; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_95; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_96; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_97; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_98; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_99; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_100; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_101; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_102; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_103; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_104; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_105; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_106; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_107; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_108; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_109; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_110; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_111; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_112; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_113; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_114; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_115; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_116; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_117; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_118; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_119; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_120; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_121; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_122; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_123; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_124; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_125; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_126; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_127; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_128; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_129; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_130; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_131; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_132; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_133; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_134; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_135; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_136; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_137; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_138; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_139; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_140; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_141; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_142; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_143; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_144; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_145; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_146; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_147; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_148; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_149; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_150; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_151; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_152; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_153; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_154; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_155; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_156; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_157; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_158; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_159; // @[ipsa.scala 56:25]
  wire [15:0] proc_7_io_pipe_phv_in_header_0; // @[ipsa.scala 56:25]
  wire [15:0] proc_7_io_pipe_phv_in_header_1; // @[ipsa.scala 56:25]
  wire [15:0] proc_7_io_pipe_phv_in_header_2; // @[ipsa.scala 56:25]
  wire [15:0] proc_7_io_pipe_phv_in_header_3; // @[ipsa.scala 56:25]
  wire [15:0] proc_7_io_pipe_phv_in_header_4; // @[ipsa.scala 56:25]
  wire [15:0] proc_7_io_pipe_phv_in_header_5; // @[ipsa.scala 56:25]
  wire [15:0] proc_7_io_pipe_phv_in_header_6; // @[ipsa.scala 56:25]
  wire [15:0] proc_7_io_pipe_phv_in_header_7; // @[ipsa.scala 56:25]
  wire [15:0] proc_7_io_pipe_phv_in_header_8; // @[ipsa.scala 56:25]
  wire [15:0] proc_7_io_pipe_phv_in_header_9; // @[ipsa.scala 56:25]
  wire [15:0] proc_7_io_pipe_phv_in_header_10; // @[ipsa.scala 56:25]
  wire [15:0] proc_7_io_pipe_phv_in_header_11; // @[ipsa.scala 56:25]
  wire [15:0] proc_7_io_pipe_phv_in_header_12; // @[ipsa.scala 56:25]
  wire [15:0] proc_7_io_pipe_phv_in_header_13; // @[ipsa.scala 56:25]
  wire [15:0] proc_7_io_pipe_phv_in_header_14; // @[ipsa.scala 56:25]
  wire [15:0] proc_7_io_pipe_phv_in_header_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_parse_current_state; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_in_parse_current_offset; // @[ipsa.scala 56:25]
  wire [15:0] proc_7_io_pipe_phv_in_parse_transition_field; // @[ipsa.scala 56:25]
  wire [3:0] proc_7_io_pipe_phv_in_next_processor_id; // @[ipsa.scala 56:25]
  wire  proc_7_io_pipe_phv_in_next_config_id; // @[ipsa.scala 56:25]
  wire  proc_7_io_pipe_phv_in_is_valid_processor; // @[ipsa.scala 56:25]
  wire  proc_7_io_pipe_phv_in_valid; // @[ipsa.scala 56:25]
  wire  proc_7_io_pipe_phv_in_last; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_0; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_1; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_2; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_3; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_4; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_5; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_6; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_7; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_8; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_9; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_10; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_11; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_12; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_13; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_14; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_16; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_17; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_18; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_19; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_20; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_21; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_22; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_23; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_24; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_25; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_26; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_27; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_28; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_29; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_30; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_31; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_32; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_33; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_34; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_35; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_36; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_37; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_38; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_39; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_40; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_41; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_42; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_43; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_44; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_45; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_46; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_47; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_48; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_49; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_50; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_51; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_52; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_53; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_54; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_55; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_56; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_57; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_58; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_59; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_60; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_61; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_62; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_63; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_64; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_65; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_66; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_67; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_68; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_69; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_70; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_71; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_72; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_73; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_74; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_75; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_76; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_77; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_78; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_79; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_80; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_81; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_82; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_83; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_84; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_85; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_86; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_87; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_88; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_89; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_90; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_91; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_92; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_93; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_94; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_95; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_96; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_97; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_98; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_99; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_100; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_101; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_102; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_103; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_104; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_105; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_106; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_107; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_108; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_109; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_110; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_111; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_112; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_113; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_114; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_115; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_116; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_117; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_118; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_119; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_120; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_121; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_122; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_123; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_124; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_125; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_126; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_127; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_128; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_129; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_130; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_131; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_132; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_133; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_134; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_135; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_136; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_137; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_138; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_139; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_140; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_141; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_142; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_143; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_144; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_145; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_146; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_147; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_148; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_149; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_150; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_151; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_152; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_153; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_154; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_155; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_156; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_157; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_158; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_159; // @[ipsa.scala 56:25]
  wire [15:0] proc_7_io_pipe_phv_out_header_0; // @[ipsa.scala 56:25]
  wire [15:0] proc_7_io_pipe_phv_out_header_1; // @[ipsa.scala 56:25]
  wire [15:0] proc_7_io_pipe_phv_out_header_2; // @[ipsa.scala 56:25]
  wire [15:0] proc_7_io_pipe_phv_out_header_3; // @[ipsa.scala 56:25]
  wire [15:0] proc_7_io_pipe_phv_out_header_4; // @[ipsa.scala 56:25]
  wire [15:0] proc_7_io_pipe_phv_out_header_5; // @[ipsa.scala 56:25]
  wire [15:0] proc_7_io_pipe_phv_out_header_6; // @[ipsa.scala 56:25]
  wire [15:0] proc_7_io_pipe_phv_out_header_7; // @[ipsa.scala 56:25]
  wire [15:0] proc_7_io_pipe_phv_out_header_8; // @[ipsa.scala 56:25]
  wire [15:0] proc_7_io_pipe_phv_out_header_9; // @[ipsa.scala 56:25]
  wire [15:0] proc_7_io_pipe_phv_out_header_10; // @[ipsa.scala 56:25]
  wire [15:0] proc_7_io_pipe_phv_out_header_11; // @[ipsa.scala 56:25]
  wire [15:0] proc_7_io_pipe_phv_out_header_12; // @[ipsa.scala 56:25]
  wire [15:0] proc_7_io_pipe_phv_out_header_13; // @[ipsa.scala 56:25]
  wire [15:0] proc_7_io_pipe_phv_out_header_14; // @[ipsa.scala 56:25]
  wire [15:0] proc_7_io_pipe_phv_out_header_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 56:25]
  wire [7:0] proc_7_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 56:25]
  wire [15:0] proc_7_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 56:25]
  wire [3:0] proc_7_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 56:25]
  wire  proc_7_io_pipe_phv_out_next_config_id; // @[ipsa.scala 56:25]
  wire  proc_7_io_pipe_phv_out_valid; // @[ipsa.scala 56:25]
  wire  proc_7_io_pipe_phv_out_last; // @[ipsa.scala 56:25]
  wire  proc_8_clock; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_0; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_1; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_2; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_3; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_4; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_5; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_6; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_7; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_8; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_9; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_10; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_11; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_12; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_13; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_14; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_16; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_17; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_18; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_19; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_20; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_21; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_22; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_23; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_24; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_25; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_26; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_27; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_28; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_29; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_30; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_31; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_32; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_33; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_34; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_35; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_36; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_37; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_38; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_39; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_40; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_41; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_42; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_43; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_44; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_45; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_46; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_47; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_48; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_49; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_50; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_51; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_52; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_53; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_54; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_55; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_56; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_57; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_58; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_59; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_60; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_61; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_62; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_63; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_64; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_65; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_66; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_67; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_68; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_69; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_70; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_71; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_72; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_73; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_74; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_75; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_76; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_77; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_78; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_79; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_80; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_81; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_82; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_83; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_84; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_85; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_86; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_87; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_88; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_89; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_90; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_91; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_92; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_93; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_94; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_95; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_96; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_97; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_98; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_99; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_100; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_101; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_102; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_103; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_104; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_105; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_106; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_107; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_108; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_109; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_110; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_111; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_112; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_113; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_114; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_115; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_116; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_117; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_118; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_119; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_120; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_121; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_122; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_123; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_124; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_125; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_126; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_127; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_128; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_129; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_130; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_131; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_132; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_133; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_134; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_135; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_136; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_137; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_138; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_139; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_140; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_141; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_142; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_143; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_144; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_145; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_146; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_147; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_148; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_149; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_150; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_151; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_152; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_153; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_154; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_155; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_156; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_157; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_158; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_159; // @[ipsa.scala 56:25]
  wire [15:0] proc_8_io_pipe_phv_in_header_0; // @[ipsa.scala 56:25]
  wire [15:0] proc_8_io_pipe_phv_in_header_1; // @[ipsa.scala 56:25]
  wire [15:0] proc_8_io_pipe_phv_in_header_2; // @[ipsa.scala 56:25]
  wire [15:0] proc_8_io_pipe_phv_in_header_3; // @[ipsa.scala 56:25]
  wire [15:0] proc_8_io_pipe_phv_in_header_4; // @[ipsa.scala 56:25]
  wire [15:0] proc_8_io_pipe_phv_in_header_5; // @[ipsa.scala 56:25]
  wire [15:0] proc_8_io_pipe_phv_in_header_6; // @[ipsa.scala 56:25]
  wire [15:0] proc_8_io_pipe_phv_in_header_7; // @[ipsa.scala 56:25]
  wire [15:0] proc_8_io_pipe_phv_in_header_8; // @[ipsa.scala 56:25]
  wire [15:0] proc_8_io_pipe_phv_in_header_9; // @[ipsa.scala 56:25]
  wire [15:0] proc_8_io_pipe_phv_in_header_10; // @[ipsa.scala 56:25]
  wire [15:0] proc_8_io_pipe_phv_in_header_11; // @[ipsa.scala 56:25]
  wire [15:0] proc_8_io_pipe_phv_in_header_12; // @[ipsa.scala 56:25]
  wire [15:0] proc_8_io_pipe_phv_in_header_13; // @[ipsa.scala 56:25]
  wire [15:0] proc_8_io_pipe_phv_in_header_14; // @[ipsa.scala 56:25]
  wire [15:0] proc_8_io_pipe_phv_in_header_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_parse_current_state; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_in_parse_current_offset; // @[ipsa.scala 56:25]
  wire [15:0] proc_8_io_pipe_phv_in_parse_transition_field; // @[ipsa.scala 56:25]
  wire [3:0] proc_8_io_pipe_phv_in_next_processor_id; // @[ipsa.scala 56:25]
  wire  proc_8_io_pipe_phv_in_next_config_id; // @[ipsa.scala 56:25]
  wire  proc_8_io_pipe_phv_in_is_valid_processor; // @[ipsa.scala 56:25]
  wire  proc_8_io_pipe_phv_in_valid; // @[ipsa.scala 56:25]
  wire  proc_8_io_pipe_phv_in_last; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_0; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_1; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_2; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_3; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_4; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_5; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_6; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_7; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_8; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_9; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_10; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_11; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_12; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_13; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_14; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_16; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_17; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_18; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_19; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_20; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_21; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_22; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_23; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_24; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_25; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_26; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_27; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_28; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_29; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_30; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_31; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_32; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_33; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_34; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_35; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_36; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_37; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_38; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_39; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_40; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_41; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_42; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_43; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_44; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_45; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_46; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_47; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_48; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_49; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_50; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_51; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_52; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_53; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_54; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_55; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_56; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_57; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_58; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_59; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_60; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_61; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_62; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_63; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_64; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_65; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_66; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_67; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_68; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_69; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_70; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_71; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_72; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_73; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_74; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_75; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_76; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_77; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_78; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_79; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_80; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_81; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_82; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_83; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_84; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_85; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_86; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_87; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_88; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_89; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_90; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_91; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_92; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_93; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_94; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_95; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_96; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_97; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_98; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_99; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_100; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_101; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_102; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_103; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_104; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_105; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_106; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_107; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_108; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_109; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_110; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_111; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_112; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_113; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_114; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_115; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_116; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_117; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_118; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_119; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_120; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_121; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_122; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_123; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_124; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_125; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_126; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_127; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_128; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_129; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_130; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_131; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_132; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_133; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_134; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_135; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_136; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_137; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_138; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_139; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_140; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_141; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_142; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_143; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_144; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_145; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_146; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_147; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_148; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_149; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_150; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_151; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_152; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_153; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_154; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_155; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_156; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_157; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_158; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_159; // @[ipsa.scala 56:25]
  wire [15:0] proc_8_io_pipe_phv_out_header_0; // @[ipsa.scala 56:25]
  wire [15:0] proc_8_io_pipe_phv_out_header_1; // @[ipsa.scala 56:25]
  wire [15:0] proc_8_io_pipe_phv_out_header_2; // @[ipsa.scala 56:25]
  wire [15:0] proc_8_io_pipe_phv_out_header_3; // @[ipsa.scala 56:25]
  wire [15:0] proc_8_io_pipe_phv_out_header_4; // @[ipsa.scala 56:25]
  wire [15:0] proc_8_io_pipe_phv_out_header_5; // @[ipsa.scala 56:25]
  wire [15:0] proc_8_io_pipe_phv_out_header_6; // @[ipsa.scala 56:25]
  wire [15:0] proc_8_io_pipe_phv_out_header_7; // @[ipsa.scala 56:25]
  wire [15:0] proc_8_io_pipe_phv_out_header_8; // @[ipsa.scala 56:25]
  wire [15:0] proc_8_io_pipe_phv_out_header_9; // @[ipsa.scala 56:25]
  wire [15:0] proc_8_io_pipe_phv_out_header_10; // @[ipsa.scala 56:25]
  wire [15:0] proc_8_io_pipe_phv_out_header_11; // @[ipsa.scala 56:25]
  wire [15:0] proc_8_io_pipe_phv_out_header_12; // @[ipsa.scala 56:25]
  wire [15:0] proc_8_io_pipe_phv_out_header_13; // @[ipsa.scala 56:25]
  wire [15:0] proc_8_io_pipe_phv_out_header_14; // @[ipsa.scala 56:25]
  wire [15:0] proc_8_io_pipe_phv_out_header_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 56:25]
  wire [7:0] proc_8_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 56:25]
  wire [15:0] proc_8_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 56:25]
  wire [3:0] proc_8_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 56:25]
  wire  proc_8_io_pipe_phv_out_next_config_id; // @[ipsa.scala 56:25]
  wire  proc_8_io_pipe_phv_out_valid; // @[ipsa.scala 56:25]
  wire  proc_8_io_pipe_phv_out_last; // @[ipsa.scala 56:25]
  wire  proc_9_clock; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_0; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_1; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_2; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_3; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_4; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_5; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_6; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_7; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_8; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_9; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_10; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_11; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_12; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_13; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_14; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_16; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_17; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_18; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_19; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_20; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_21; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_22; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_23; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_24; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_25; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_26; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_27; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_28; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_29; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_30; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_31; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_32; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_33; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_34; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_35; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_36; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_37; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_38; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_39; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_40; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_41; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_42; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_43; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_44; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_45; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_46; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_47; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_48; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_49; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_50; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_51; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_52; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_53; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_54; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_55; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_56; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_57; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_58; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_59; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_60; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_61; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_62; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_63; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_64; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_65; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_66; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_67; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_68; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_69; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_70; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_71; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_72; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_73; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_74; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_75; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_76; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_77; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_78; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_79; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_80; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_81; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_82; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_83; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_84; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_85; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_86; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_87; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_88; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_89; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_90; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_91; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_92; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_93; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_94; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_95; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_96; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_97; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_98; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_99; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_100; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_101; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_102; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_103; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_104; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_105; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_106; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_107; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_108; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_109; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_110; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_111; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_112; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_113; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_114; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_115; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_116; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_117; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_118; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_119; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_120; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_121; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_122; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_123; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_124; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_125; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_126; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_127; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_128; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_129; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_130; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_131; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_132; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_133; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_134; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_135; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_136; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_137; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_138; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_139; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_140; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_141; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_142; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_143; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_144; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_145; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_146; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_147; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_148; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_149; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_150; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_151; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_152; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_153; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_154; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_155; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_156; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_157; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_158; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_159; // @[ipsa.scala 56:25]
  wire [15:0] proc_9_io_pipe_phv_in_header_0; // @[ipsa.scala 56:25]
  wire [15:0] proc_9_io_pipe_phv_in_header_1; // @[ipsa.scala 56:25]
  wire [15:0] proc_9_io_pipe_phv_in_header_2; // @[ipsa.scala 56:25]
  wire [15:0] proc_9_io_pipe_phv_in_header_3; // @[ipsa.scala 56:25]
  wire [15:0] proc_9_io_pipe_phv_in_header_4; // @[ipsa.scala 56:25]
  wire [15:0] proc_9_io_pipe_phv_in_header_5; // @[ipsa.scala 56:25]
  wire [15:0] proc_9_io_pipe_phv_in_header_6; // @[ipsa.scala 56:25]
  wire [15:0] proc_9_io_pipe_phv_in_header_7; // @[ipsa.scala 56:25]
  wire [15:0] proc_9_io_pipe_phv_in_header_8; // @[ipsa.scala 56:25]
  wire [15:0] proc_9_io_pipe_phv_in_header_9; // @[ipsa.scala 56:25]
  wire [15:0] proc_9_io_pipe_phv_in_header_10; // @[ipsa.scala 56:25]
  wire [15:0] proc_9_io_pipe_phv_in_header_11; // @[ipsa.scala 56:25]
  wire [15:0] proc_9_io_pipe_phv_in_header_12; // @[ipsa.scala 56:25]
  wire [15:0] proc_9_io_pipe_phv_in_header_13; // @[ipsa.scala 56:25]
  wire [15:0] proc_9_io_pipe_phv_in_header_14; // @[ipsa.scala 56:25]
  wire [15:0] proc_9_io_pipe_phv_in_header_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_parse_current_state; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_in_parse_current_offset; // @[ipsa.scala 56:25]
  wire [15:0] proc_9_io_pipe_phv_in_parse_transition_field; // @[ipsa.scala 56:25]
  wire [3:0] proc_9_io_pipe_phv_in_next_processor_id; // @[ipsa.scala 56:25]
  wire  proc_9_io_pipe_phv_in_next_config_id; // @[ipsa.scala 56:25]
  wire  proc_9_io_pipe_phv_in_is_valid_processor; // @[ipsa.scala 56:25]
  wire  proc_9_io_pipe_phv_in_valid; // @[ipsa.scala 56:25]
  wire  proc_9_io_pipe_phv_in_last; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_0; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_1; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_2; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_3; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_4; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_5; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_6; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_7; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_8; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_9; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_10; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_11; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_12; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_13; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_14; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_16; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_17; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_18; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_19; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_20; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_21; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_22; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_23; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_24; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_25; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_26; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_27; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_28; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_29; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_30; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_31; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_32; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_33; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_34; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_35; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_36; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_37; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_38; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_39; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_40; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_41; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_42; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_43; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_44; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_45; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_46; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_47; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_48; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_49; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_50; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_51; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_52; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_53; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_54; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_55; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_56; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_57; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_58; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_59; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_60; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_61; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_62; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_63; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_64; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_65; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_66; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_67; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_68; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_69; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_70; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_71; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_72; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_73; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_74; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_75; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_76; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_77; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_78; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_79; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_80; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_81; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_82; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_83; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_84; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_85; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_86; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_87; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_88; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_89; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_90; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_91; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_92; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_93; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_94; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_95; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_96; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_97; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_98; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_99; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_100; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_101; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_102; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_103; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_104; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_105; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_106; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_107; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_108; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_109; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_110; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_111; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_112; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_113; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_114; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_115; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_116; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_117; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_118; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_119; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_120; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_121; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_122; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_123; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_124; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_125; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_126; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_127; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_128; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_129; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_130; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_131; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_132; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_133; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_134; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_135; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_136; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_137; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_138; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_139; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_140; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_141; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_142; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_143; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_144; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_145; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_146; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_147; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_148; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_149; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_150; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_151; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_152; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_153; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_154; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_155; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_156; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_157; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_158; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_159; // @[ipsa.scala 56:25]
  wire [15:0] proc_9_io_pipe_phv_out_header_0; // @[ipsa.scala 56:25]
  wire [15:0] proc_9_io_pipe_phv_out_header_1; // @[ipsa.scala 56:25]
  wire [15:0] proc_9_io_pipe_phv_out_header_2; // @[ipsa.scala 56:25]
  wire [15:0] proc_9_io_pipe_phv_out_header_3; // @[ipsa.scala 56:25]
  wire [15:0] proc_9_io_pipe_phv_out_header_4; // @[ipsa.scala 56:25]
  wire [15:0] proc_9_io_pipe_phv_out_header_5; // @[ipsa.scala 56:25]
  wire [15:0] proc_9_io_pipe_phv_out_header_6; // @[ipsa.scala 56:25]
  wire [15:0] proc_9_io_pipe_phv_out_header_7; // @[ipsa.scala 56:25]
  wire [15:0] proc_9_io_pipe_phv_out_header_8; // @[ipsa.scala 56:25]
  wire [15:0] proc_9_io_pipe_phv_out_header_9; // @[ipsa.scala 56:25]
  wire [15:0] proc_9_io_pipe_phv_out_header_10; // @[ipsa.scala 56:25]
  wire [15:0] proc_9_io_pipe_phv_out_header_11; // @[ipsa.scala 56:25]
  wire [15:0] proc_9_io_pipe_phv_out_header_12; // @[ipsa.scala 56:25]
  wire [15:0] proc_9_io_pipe_phv_out_header_13; // @[ipsa.scala 56:25]
  wire [15:0] proc_9_io_pipe_phv_out_header_14; // @[ipsa.scala 56:25]
  wire [15:0] proc_9_io_pipe_phv_out_header_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 56:25]
  wire [7:0] proc_9_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 56:25]
  wire [15:0] proc_9_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 56:25]
  wire [3:0] proc_9_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 56:25]
  wire  proc_9_io_pipe_phv_out_next_config_id; // @[ipsa.scala 56:25]
  wire  proc_9_io_pipe_phv_out_valid; // @[ipsa.scala 56:25]
  wire  proc_9_io_pipe_phv_out_last; // @[ipsa.scala 56:25]
  wire  proc_10_clock; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_0; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_1; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_2; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_3; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_4; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_5; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_6; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_7; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_8; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_9; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_10; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_11; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_12; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_13; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_14; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_16; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_17; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_18; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_19; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_20; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_21; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_22; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_23; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_24; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_25; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_26; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_27; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_28; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_29; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_30; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_31; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_32; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_33; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_34; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_35; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_36; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_37; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_38; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_39; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_40; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_41; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_42; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_43; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_44; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_45; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_46; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_47; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_48; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_49; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_50; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_51; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_52; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_53; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_54; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_55; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_56; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_57; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_58; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_59; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_60; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_61; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_62; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_63; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_64; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_65; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_66; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_67; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_68; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_69; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_70; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_71; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_72; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_73; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_74; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_75; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_76; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_77; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_78; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_79; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_80; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_81; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_82; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_83; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_84; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_85; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_86; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_87; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_88; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_89; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_90; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_91; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_92; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_93; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_94; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_95; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_96; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_97; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_98; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_99; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_100; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_101; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_102; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_103; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_104; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_105; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_106; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_107; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_108; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_109; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_110; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_111; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_112; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_113; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_114; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_115; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_116; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_117; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_118; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_119; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_120; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_121; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_122; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_123; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_124; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_125; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_126; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_127; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_128; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_129; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_130; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_131; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_132; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_133; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_134; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_135; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_136; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_137; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_138; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_139; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_140; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_141; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_142; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_143; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_144; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_145; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_146; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_147; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_148; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_149; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_150; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_151; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_152; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_153; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_154; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_155; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_156; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_157; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_158; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_159; // @[ipsa.scala 56:25]
  wire [15:0] proc_10_io_pipe_phv_in_header_0; // @[ipsa.scala 56:25]
  wire [15:0] proc_10_io_pipe_phv_in_header_1; // @[ipsa.scala 56:25]
  wire [15:0] proc_10_io_pipe_phv_in_header_2; // @[ipsa.scala 56:25]
  wire [15:0] proc_10_io_pipe_phv_in_header_3; // @[ipsa.scala 56:25]
  wire [15:0] proc_10_io_pipe_phv_in_header_4; // @[ipsa.scala 56:25]
  wire [15:0] proc_10_io_pipe_phv_in_header_5; // @[ipsa.scala 56:25]
  wire [15:0] proc_10_io_pipe_phv_in_header_6; // @[ipsa.scala 56:25]
  wire [15:0] proc_10_io_pipe_phv_in_header_7; // @[ipsa.scala 56:25]
  wire [15:0] proc_10_io_pipe_phv_in_header_8; // @[ipsa.scala 56:25]
  wire [15:0] proc_10_io_pipe_phv_in_header_9; // @[ipsa.scala 56:25]
  wire [15:0] proc_10_io_pipe_phv_in_header_10; // @[ipsa.scala 56:25]
  wire [15:0] proc_10_io_pipe_phv_in_header_11; // @[ipsa.scala 56:25]
  wire [15:0] proc_10_io_pipe_phv_in_header_12; // @[ipsa.scala 56:25]
  wire [15:0] proc_10_io_pipe_phv_in_header_13; // @[ipsa.scala 56:25]
  wire [15:0] proc_10_io_pipe_phv_in_header_14; // @[ipsa.scala 56:25]
  wire [15:0] proc_10_io_pipe_phv_in_header_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_parse_current_state; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_in_parse_current_offset; // @[ipsa.scala 56:25]
  wire [15:0] proc_10_io_pipe_phv_in_parse_transition_field; // @[ipsa.scala 56:25]
  wire [3:0] proc_10_io_pipe_phv_in_next_processor_id; // @[ipsa.scala 56:25]
  wire  proc_10_io_pipe_phv_in_next_config_id; // @[ipsa.scala 56:25]
  wire  proc_10_io_pipe_phv_in_is_valid_processor; // @[ipsa.scala 56:25]
  wire  proc_10_io_pipe_phv_in_valid; // @[ipsa.scala 56:25]
  wire  proc_10_io_pipe_phv_in_last; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_0; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_1; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_2; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_3; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_4; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_5; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_6; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_7; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_8; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_9; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_10; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_11; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_12; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_13; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_14; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_16; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_17; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_18; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_19; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_20; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_21; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_22; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_23; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_24; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_25; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_26; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_27; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_28; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_29; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_30; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_31; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_32; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_33; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_34; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_35; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_36; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_37; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_38; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_39; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_40; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_41; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_42; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_43; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_44; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_45; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_46; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_47; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_48; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_49; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_50; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_51; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_52; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_53; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_54; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_55; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_56; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_57; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_58; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_59; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_60; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_61; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_62; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_63; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_64; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_65; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_66; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_67; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_68; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_69; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_70; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_71; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_72; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_73; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_74; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_75; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_76; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_77; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_78; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_79; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_80; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_81; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_82; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_83; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_84; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_85; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_86; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_87; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_88; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_89; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_90; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_91; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_92; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_93; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_94; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_95; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_96; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_97; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_98; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_99; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_100; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_101; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_102; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_103; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_104; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_105; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_106; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_107; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_108; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_109; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_110; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_111; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_112; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_113; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_114; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_115; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_116; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_117; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_118; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_119; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_120; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_121; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_122; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_123; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_124; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_125; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_126; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_127; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_128; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_129; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_130; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_131; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_132; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_133; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_134; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_135; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_136; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_137; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_138; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_139; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_140; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_141; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_142; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_143; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_144; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_145; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_146; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_147; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_148; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_149; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_150; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_151; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_152; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_153; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_154; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_155; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_156; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_157; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_158; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_159; // @[ipsa.scala 56:25]
  wire [15:0] proc_10_io_pipe_phv_out_header_0; // @[ipsa.scala 56:25]
  wire [15:0] proc_10_io_pipe_phv_out_header_1; // @[ipsa.scala 56:25]
  wire [15:0] proc_10_io_pipe_phv_out_header_2; // @[ipsa.scala 56:25]
  wire [15:0] proc_10_io_pipe_phv_out_header_3; // @[ipsa.scala 56:25]
  wire [15:0] proc_10_io_pipe_phv_out_header_4; // @[ipsa.scala 56:25]
  wire [15:0] proc_10_io_pipe_phv_out_header_5; // @[ipsa.scala 56:25]
  wire [15:0] proc_10_io_pipe_phv_out_header_6; // @[ipsa.scala 56:25]
  wire [15:0] proc_10_io_pipe_phv_out_header_7; // @[ipsa.scala 56:25]
  wire [15:0] proc_10_io_pipe_phv_out_header_8; // @[ipsa.scala 56:25]
  wire [15:0] proc_10_io_pipe_phv_out_header_9; // @[ipsa.scala 56:25]
  wire [15:0] proc_10_io_pipe_phv_out_header_10; // @[ipsa.scala 56:25]
  wire [15:0] proc_10_io_pipe_phv_out_header_11; // @[ipsa.scala 56:25]
  wire [15:0] proc_10_io_pipe_phv_out_header_12; // @[ipsa.scala 56:25]
  wire [15:0] proc_10_io_pipe_phv_out_header_13; // @[ipsa.scala 56:25]
  wire [15:0] proc_10_io_pipe_phv_out_header_14; // @[ipsa.scala 56:25]
  wire [15:0] proc_10_io_pipe_phv_out_header_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 56:25]
  wire [7:0] proc_10_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 56:25]
  wire [15:0] proc_10_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 56:25]
  wire [3:0] proc_10_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 56:25]
  wire  proc_10_io_pipe_phv_out_next_config_id; // @[ipsa.scala 56:25]
  wire  proc_10_io_pipe_phv_out_valid; // @[ipsa.scala 56:25]
  wire  proc_10_io_pipe_phv_out_last; // @[ipsa.scala 56:25]
  wire  proc_11_clock; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_0; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_1; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_2; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_3; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_4; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_5; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_6; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_7; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_8; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_9; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_10; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_11; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_12; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_13; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_14; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_16; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_17; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_18; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_19; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_20; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_21; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_22; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_23; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_24; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_25; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_26; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_27; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_28; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_29; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_30; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_31; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_32; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_33; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_34; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_35; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_36; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_37; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_38; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_39; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_40; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_41; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_42; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_43; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_44; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_45; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_46; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_47; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_48; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_49; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_50; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_51; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_52; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_53; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_54; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_55; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_56; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_57; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_58; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_59; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_60; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_61; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_62; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_63; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_64; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_65; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_66; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_67; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_68; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_69; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_70; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_71; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_72; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_73; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_74; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_75; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_76; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_77; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_78; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_79; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_80; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_81; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_82; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_83; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_84; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_85; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_86; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_87; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_88; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_89; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_90; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_91; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_92; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_93; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_94; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_95; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_96; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_97; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_98; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_99; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_100; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_101; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_102; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_103; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_104; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_105; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_106; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_107; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_108; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_109; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_110; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_111; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_112; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_113; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_114; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_115; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_116; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_117; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_118; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_119; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_120; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_121; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_122; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_123; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_124; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_125; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_126; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_127; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_128; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_129; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_130; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_131; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_132; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_133; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_134; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_135; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_136; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_137; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_138; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_139; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_140; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_141; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_142; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_143; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_144; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_145; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_146; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_147; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_148; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_149; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_150; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_151; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_152; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_153; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_154; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_155; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_156; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_157; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_158; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_159; // @[ipsa.scala 56:25]
  wire [15:0] proc_11_io_pipe_phv_in_header_0; // @[ipsa.scala 56:25]
  wire [15:0] proc_11_io_pipe_phv_in_header_1; // @[ipsa.scala 56:25]
  wire [15:0] proc_11_io_pipe_phv_in_header_2; // @[ipsa.scala 56:25]
  wire [15:0] proc_11_io_pipe_phv_in_header_3; // @[ipsa.scala 56:25]
  wire [15:0] proc_11_io_pipe_phv_in_header_4; // @[ipsa.scala 56:25]
  wire [15:0] proc_11_io_pipe_phv_in_header_5; // @[ipsa.scala 56:25]
  wire [15:0] proc_11_io_pipe_phv_in_header_6; // @[ipsa.scala 56:25]
  wire [15:0] proc_11_io_pipe_phv_in_header_7; // @[ipsa.scala 56:25]
  wire [15:0] proc_11_io_pipe_phv_in_header_8; // @[ipsa.scala 56:25]
  wire [15:0] proc_11_io_pipe_phv_in_header_9; // @[ipsa.scala 56:25]
  wire [15:0] proc_11_io_pipe_phv_in_header_10; // @[ipsa.scala 56:25]
  wire [15:0] proc_11_io_pipe_phv_in_header_11; // @[ipsa.scala 56:25]
  wire [15:0] proc_11_io_pipe_phv_in_header_12; // @[ipsa.scala 56:25]
  wire [15:0] proc_11_io_pipe_phv_in_header_13; // @[ipsa.scala 56:25]
  wire [15:0] proc_11_io_pipe_phv_in_header_14; // @[ipsa.scala 56:25]
  wire [15:0] proc_11_io_pipe_phv_in_header_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_parse_current_state; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_in_parse_current_offset; // @[ipsa.scala 56:25]
  wire [15:0] proc_11_io_pipe_phv_in_parse_transition_field; // @[ipsa.scala 56:25]
  wire [3:0] proc_11_io_pipe_phv_in_next_processor_id; // @[ipsa.scala 56:25]
  wire  proc_11_io_pipe_phv_in_next_config_id; // @[ipsa.scala 56:25]
  wire  proc_11_io_pipe_phv_in_is_valid_processor; // @[ipsa.scala 56:25]
  wire  proc_11_io_pipe_phv_in_valid; // @[ipsa.scala 56:25]
  wire  proc_11_io_pipe_phv_in_last; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_0; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_1; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_2; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_3; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_4; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_5; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_6; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_7; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_8; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_9; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_10; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_11; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_12; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_13; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_14; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_16; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_17; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_18; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_19; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_20; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_21; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_22; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_23; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_24; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_25; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_26; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_27; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_28; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_29; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_30; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_31; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_32; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_33; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_34; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_35; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_36; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_37; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_38; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_39; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_40; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_41; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_42; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_43; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_44; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_45; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_46; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_47; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_48; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_49; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_50; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_51; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_52; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_53; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_54; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_55; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_56; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_57; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_58; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_59; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_60; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_61; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_62; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_63; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_64; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_65; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_66; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_67; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_68; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_69; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_70; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_71; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_72; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_73; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_74; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_75; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_76; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_77; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_78; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_79; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_80; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_81; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_82; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_83; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_84; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_85; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_86; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_87; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_88; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_89; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_90; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_91; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_92; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_93; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_94; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_95; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_96; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_97; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_98; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_99; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_100; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_101; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_102; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_103; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_104; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_105; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_106; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_107; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_108; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_109; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_110; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_111; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_112; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_113; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_114; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_115; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_116; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_117; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_118; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_119; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_120; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_121; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_122; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_123; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_124; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_125; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_126; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_127; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_128; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_129; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_130; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_131; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_132; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_133; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_134; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_135; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_136; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_137; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_138; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_139; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_140; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_141; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_142; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_143; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_144; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_145; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_146; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_147; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_148; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_149; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_150; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_151; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_152; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_153; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_154; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_155; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_156; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_157; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_158; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_159; // @[ipsa.scala 56:25]
  wire [15:0] proc_11_io_pipe_phv_out_header_0; // @[ipsa.scala 56:25]
  wire [15:0] proc_11_io_pipe_phv_out_header_1; // @[ipsa.scala 56:25]
  wire [15:0] proc_11_io_pipe_phv_out_header_2; // @[ipsa.scala 56:25]
  wire [15:0] proc_11_io_pipe_phv_out_header_3; // @[ipsa.scala 56:25]
  wire [15:0] proc_11_io_pipe_phv_out_header_4; // @[ipsa.scala 56:25]
  wire [15:0] proc_11_io_pipe_phv_out_header_5; // @[ipsa.scala 56:25]
  wire [15:0] proc_11_io_pipe_phv_out_header_6; // @[ipsa.scala 56:25]
  wire [15:0] proc_11_io_pipe_phv_out_header_7; // @[ipsa.scala 56:25]
  wire [15:0] proc_11_io_pipe_phv_out_header_8; // @[ipsa.scala 56:25]
  wire [15:0] proc_11_io_pipe_phv_out_header_9; // @[ipsa.scala 56:25]
  wire [15:0] proc_11_io_pipe_phv_out_header_10; // @[ipsa.scala 56:25]
  wire [15:0] proc_11_io_pipe_phv_out_header_11; // @[ipsa.scala 56:25]
  wire [15:0] proc_11_io_pipe_phv_out_header_12; // @[ipsa.scala 56:25]
  wire [15:0] proc_11_io_pipe_phv_out_header_13; // @[ipsa.scala 56:25]
  wire [15:0] proc_11_io_pipe_phv_out_header_14; // @[ipsa.scala 56:25]
  wire [15:0] proc_11_io_pipe_phv_out_header_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 56:25]
  wire [7:0] proc_11_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 56:25]
  wire [15:0] proc_11_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 56:25]
  wire [3:0] proc_11_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 56:25]
  wire  proc_11_io_pipe_phv_out_next_config_id; // @[ipsa.scala 56:25]
  wire  proc_11_io_pipe_phv_out_valid; // @[ipsa.scala 56:25]
  wire  proc_11_io_pipe_phv_out_last; // @[ipsa.scala 56:25]
  wire  proc_12_clock; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_0; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_1; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_2; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_3; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_4; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_5; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_6; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_7; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_8; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_9; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_10; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_11; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_12; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_13; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_14; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_16; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_17; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_18; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_19; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_20; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_21; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_22; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_23; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_24; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_25; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_26; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_27; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_28; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_29; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_30; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_31; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_32; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_33; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_34; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_35; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_36; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_37; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_38; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_39; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_40; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_41; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_42; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_43; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_44; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_45; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_46; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_47; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_48; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_49; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_50; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_51; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_52; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_53; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_54; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_55; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_56; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_57; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_58; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_59; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_60; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_61; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_62; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_63; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_64; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_65; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_66; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_67; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_68; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_69; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_70; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_71; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_72; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_73; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_74; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_75; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_76; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_77; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_78; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_79; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_80; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_81; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_82; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_83; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_84; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_85; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_86; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_87; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_88; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_89; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_90; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_91; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_92; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_93; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_94; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_95; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_96; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_97; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_98; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_99; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_100; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_101; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_102; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_103; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_104; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_105; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_106; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_107; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_108; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_109; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_110; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_111; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_112; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_113; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_114; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_115; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_116; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_117; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_118; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_119; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_120; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_121; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_122; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_123; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_124; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_125; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_126; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_127; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_128; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_129; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_130; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_131; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_132; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_133; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_134; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_135; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_136; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_137; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_138; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_139; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_140; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_141; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_142; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_143; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_144; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_145; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_146; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_147; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_148; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_149; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_150; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_151; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_152; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_153; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_154; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_155; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_156; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_157; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_158; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_159; // @[ipsa.scala 56:25]
  wire [15:0] proc_12_io_pipe_phv_in_header_0; // @[ipsa.scala 56:25]
  wire [15:0] proc_12_io_pipe_phv_in_header_1; // @[ipsa.scala 56:25]
  wire [15:0] proc_12_io_pipe_phv_in_header_2; // @[ipsa.scala 56:25]
  wire [15:0] proc_12_io_pipe_phv_in_header_3; // @[ipsa.scala 56:25]
  wire [15:0] proc_12_io_pipe_phv_in_header_4; // @[ipsa.scala 56:25]
  wire [15:0] proc_12_io_pipe_phv_in_header_5; // @[ipsa.scala 56:25]
  wire [15:0] proc_12_io_pipe_phv_in_header_6; // @[ipsa.scala 56:25]
  wire [15:0] proc_12_io_pipe_phv_in_header_7; // @[ipsa.scala 56:25]
  wire [15:0] proc_12_io_pipe_phv_in_header_8; // @[ipsa.scala 56:25]
  wire [15:0] proc_12_io_pipe_phv_in_header_9; // @[ipsa.scala 56:25]
  wire [15:0] proc_12_io_pipe_phv_in_header_10; // @[ipsa.scala 56:25]
  wire [15:0] proc_12_io_pipe_phv_in_header_11; // @[ipsa.scala 56:25]
  wire [15:0] proc_12_io_pipe_phv_in_header_12; // @[ipsa.scala 56:25]
  wire [15:0] proc_12_io_pipe_phv_in_header_13; // @[ipsa.scala 56:25]
  wire [15:0] proc_12_io_pipe_phv_in_header_14; // @[ipsa.scala 56:25]
  wire [15:0] proc_12_io_pipe_phv_in_header_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_parse_current_state; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_in_parse_current_offset; // @[ipsa.scala 56:25]
  wire [15:0] proc_12_io_pipe_phv_in_parse_transition_field; // @[ipsa.scala 56:25]
  wire [3:0] proc_12_io_pipe_phv_in_next_processor_id; // @[ipsa.scala 56:25]
  wire  proc_12_io_pipe_phv_in_next_config_id; // @[ipsa.scala 56:25]
  wire  proc_12_io_pipe_phv_in_is_valid_processor; // @[ipsa.scala 56:25]
  wire  proc_12_io_pipe_phv_in_valid; // @[ipsa.scala 56:25]
  wire  proc_12_io_pipe_phv_in_last; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_0; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_1; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_2; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_3; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_4; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_5; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_6; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_7; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_8; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_9; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_10; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_11; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_12; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_13; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_14; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_16; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_17; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_18; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_19; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_20; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_21; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_22; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_23; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_24; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_25; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_26; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_27; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_28; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_29; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_30; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_31; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_32; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_33; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_34; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_35; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_36; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_37; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_38; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_39; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_40; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_41; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_42; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_43; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_44; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_45; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_46; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_47; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_48; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_49; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_50; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_51; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_52; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_53; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_54; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_55; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_56; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_57; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_58; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_59; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_60; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_61; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_62; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_63; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_64; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_65; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_66; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_67; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_68; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_69; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_70; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_71; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_72; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_73; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_74; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_75; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_76; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_77; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_78; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_79; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_80; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_81; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_82; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_83; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_84; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_85; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_86; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_87; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_88; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_89; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_90; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_91; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_92; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_93; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_94; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_95; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_96; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_97; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_98; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_99; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_100; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_101; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_102; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_103; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_104; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_105; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_106; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_107; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_108; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_109; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_110; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_111; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_112; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_113; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_114; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_115; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_116; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_117; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_118; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_119; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_120; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_121; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_122; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_123; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_124; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_125; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_126; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_127; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_128; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_129; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_130; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_131; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_132; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_133; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_134; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_135; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_136; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_137; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_138; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_139; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_140; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_141; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_142; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_143; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_144; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_145; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_146; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_147; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_148; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_149; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_150; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_151; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_152; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_153; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_154; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_155; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_156; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_157; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_158; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_159; // @[ipsa.scala 56:25]
  wire [15:0] proc_12_io_pipe_phv_out_header_0; // @[ipsa.scala 56:25]
  wire [15:0] proc_12_io_pipe_phv_out_header_1; // @[ipsa.scala 56:25]
  wire [15:0] proc_12_io_pipe_phv_out_header_2; // @[ipsa.scala 56:25]
  wire [15:0] proc_12_io_pipe_phv_out_header_3; // @[ipsa.scala 56:25]
  wire [15:0] proc_12_io_pipe_phv_out_header_4; // @[ipsa.scala 56:25]
  wire [15:0] proc_12_io_pipe_phv_out_header_5; // @[ipsa.scala 56:25]
  wire [15:0] proc_12_io_pipe_phv_out_header_6; // @[ipsa.scala 56:25]
  wire [15:0] proc_12_io_pipe_phv_out_header_7; // @[ipsa.scala 56:25]
  wire [15:0] proc_12_io_pipe_phv_out_header_8; // @[ipsa.scala 56:25]
  wire [15:0] proc_12_io_pipe_phv_out_header_9; // @[ipsa.scala 56:25]
  wire [15:0] proc_12_io_pipe_phv_out_header_10; // @[ipsa.scala 56:25]
  wire [15:0] proc_12_io_pipe_phv_out_header_11; // @[ipsa.scala 56:25]
  wire [15:0] proc_12_io_pipe_phv_out_header_12; // @[ipsa.scala 56:25]
  wire [15:0] proc_12_io_pipe_phv_out_header_13; // @[ipsa.scala 56:25]
  wire [15:0] proc_12_io_pipe_phv_out_header_14; // @[ipsa.scala 56:25]
  wire [15:0] proc_12_io_pipe_phv_out_header_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 56:25]
  wire [7:0] proc_12_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 56:25]
  wire [15:0] proc_12_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 56:25]
  wire [3:0] proc_12_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 56:25]
  wire  proc_12_io_pipe_phv_out_next_config_id; // @[ipsa.scala 56:25]
  wire  proc_12_io_pipe_phv_out_valid; // @[ipsa.scala 56:25]
  wire  proc_12_io_pipe_phv_out_last; // @[ipsa.scala 56:25]
  wire  proc_13_clock; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_0; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_1; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_2; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_3; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_4; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_5; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_6; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_7; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_8; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_9; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_10; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_11; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_12; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_13; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_14; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_16; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_17; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_18; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_19; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_20; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_21; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_22; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_23; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_24; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_25; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_26; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_27; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_28; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_29; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_30; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_31; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_32; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_33; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_34; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_35; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_36; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_37; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_38; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_39; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_40; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_41; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_42; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_43; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_44; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_45; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_46; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_47; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_48; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_49; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_50; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_51; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_52; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_53; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_54; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_55; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_56; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_57; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_58; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_59; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_60; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_61; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_62; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_63; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_64; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_65; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_66; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_67; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_68; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_69; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_70; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_71; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_72; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_73; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_74; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_75; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_76; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_77; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_78; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_79; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_80; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_81; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_82; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_83; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_84; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_85; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_86; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_87; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_88; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_89; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_90; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_91; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_92; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_93; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_94; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_95; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_96; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_97; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_98; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_99; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_100; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_101; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_102; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_103; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_104; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_105; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_106; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_107; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_108; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_109; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_110; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_111; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_112; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_113; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_114; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_115; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_116; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_117; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_118; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_119; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_120; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_121; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_122; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_123; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_124; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_125; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_126; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_127; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_128; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_129; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_130; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_131; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_132; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_133; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_134; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_135; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_136; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_137; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_138; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_139; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_140; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_141; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_142; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_143; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_144; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_145; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_146; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_147; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_148; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_149; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_150; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_151; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_152; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_153; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_154; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_155; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_156; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_157; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_158; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_159; // @[ipsa.scala 56:25]
  wire [15:0] proc_13_io_pipe_phv_in_header_0; // @[ipsa.scala 56:25]
  wire [15:0] proc_13_io_pipe_phv_in_header_1; // @[ipsa.scala 56:25]
  wire [15:0] proc_13_io_pipe_phv_in_header_2; // @[ipsa.scala 56:25]
  wire [15:0] proc_13_io_pipe_phv_in_header_3; // @[ipsa.scala 56:25]
  wire [15:0] proc_13_io_pipe_phv_in_header_4; // @[ipsa.scala 56:25]
  wire [15:0] proc_13_io_pipe_phv_in_header_5; // @[ipsa.scala 56:25]
  wire [15:0] proc_13_io_pipe_phv_in_header_6; // @[ipsa.scala 56:25]
  wire [15:0] proc_13_io_pipe_phv_in_header_7; // @[ipsa.scala 56:25]
  wire [15:0] proc_13_io_pipe_phv_in_header_8; // @[ipsa.scala 56:25]
  wire [15:0] proc_13_io_pipe_phv_in_header_9; // @[ipsa.scala 56:25]
  wire [15:0] proc_13_io_pipe_phv_in_header_10; // @[ipsa.scala 56:25]
  wire [15:0] proc_13_io_pipe_phv_in_header_11; // @[ipsa.scala 56:25]
  wire [15:0] proc_13_io_pipe_phv_in_header_12; // @[ipsa.scala 56:25]
  wire [15:0] proc_13_io_pipe_phv_in_header_13; // @[ipsa.scala 56:25]
  wire [15:0] proc_13_io_pipe_phv_in_header_14; // @[ipsa.scala 56:25]
  wire [15:0] proc_13_io_pipe_phv_in_header_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_parse_current_state; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_in_parse_current_offset; // @[ipsa.scala 56:25]
  wire [15:0] proc_13_io_pipe_phv_in_parse_transition_field; // @[ipsa.scala 56:25]
  wire [3:0] proc_13_io_pipe_phv_in_next_processor_id; // @[ipsa.scala 56:25]
  wire  proc_13_io_pipe_phv_in_next_config_id; // @[ipsa.scala 56:25]
  wire  proc_13_io_pipe_phv_in_is_valid_processor; // @[ipsa.scala 56:25]
  wire  proc_13_io_pipe_phv_in_valid; // @[ipsa.scala 56:25]
  wire  proc_13_io_pipe_phv_in_last; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_0; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_1; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_2; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_3; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_4; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_5; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_6; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_7; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_8; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_9; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_10; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_11; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_12; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_13; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_14; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_16; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_17; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_18; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_19; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_20; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_21; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_22; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_23; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_24; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_25; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_26; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_27; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_28; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_29; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_30; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_31; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_32; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_33; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_34; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_35; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_36; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_37; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_38; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_39; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_40; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_41; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_42; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_43; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_44; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_45; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_46; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_47; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_48; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_49; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_50; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_51; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_52; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_53; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_54; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_55; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_56; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_57; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_58; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_59; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_60; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_61; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_62; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_63; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_64; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_65; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_66; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_67; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_68; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_69; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_70; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_71; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_72; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_73; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_74; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_75; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_76; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_77; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_78; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_79; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_80; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_81; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_82; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_83; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_84; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_85; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_86; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_87; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_88; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_89; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_90; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_91; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_92; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_93; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_94; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_95; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_96; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_97; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_98; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_99; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_100; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_101; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_102; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_103; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_104; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_105; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_106; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_107; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_108; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_109; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_110; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_111; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_112; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_113; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_114; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_115; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_116; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_117; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_118; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_119; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_120; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_121; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_122; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_123; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_124; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_125; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_126; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_127; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_128; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_129; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_130; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_131; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_132; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_133; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_134; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_135; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_136; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_137; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_138; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_139; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_140; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_141; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_142; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_143; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_144; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_145; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_146; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_147; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_148; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_149; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_150; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_151; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_152; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_153; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_154; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_155; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_156; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_157; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_158; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_159; // @[ipsa.scala 56:25]
  wire [15:0] proc_13_io_pipe_phv_out_header_0; // @[ipsa.scala 56:25]
  wire [15:0] proc_13_io_pipe_phv_out_header_1; // @[ipsa.scala 56:25]
  wire [15:0] proc_13_io_pipe_phv_out_header_2; // @[ipsa.scala 56:25]
  wire [15:0] proc_13_io_pipe_phv_out_header_3; // @[ipsa.scala 56:25]
  wire [15:0] proc_13_io_pipe_phv_out_header_4; // @[ipsa.scala 56:25]
  wire [15:0] proc_13_io_pipe_phv_out_header_5; // @[ipsa.scala 56:25]
  wire [15:0] proc_13_io_pipe_phv_out_header_6; // @[ipsa.scala 56:25]
  wire [15:0] proc_13_io_pipe_phv_out_header_7; // @[ipsa.scala 56:25]
  wire [15:0] proc_13_io_pipe_phv_out_header_8; // @[ipsa.scala 56:25]
  wire [15:0] proc_13_io_pipe_phv_out_header_9; // @[ipsa.scala 56:25]
  wire [15:0] proc_13_io_pipe_phv_out_header_10; // @[ipsa.scala 56:25]
  wire [15:0] proc_13_io_pipe_phv_out_header_11; // @[ipsa.scala 56:25]
  wire [15:0] proc_13_io_pipe_phv_out_header_12; // @[ipsa.scala 56:25]
  wire [15:0] proc_13_io_pipe_phv_out_header_13; // @[ipsa.scala 56:25]
  wire [15:0] proc_13_io_pipe_phv_out_header_14; // @[ipsa.scala 56:25]
  wire [15:0] proc_13_io_pipe_phv_out_header_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 56:25]
  wire [7:0] proc_13_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 56:25]
  wire [15:0] proc_13_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 56:25]
  wire [3:0] proc_13_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 56:25]
  wire  proc_13_io_pipe_phv_out_next_config_id; // @[ipsa.scala 56:25]
  wire  proc_13_io_pipe_phv_out_valid; // @[ipsa.scala 56:25]
  wire  proc_13_io_pipe_phv_out_last; // @[ipsa.scala 56:25]
  wire  proc_14_clock; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_0; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_1; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_2; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_3; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_4; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_5; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_6; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_7; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_8; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_9; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_10; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_11; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_12; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_13; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_14; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_16; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_17; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_18; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_19; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_20; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_21; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_22; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_23; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_24; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_25; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_26; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_27; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_28; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_29; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_30; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_31; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_32; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_33; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_34; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_35; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_36; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_37; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_38; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_39; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_40; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_41; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_42; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_43; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_44; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_45; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_46; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_47; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_48; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_49; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_50; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_51; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_52; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_53; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_54; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_55; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_56; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_57; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_58; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_59; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_60; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_61; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_62; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_63; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_64; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_65; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_66; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_67; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_68; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_69; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_70; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_71; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_72; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_73; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_74; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_75; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_76; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_77; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_78; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_79; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_80; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_81; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_82; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_83; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_84; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_85; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_86; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_87; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_88; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_89; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_90; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_91; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_92; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_93; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_94; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_95; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_96; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_97; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_98; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_99; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_100; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_101; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_102; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_103; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_104; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_105; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_106; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_107; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_108; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_109; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_110; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_111; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_112; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_113; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_114; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_115; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_116; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_117; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_118; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_119; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_120; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_121; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_122; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_123; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_124; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_125; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_126; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_127; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_128; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_129; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_130; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_131; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_132; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_133; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_134; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_135; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_136; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_137; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_138; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_139; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_140; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_141; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_142; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_143; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_144; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_145; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_146; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_147; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_148; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_149; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_150; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_151; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_152; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_153; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_154; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_155; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_156; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_157; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_158; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_159; // @[ipsa.scala 56:25]
  wire [15:0] proc_14_io_pipe_phv_in_header_0; // @[ipsa.scala 56:25]
  wire [15:0] proc_14_io_pipe_phv_in_header_1; // @[ipsa.scala 56:25]
  wire [15:0] proc_14_io_pipe_phv_in_header_2; // @[ipsa.scala 56:25]
  wire [15:0] proc_14_io_pipe_phv_in_header_3; // @[ipsa.scala 56:25]
  wire [15:0] proc_14_io_pipe_phv_in_header_4; // @[ipsa.scala 56:25]
  wire [15:0] proc_14_io_pipe_phv_in_header_5; // @[ipsa.scala 56:25]
  wire [15:0] proc_14_io_pipe_phv_in_header_6; // @[ipsa.scala 56:25]
  wire [15:0] proc_14_io_pipe_phv_in_header_7; // @[ipsa.scala 56:25]
  wire [15:0] proc_14_io_pipe_phv_in_header_8; // @[ipsa.scala 56:25]
  wire [15:0] proc_14_io_pipe_phv_in_header_9; // @[ipsa.scala 56:25]
  wire [15:0] proc_14_io_pipe_phv_in_header_10; // @[ipsa.scala 56:25]
  wire [15:0] proc_14_io_pipe_phv_in_header_11; // @[ipsa.scala 56:25]
  wire [15:0] proc_14_io_pipe_phv_in_header_12; // @[ipsa.scala 56:25]
  wire [15:0] proc_14_io_pipe_phv_in_header_13; // @[ipsa.scala 56:25]
  wire [15:0] proc_14_io_pipe_phv_in_header_14; // @[ipsa.scala 56:25]
  wire [15:0] proc_14_io_pipe_phv_in_header_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_parse_current_state; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_in_parse_current_offset; // @[ipsa.scala 56:25]
  wire [15:0] proc_14_io_pipe_phv_in_parse_transition_field; // @[ipsa.scala 56:25]
  wire [3:0] proc_14_io_pipe_phv_in_next_processor_id; // @[ipsa.scala 56:25]
  wire  proc_14_io_pipe_phv_in_next_config_id; // @[ipsa.scala 56:25]
  wire  proc_14_io_pipe_phv_in_is_valid_processor; // @[ipsa.scala 56:25]
  wire  proc_14_io_pipe_phv_in_valid; // @[ipsa.scala 56:25]
  wire  proc_14_io_pipe_phv_in_last; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_0; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_1; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_2; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_3; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_4; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_5; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_6; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_7; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_8; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_9; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_10; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_11; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_12; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_13; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_14; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_16; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_17; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_18; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_19; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_20; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_21; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_22; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_23; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_24; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_25; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_26; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_27; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_28; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_29; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_30; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_31; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_32; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_33; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_34; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_35; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_36; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_37; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_38; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_39; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_40; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_41; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_42; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_43; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_44; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_45; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_46; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_47; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_48; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_49; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_50; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_51; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_52; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_53; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_54; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_55; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_56; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_57; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_58; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_59; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_60; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_61; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_62; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_63; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_64; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_65; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_66; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_67; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_68; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_69; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_70; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_71; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_72; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_73; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_74; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_75; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_76; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_77; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_78; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_79; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_80; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_81; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_82; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_83; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_84; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_85; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_86; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_87; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_88; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_89; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_90; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_91; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_92; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_93; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_94; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_95; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_96; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_97; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_98; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_99; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_100; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_101; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_102; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_103; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_104; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_105; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_106; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_107; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_108; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_109; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_110; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_111; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_112; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_113; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_114; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_115; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_116; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_117; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_118; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_119; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_120; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_121; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_122; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_123; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_124; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_125; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_126; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_127; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_128; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_129; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_130; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_131; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_132; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_133; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_134; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_135; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_136; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_137; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_138; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_139; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_140; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_141; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_142; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_143; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_144; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_145; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_146; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_147; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_148; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_149; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_150; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_151; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_152; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_153; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_154; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_155; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_156; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_157; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_158; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_159; // @[ipsa.scala 56:25]
  wire [15:0] proc_14_io_pipe_phv_out_header_0; // @[ipsa.scala 56:25]
  wire [15:0] proc_14_io_pipe_phv_out_header_1; // @[ipsa.scala 56:25]
  wire [15:0] proc_14_io_pipe_phv_out_header_2; // @[ipsa.scala 56:25]
  wire [15:0] proc_14_io_pipe_phv_out_header_3; // @[ipsa.scala 56:25]
  wire [15:0] proc_14_io_pipe_phv_out_header_4; // @[ipsa.scala 56:25]
  wire [15:0] proc_14_io_pipe_phv_out_header_5; // @[ipsa.scala 56:25]
  wire [15:0] proc_14_io_pipe_phv_out_header_6; // @[ipsa.scala 56:25]
  wire [15:0] proc_14_io_pipe_phv_out_header_7; // @[ipsa.scala 56:25]
  wire [15:0] proc_14_io_pipe_phv_out_header_8; // @[ipsa.scala 56:25]
  wire [15:0] proc_14_io_pipe_phv_out_header_9; // @[ipsa.scala 56:25]
  wire [15:0] proc_14_io_pipe_phv_out_header_10; // @[ipsa.scala 56:25]
  wire [15:0] proc_14_io_pipe_phv_out_header_11; // @[ipsa.scala 56:25]
  wire [15:0] proc_14_io_pipe_phv_out_header_12; // @[ipsa.scala 56:25]
  wire [15:0] proc_14_io_pipe_phv_out_header_13; // @[ipsa.scala 56:25]
  wire [15:0] proc_14_io_pipe_phv_out_header_14; // @[ipsa.scala 56:25]
  wire [15:0] proc_14_io_pipe_phv_out_header_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 56:25]
  wire [7:0] proc_14_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 56:25]
  wire [15:0] proc_14_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 56:25]
  wire [3:0] proc_14_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 56:25]
  wire  proc_14_io_pipe_phv_out_next_config_id; // @[ipsa.scala 56:25]
  wire  proc_14_io_pipe_phv_out_valid; // @[ipsa.scala 56:25]
  wire  proc_14_io_pipe_phv_out_last; // @[ipsa.scala 56:25]
  wire  proc_15_clock; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_0; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_1; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_2; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_3; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_4; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_5; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_6; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_7; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_8; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_9; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_10; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_11; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_12; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_13; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_14; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_16; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_17; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_18; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_19; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_20; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_21; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_22; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_23; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_24; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_25; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_26; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_27; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_28; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_29; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_30; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_31; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_32; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_33; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_34; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_35; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_36; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_37; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_38; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_39; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_40; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_41; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_42; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_43; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_44; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_45; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_46; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_47; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_48; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_49; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_50; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_51; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_52; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_53; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_54; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_55; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_56; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_57; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_58; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_59; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_60; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_61; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_62; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_63; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_64; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_65; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_66; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_67; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_68; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_69; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_70; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_71; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_72; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_73; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_74; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_75; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_76; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_77; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_78; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_79; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_80; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_81; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_82; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_83; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_84; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_85; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_86; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_87; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_88; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_89; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_90; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_91; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_92; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_93; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_94; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_95; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_96; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_97; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_98; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_99; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_100; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_101; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_102; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_103; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_104; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_105; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_106; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_107; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_108; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_109; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_110; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_111; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_112; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_113; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_114; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_115; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_116; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_117; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_118; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_119; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_120; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_121; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_122; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_123; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_124; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_125; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_126; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_127; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_128; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_129; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_130; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_131; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_132; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_133; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_134; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_135; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_136; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_137; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_138; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_139; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_140; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_141; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_142; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_143; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_144; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_145; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_146; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_147; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_148; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_149; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_150; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_151; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_152; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_153; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_154; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_155; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_156; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_157; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_158; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_159; // @[ipsa.scala 56:25]
  wire [15:0] proc_15_io_pipe_phv_in_header_0; // @[ipsa.scala 56:25]
  wire [15:0] proc_15_io_pipe_phv_in_header_1; // @[ipsa.scala 56:25]
  wire [15:0] proc_15_io_pipe_phv_in_header_2; // @[ipsa.scala 56:25]
  wire [15:0] proc_15_io_pipe_phv_in_header_3; // @[ipsa.scala 56:25]
  wire [15:0] proc_15_io_pipe_phv_in_header_4; // @[ipsa.scala 56:25]
  wire [15:0] proc_15_io_pipe_phv_in_header_5; // @[ipsa.scala 56:25]
  wire [15:0] proc_15_io_pipe_phv_in_header_6; // @[ipsa.scala 56:25]
  wire [15:0] proc_15_io_pipe_phv_in_header_7; // @[ipsa.scala 56:25]
  wire [15:0] proc_15_io_pipe_phv_in_header_8; // @[ipsa.scala 56:25]
  wire [15:0] proc_15_io_pipe_phv_in_header_9; // @[ipsa.scala 56:25]
  wire [15:0] proc_15_io_pipe_phv_in_header_10; // @[ipsa.scala 56:25]
  wire [15:0] proc_15_io_pipe_phv_in_header_11; // @[ipsa.scala 56:25]
  wire [15:0] proc_15_io_pipe_phv_in_header_12; // @[ipsa.scala 56:25]
  wire [15:0] proc_15_io_pipe_phv_in_header_13; // @[ipsa.scala 56:25]
  wire [15:0] proc_15_io_pipe_phv_in_header_14; // @[ipsa.scala 56:25]
  wire [15:0] proc_15_io_pipe_phv_in_header_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_parse_current_state; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_in_parse_current_offset; // @[ipsa.scala 56:25]
  wire [15:0] proc_15_io_pipe_phv_in_parse_transition_field; // @[ipsa.scala 56:25]
  wire [3:0] proc_15_io_pipe_phv_in_next_processor_id; // @[ipsa.scala 56:25]
  wire  proc_15_io_pipe_phv_in_next_config_id; // @[ipsa.scala 56:25]
  wire  proc_15_io_pipe_phv_in_is_valid_processor; // @[ipsa.scala 56:25]
  wire  proc_15_io_pipe_phv_in_valid; // @[ipsa.scala 56:25]
  wire  proc_15_io_pipe_phv_in_last; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_0; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_1; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_2; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_3; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_4; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_5; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_6; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_7; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_8; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_9; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_10; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_11; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_12; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_13; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_14; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_16; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_17; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_18; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_19; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_20; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_21; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_22; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_23; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_24; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_25; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_26; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_27; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_28; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_29; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_30; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_31; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_32; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_33; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_34; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_35; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_36; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_37; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_38; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_39; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_40; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_41; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_42; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_43; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_44; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_45; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_46; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_47; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_48; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_49; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_50; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_51; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_52; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_53; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_54; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_55; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_56; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_57; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_58; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_59; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_60; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_61; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_62; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_63; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_64; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_65; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_66; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_67; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_68; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_69; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_70; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_71; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_72; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_73; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_74; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_75; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_76; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_77; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_78; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_79; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_80; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_81; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_82; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_83; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_84; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_85; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_86; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_87; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_88; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_89; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_90; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_91; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_92; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_93; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_94; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_95; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_96; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_97; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_98; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_99; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_100; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_101; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_102; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_103; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_104; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_105; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_106; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_107; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_108; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_109; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_110; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_111; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_112; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_113; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_114; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_115; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_116; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_117; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_118; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_119; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_120; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_121; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_122; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_123; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_124; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_125; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_126; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_127; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_128; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_129; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_130; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_131; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_132; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_133; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_134; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_135; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_136; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_137; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_138; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_139; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_140; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_141; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_142; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_143; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_144; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_145; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_146; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_147; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_148; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_149; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_150; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_151; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_152; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_153; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_154; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_155; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_156; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_157; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_158; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_159; // @[ipsa.scala 56:25]
  wire [15:0] proc_15_io_pipe_phv_out_header_0; // @[ipsa.scala 56:25]
  wire [15:0] proc_15_io_pipe_phv_out_header_1; // @[ipsa.scala 56:25]
  wire [15:0] proc_15_io_pipe_phv_out_header_2; // @[ipsa.scala 56:25]
  wire [15:0] proc_15_io_pipe_phv_out_header_3; // @[ipsa.scala 56:25]
  wire [15:0] proc_15_io_pipe_phv_out_header_4; // @[ipsa.scala 56:25]
  wire [15:0] proc_15_io_pipe_phv_out_header_5; // @[ipsa.scala 56:25]
  wire [15:0] proc_15_io_pipe_phv_out_header_6; // @[ipsa.scala 56:25]
  wire [15:0] proc_15_io_pipe_phv_out_header_7; // @[ipsa.scala 56:25]
  wire [15:0] proc_15_io_pipe_phv_out_header_8; // @[ipsa.scala 56:25]
  wire [15:0] proc_15_io_pipe_phv_out_header_9; // @[ipsa.scala 56:25]
  wire [15:0] proc_15_io_pipe_phv_out_header_10; // @[ipsa.scala 56:25]
  wire [15:0] proc_15_io_pipe_phv_out_header_11; // @[ipsa.scala 56:25]
  wire [15:0] proc_15_io_pipe_phv_out_header_12; // @[ipsa.scala 56:25]
  wire [15:0] proc_15_io_pipe_phv_out_header_13; // @[ipsa.scala 56:25]
  wire [15:0] proc_15_io_pipe_phv_out_header_14; // @[ipsa.scala 56:25]
  wire [15:0] proc_15_io_pipe_phv_out_header_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 56:25]
  wire [7:0] proc_15_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 56:25]
  wire [15:0] proc_15_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 56:25]
  wire [3:0] proc_15_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 56:25]
  wire  proc_15_io_pipe_phv_out_next_config_id; // @[ipsa.scala 56:25]
  wire  proc_15_io_pipe_phv_out_valid; // @[ipsa.scala 56:25]
  wire  proc_15_io_pipe_phv_out_last; // @[ipsa.scala 56:25]
  wire  sram_cluster_0_clock; // @[ipsa.scala 62:25]
  wire  sram_cluster_1_clock; // @[ipsa.scala 62:25]
  wire  sram_cluster_2_clock; // @[ipsa.scala 62:25]
  wire  sram_cluster_3_clock; // @[ipsa.scala 62:25]
  wire  sram_cluster_4_clock; // @[ipsa.scala 62:25]
  wire  sram_cluster_5_clock; // @[ipsa.scala 62:25]
  wire  sram_cluster_6_clock; // @[ipsa.scala 62:25]
  wire  sram_cluster_7_clock; // @[ipsa.scala 62:25]
  wire  init_clock; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_0; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_1; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_2; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_3; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_4; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_5; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_6; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_7; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_8; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_9; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_10; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_11; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_12; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_13; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_14; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_15; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_16; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_17; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_18; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_19; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_20; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_21; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_22; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_23; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_24; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_25; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_26; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_27; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_28; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_29; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_30; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_31; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_32; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_33; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_34; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_35; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_36; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_37; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_38; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_39; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_40; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_41; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_42; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_43; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_44; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_45; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_46; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_47; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_48; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_49; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_50; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_51; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_52; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_53; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_54; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_55; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_56; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_57; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_58; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_59; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_60; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_61; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_62; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_63; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_64; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_65; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_66; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_67; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_68; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_69; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_70; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_71; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_72; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_73; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_74; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_75; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_76; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_77; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_78; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_79; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_80; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_81; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_82; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_83; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_84; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_85; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_86; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_87; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_88; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_89; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_90; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_91; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_92; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_93; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_94; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_95; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_96; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_97; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_98; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_99; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_100; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_101; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_102; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_103; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_104; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_105; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_106; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_107; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_108; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_109; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_110; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_111; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_112; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_113; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_114; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_115; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_116; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_117; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_118; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_119; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_120; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_121; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_122; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_123; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_124; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_125; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_126; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_127; // @[ipsa.scala 74:22]
  wire  init_io_pipe_phv_in_valid; // @[ipsa.scala 74:22]
  wire  init_io_pipe_phv_in_last; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_0; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_1; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_2; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_3; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_4; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_5; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_6; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_7; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_8; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_9; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_10; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_11; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_12; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_13; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_14; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_15; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_16; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_17; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_18; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_19; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_20; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_21; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_22; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_23; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_24; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_25; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_26; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_27; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_28; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_29; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_30; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_31; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_32; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_33; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_34; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_35; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_36; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_37; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_38; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_39; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_40; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_41; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_42; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_43; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_44; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_45; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_46; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_47; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_48; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_49; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_50; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_51; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_52; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_53; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_54; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_55; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_56; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_57; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_58; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_59; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_60; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_61; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_62; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_63; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_64; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_65; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_66; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_67; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_68; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_69; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_70; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_71; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_72; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_73; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_74; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_75; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_76; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_77; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_78; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_79; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_80; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_81; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_82; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_83; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_84; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_85; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_86; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_87; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_88; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_89; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_90; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_91; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_92; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_93; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_94; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_95; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_96; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_97; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_98; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_99; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_100; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_101; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_102; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_103; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_104; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_105; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_106; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_107; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_108; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_109; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_110; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_111; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_112; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_113; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_114; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_115; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_116; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_117; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_118; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_119; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_120; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_121; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_122; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_123; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_124; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_125; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_126; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_127; // @[ipsa.scala 74:22]
  wire  init_io_pipe_phv_out_valid; // @[ipsa.scala 74:22]
  wire  init_io_pipe_phv_out_last; // @[ipsa.scala 74:22]
  wire  trans_0_clock; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_0; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_1; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_2; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_3; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_4; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_5; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_6; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_7; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_8; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_9; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_10; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_11; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_12; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_13; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_14; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_16; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_17; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_18; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_19; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_20; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_21; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_22; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_23; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_24; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_25; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_26; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_27; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_28; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_29; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_30; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_31; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_32; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_33; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_34; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_35; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_36; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_37; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_38; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_39; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_40; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_41; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_42; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_43; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_44; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_45; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_46; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_47; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_48; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_49; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_50; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_51; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_52; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_53; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_54; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_55; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_56; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_57; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_58; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_59; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_60; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_61; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_62; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_63; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_64; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_65; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_66; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_67; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_68; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_69; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_70; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_71; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_72; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_73; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_74; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_75; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_76; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_77; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_78; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_79; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_80; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_81; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_82; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_83; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_84; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_85; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_86; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_87; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_88; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_89; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_90; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_91; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_92; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_93; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_94; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_95; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_96; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_97; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_98; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_99; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_100; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_101; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_102; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_103; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_104; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_105; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_106; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_107; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_108; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_109; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_110; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_111; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_112; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_113; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_114; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_115; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_116; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_117; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_118; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_119; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_120; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_121; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_122; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_123; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_124; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_125; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_126; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_127; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_128; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_129; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_130; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_131; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_132; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_133; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_134; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_135; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_136; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_137; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_138; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_139; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_140; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_141; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_142; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_143; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_144; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_145; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_146; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_147; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_148; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_149; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_150; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_151; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_152; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_153; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_154; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_155; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_156; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_157; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_158; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_159; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_in_header_0; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_in_header_1; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_in_header_2; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_in_header_3; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_in_header_4; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_in_header_5; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_in_header_6; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_in_header_7; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_in_header_8; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_in_header_9; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_in_header_10; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_in_header_11; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_in_header_12; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_in_header_13; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_in_header_14; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_in_header_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_parse_current_state; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_parse_current_offset; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_in_parse_transition_field; // @[ipsa.scala 79:25]
  wire [3:0] trans_0_io_pipe_phv_in_next_processor_id; // @[ipsa.scala 79:25]
  wire  trans_0_io_pipe_phv_in_next_config_id; // @[ipsa.scala 79:25]
  wire  trans_0_io_pipe_phv_in_valid; // @[ipsa.scala 79:25]
  wire  trans_0_io_pipe_phv_in_last; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_0; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_1; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_2; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_3; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_4; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_5; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_6; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_7; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_8; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_9; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_10; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_11; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_12; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_13; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_14; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_16; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_17; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_18; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_19; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_20; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_21; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_22; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_23; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_24; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_25; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_26; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_27; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_28; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_29; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_30; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_31; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_32; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_33; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_34; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_35; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_36; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_37; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_38; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_39; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_40; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_41; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_42; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_43; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_44; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_45; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_46; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_47; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_48; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_49; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_50; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_51; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_52; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_53; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_54; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_55; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_56; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_57; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_58; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_59; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_60; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_61; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_62; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_63; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_64; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_65; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_66; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_67; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_68; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_69; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_70; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_71; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_72; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_73; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_74; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_75; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_76; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_77; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_78; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_79; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_80; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_81; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_82; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_83; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_84; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_85; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_86; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_87; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_88; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_89; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_90; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_91; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_92; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_93; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_94; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_95; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_96; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_97; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_98; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_99; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_100; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_101; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_102; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_103; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_104; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_105; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_106; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_107; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_108; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_109; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_110; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_111; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_112; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_113; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_114; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_115; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_116; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_117; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_118; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_119; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_120; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_121; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_122; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_123; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_124; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_125; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_126; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_127; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_128; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_129; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_130; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_131; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_132; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_133; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_134; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_135; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_136; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_137; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_138; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_139; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_140; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_141; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_142; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_143; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_144; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_145; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_146; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_147; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_148; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_149; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_150; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_151; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_152; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_153; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_154; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_155; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_156; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_157; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_158; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_159; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_out_header_0; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_out_header_1; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_out_header_2; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_out_header_3; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_out_header_4; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_out_header_5; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_out_header_6; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_out_header_7; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_out_header_8; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_out_header_9; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_out_header_10; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_out_header_11; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_out_header_12; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_out_header_13; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_out_header_14; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_out_header_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 79:25]
  wire [3:0] trans_0_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 79:25]
  wire  trans_0_io_pipe_phv_out_next_config_id; // @[ipsa.scala 79:25]
  wire  trans_0_io_pipe_phv_out_is_valid_processor; // @[ipsa.scala 79:25]
  wire  trans_0_io_pipe_phv_out_valid; // @[ipsa.scala 79:25]
  wire  trans_0_io_pipe_phv_out_last; // @[ipsa.scala 79:25]
  wire  trans_0_io_next_proc_exist; // @[ipsa.scala 79:25]
  wire  trans_1_clock; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_0; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_1; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_2; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_3; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_4; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_5; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_6; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_7; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_8; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_9; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_10; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_11; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_12; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_13; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_14; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_16; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_17; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_18; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_19; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_20; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_21; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_22; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_23; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_24; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_25; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_26; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_27; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_28; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_29; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_30; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_31; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_32; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_33; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_34; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_35; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_36; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_37; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_38; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_39; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_40; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_41; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_42; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_43; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_44; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_45; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_46; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_47; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_48; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_49; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_50; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_51; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_52; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_53; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_54; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_55; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_56; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_57; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_58; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_59; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_60; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_61; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_62; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_63; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_64; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_65; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_66; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_67; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_68; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_69; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_70; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_71; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_72; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_73; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_74; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_75; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_76; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_77; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_78; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_79; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_80; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_81; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_82; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_83; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_84; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_85; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_86; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_87; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_88; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_89; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_90; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_91; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_92; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_93; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_94; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_95; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_96; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_97; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_98; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_99; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_100; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_101; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_102; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_103; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_104; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_105; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_106; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_107; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_108; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_109; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_110; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_111; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_112; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_113; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_114; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_115; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_116; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_117; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_118; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_119; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_120; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_121; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_122; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_123; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_124; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_125; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_126; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_127; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_128; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_129; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_130; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_131; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_132; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_133; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_134; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_135; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_136; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_137; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_138; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_139; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_140; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_141; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_142; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_143; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_144; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_145; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_146; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_147; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_148; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_149; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_150; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_151; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_152; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_153; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_154; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_155; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_156; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_157; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_158; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_159; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_in_header_0; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_in_header_1; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_in_header_2; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_in_header_3; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_in_header_4; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_in_header_5; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_in_header_6; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_in_header_7; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_in_header_8; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_in_header_9; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_in_header_10; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_in_header_11; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_in_header_12; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_in_header_13; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_in_header_14; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_in_header_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_parse_current_state; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_parse_current_offset; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_in_parse_transition_field; // @[ipsa.scala 79:25]
  wire [3:0] trans_1_io_pipe_phv_in_next_processor_id; // @[ipsa.scala 79:25]
  wire  trans_1_io_pipe_phv_in_next_config_id; // @[ipsa.scala 79:25]
  wire  trans_1_io_pipe_phv_in_valid; // @[ipsa.scala 79:25]
  wire  trans_1_io_pipe_phv_in_last; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_0; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_1; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_2; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_3; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_4; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_5; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_6; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_7; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_8; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_9; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_10; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_11; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_12; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_13; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_14; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_16; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_17; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_18; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_19; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_20; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_21; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_22; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_23; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_24; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_25; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_26; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_27; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_28; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_29; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_30; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_31; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_32; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_33; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_34; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_35; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_36; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_37; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_38; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_39; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_40; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_41; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_42; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_43; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_44; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_45; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_46; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_47; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_48; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_49; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_50; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_51; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_52; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_53; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_54; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_55; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_56; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_57; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_58; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_59; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_60; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_61; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_62; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_63; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_64; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_65; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_66; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_67; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_68; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_69; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_70; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_71; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_72; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_73; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_74; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_75; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_76; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_77; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_78; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_79; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_80; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_81; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_82; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_83; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_84; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_85; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_86; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_87; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_88; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_89; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_90; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_91; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_92; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_93; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_94; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_95; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_96; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_97; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_98; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_99; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_100; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_101; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_102; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_103; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_104; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_105; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_106; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_107; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_108; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_109; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_110; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_111; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_112; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_113; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_114; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_115; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_116; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_117; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_118; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_119; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_120; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_121; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_122; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_123; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_124; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_125; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_126; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_127; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_128; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_129; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_130; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_131; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_132; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_133; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_134; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_135; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_136; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_137; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_138; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_139; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_140; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_141; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_142; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_143; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_144; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_145; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_146; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_147; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_148; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_149; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_150; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_151; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_152; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_153; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_154; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_155; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_156; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_157; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_158; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_159; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_out_header_0; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_out_header_1; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_out_header_2; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_out_header_3; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_out_header_4; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_out_header_5; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_out_header_6; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_out_header_7; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_out_header_8; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_out_header_9; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_out_header_10; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_out_header_11; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_out_header_12; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_out_header_13; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_out_header_14; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_out_header_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 79:25]
  wire [3:0] trans_1_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 79:25]
  wire  trans_1_io_pipe_phv_out_next_config_id; // @[ipsa.scala 79:25]
  wire  trans_1_io_pipe_phv_out_is_valid_processor; // @[ipsa.scala 79:25]
  wire  trans_1_io_pipe_phv_out_valid; // @[ipsa.scala 79:25]
  wire  trans_1_io_pipe_phv_out_last; // @[ipsa.scala 79:25]
  wire  trans_1_io_next_proc_exist; // @[ipsa.scala 79:25]
  wire  trans_2_clock; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_0; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_1; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_2; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_3; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_4; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_5; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_6; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_7; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_8; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_9; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_10; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_11; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_12; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_13; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_14; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_16; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_17; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_18; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_19; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_20; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_21; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_22; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_23; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_24; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_25; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_26; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_27; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_28; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_29; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_30; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_31; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_32; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_33; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_34; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_35; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_36; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_37; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_38; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_39; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_40; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_41; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_42; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_43; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_44; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_45; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_46; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_47; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_48; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_49; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_50; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_51; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_52; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_53; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_54; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_55; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_56; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_57; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_58; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_59; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_60; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_61; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_62; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_63; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_64; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_65; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_66; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_67; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_68; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_69; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_70; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_71; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_72; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_73; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_74; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_75; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_76; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_77; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_78; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_79; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_80; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_81; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_82; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_83; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_84; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_85; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_86; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_87; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_88; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_89; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_90; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_91; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_92; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_93; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_94; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_95; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_96; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_97; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_98; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_99; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_100; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_101; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_102; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_103; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_104; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_105; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_106; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_107; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_108; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_109; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_110; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_111; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_112; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_113; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_114; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_115; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_116; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_117; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_118; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_119; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_120; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_121; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_122; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_123; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_124; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_125; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_126; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_127; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_128; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_129; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_130; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_131; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_132; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_133; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_134; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_135; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_136; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_137; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_138; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_139; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_140; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_141; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_142; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_143; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_144; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_145; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_146; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_147; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_148; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_149; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_150; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_151; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_152; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_153; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_154; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_155; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_156; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_157; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_158; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_159; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_in_header_0; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_in_header_1; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_in_header_2; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_in_header_3; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_in_header_4; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_in_header_5; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_in_header_6; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_in_header_7; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_in_header_8; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_in_header_9; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_in_header_10; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_in_header_11; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_in_header_12; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_in_header_13; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_in_header_14; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_in_header_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_parse_current_state; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_parse_current_offset; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_in_parse_transition_field; // @[ipsa.scala 79:25]
  wire [3:0] trans_2_io_pipe_phv_in_next_processor_id; // @[ipsa.scala 79:25]
  wire  trans_2_io_pipe_phv_in_next_config_id; // @[ipsa.scala 79:25]
  wire  trans_2_io_pipe_phv_in_valid; // @[ipsa.scala 79:25]
  wire  trans_2_io_pipe_phv_in_last; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_0; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_1; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_2; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_3; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_4; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_5; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_6; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_7; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_8; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_9; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_10; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_11; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_12; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_13; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_14; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_16; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_17; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_18; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_19; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_20; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_21; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_22; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_23; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_24; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_25; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_26; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_27; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_28; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_29; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_30; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_31; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_32; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_33; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_34; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_35; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_36; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_37; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_38; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_39; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_40; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_41; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_42; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_43; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_44; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_45; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_46; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_47; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_48; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_49; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_50; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_51; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_52; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_53; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_54; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_55; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_56; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_57; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_58; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_59; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_60; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_61; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_62; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_63; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_64; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_65; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_66; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_67; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_68; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_69; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_70; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_71; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_72; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_73; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_74; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_75; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_76; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_77; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_78; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_79; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_80; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_81; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_82; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_83; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_84; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_85; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_86; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_87; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_88; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_89; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_90; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_91; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_92; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_93; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_94; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_95; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_96; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_97; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_98; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_99; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_100; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_101; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_102; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_103; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_104; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_105; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_106; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_107; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_108; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_109; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_110; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_111; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_112; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_113; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_114; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_115; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_116; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_117; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_118; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_119; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_120; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_121; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_122; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_123; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_124; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_125; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_126; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_127; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_128; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_129; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_130; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_131; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_132; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_133; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_134; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_135; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_136; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_137; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_138; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_139; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_140; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_141; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_142; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_143; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_144; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_145; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_146; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_147; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_148; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_149; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_150; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_151; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_152; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_153; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_154; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_155; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_156; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_157; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_158; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_159; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_out_header_0; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_out_header_1; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_out_header_2; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_out_header_3; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_out_header_4; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_out_header_5; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_out_header_6; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_out_header_7; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_out_header_8; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_out_header_9; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_out_header_10; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_out_header_11; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_out_header_12; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_out_header_13; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_out_header_14; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_out_header_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 79:25]
  wire [3:0] trans_2_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 79:25]
  wire  trans_2_io_pipe_phv_out_next_config_id; // @[ipsa.scala 79:25]
  wire  trans_2_io_pipe_phv_out_is_valid_processor; // @[ipsa.scala 79:25]
  wire  trans_2_io_pipe_phv_out_valid; // @[ipsa.scala 79:25]
  wire  trans_2_io_pipe_phv_out_last; // @[ipsa.scala 79:25]
  wire  trans_2_io_next_proc_exist; // @[ipsa.scala 79:25]
  wire  trans_3_clock; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_0; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_1; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_2; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_3; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_4; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_5; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_6; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_7; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_8; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_9; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_10; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_11; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_12; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_13; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_14; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_16; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_17; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_18; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_19; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_20; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_21; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_22; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_23; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_24; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_25; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_26; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_27; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_28; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_29; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_30; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_31; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_32; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_33; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_34; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_35; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_36; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_37; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_38; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_39; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_40; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_41; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_42; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_43; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_44; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_45; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_46; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_47; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_48; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_49; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_50; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_51; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_52; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_53; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_54; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_55; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_56; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_57; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_58; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_59; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_60; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_61; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_62; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_63; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_64; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_65; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_66; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_67; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_68; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_69; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_70; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_71; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_72; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_73; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_74; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_75; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_76; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_77; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_78; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_79; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_80; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_81; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_82; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_83; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_84; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_85; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_86; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_87; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_88; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_89; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_90; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_91; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_92; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_93; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_94; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_95; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_96; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_97; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_98; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_99; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_100; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_101; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_102; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_103; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_104; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_105; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_106; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_107; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_108; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_109; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_110; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_111; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_112; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_113; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_114; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_115; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_116; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_117; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_118; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_119; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_120; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_121; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_122; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_123; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_124; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_125; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_126; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_127; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_128; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_129; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_130; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_131; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_132; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_133; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_134; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_135; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_136; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_137; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_138; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_139; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_140; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_141; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_142; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_143; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_144; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_145; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_146; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_147; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_148; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_149; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_150; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_151; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_152; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_153; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_154; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_155; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_156; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_157; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_158; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_159; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_in_header_0; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_in_header_1; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_in_header_2; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_in_header_3; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_in_header_4; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_in_header_5; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_in_header_6; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_in_header_7; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_in_header_8; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_in_header_9; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_in_header_10; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_in_header_11; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_in_header_12; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_in_header_13; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_in_header_14; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_in_header_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_parse_current_state; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_parse_current_offset; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_in_parse_transition_field; // @[ipsa.scala 79:25]
  wire [3:0] trans_3_io_pipe_phv_in_next_processor_id; // @[ipsa.scala 79:25]
  wire  trans_3_io_pipe_phv_in_next_config_id; // @[ipsa.scala 79:25]
  wire  trans_3_io_pipe_phv_in_valid; // @[ipsa.scala 79:25]
  wire  trans_3_io_pipe_phv_in_last; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_0; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_1; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_2; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_3; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_4; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_5; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_6; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_7; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_8; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_9; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_10; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_11; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_12; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_13; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_14; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_16; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_17; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_18; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_19; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_20; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_21; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_22; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_23; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_24; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_25; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_26; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_27; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_28; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_29; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_30; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_31; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_32; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_33; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_34; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_35; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_36; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_37; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_38; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_39; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_40; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_41; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_42; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_43; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_44; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_45; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_46; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_47; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_48; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_49; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_50; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_51; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_52; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_53; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_54; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_55; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_56; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_57; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_58; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_59; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_60; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_61; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_62; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_63; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_64; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_65; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_66; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_67; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_68; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_69; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_70; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_71; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_72; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_73; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_74; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_75; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_76; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_77; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_78; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_79; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_80; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_81; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_82; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_83; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_84; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_85; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_86; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_87; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_88; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_89; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_90; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_91; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_92; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_93; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_94; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_95; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_96; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_97; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_98; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_99; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_100; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_101; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_102; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_103; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_104; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_105; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_106; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_107; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_108; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_109; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_110; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_111; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_112; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_113; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_114; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_115; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_116; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_117; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_118; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_119; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_120; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_121; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_122; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_123; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_124; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_125; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_126; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_127; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_128; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_129; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_130; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_131; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_132; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_133; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_134; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_135; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_136; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_137; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_138; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_139; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_140; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_141; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_142; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_143; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_144; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_145; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_146; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_147; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_148; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_149; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_150; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_151; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_152; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_153; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_154; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_155; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_156; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_157; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_158; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_159; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_out_header_0; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_out_header_1; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_out_header_2; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_out_header_3; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_out_header_4; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_out_header_5; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_out_header_6; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_out_header_7; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_out_header_8; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_out_header_9; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_out_header_10; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_out_header_11; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_out_header_12; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_out_header_13; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_out_header_14; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_out_header_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 79:25]
  wire [3:0] trans_3_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 79:25]
  wire  trans_3_io_pipe_phv_out_next_config_id; // @[ipsa.scala 79:25]
  wire  trans_3_io_pipe_phv_out_is_valid_processor; // @[ipsa.scala 79:25]
  wire  trans_3_io_pipe_phv_out_valid; // @[ipsa.scala 79:25]
  wire  trans_3_io_pipe_phv_out_last; // @[ipsa.scala 79:25]
  wire  trans_3_io_next_proc_exist; // @[ipsa.scala 79:25]
  wire  trans_4_clock; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_0; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_1; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_2; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_3; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_4; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_5; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_6; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_7; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_8; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_9; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_10; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_11; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_12; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_13; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_14; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_16; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_17; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_18; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_19; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_20; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_21; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_22; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_23; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_24; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_25; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_26; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_27; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_28; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_29; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_30; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_31; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_32; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_33; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_34; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_35; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_36; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_37; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_38; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_39; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_40; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_41; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_42; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_43; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_44; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_45; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_46; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_47; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_48; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_49; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_50; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_51; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_52; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_53; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_54; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_55; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_56; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_57; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_58; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_59; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_60; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_61; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_62; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_63; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_64; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_65; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_66; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_67; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_68; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_69; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_70; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_71; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_72; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_73; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_74; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_75; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_76; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_77; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_78; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_79; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_80; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_81; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_82; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_83; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_84; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_85; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_86; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_87; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_88; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_89; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_90; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_91; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_92; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_93; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_94; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_95; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_96; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_97; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_98; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_99; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_100; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_101; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_102; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_103; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_104; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_105; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_106; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_107; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_108; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_109; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_110; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_111; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_112; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_113; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_114; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_115; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_116; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_117; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_118; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_119; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_120; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_121; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_122; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_123; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_124; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_125; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_126; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_127; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_128; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_129; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_130; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_131; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_132; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_133; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_134; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_135; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_136; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_137; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_138; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_139; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_140; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_141; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_142; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_143; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_144; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_145; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_146; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_147; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_148; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_149; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_150; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_151; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_152; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_153; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_154; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_155; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_156; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_157; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_158; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_data_159; // @[ipsa.scala 79:25]
  wire [15:0] trans_4_io_pipe_phv_in_header_0; // @[ipsa.scala 79:25]
  wire [15:0] trans_4_io_pipe_phv_in_header_1; // @[ipsa.scala 79:25]
  wire [15:0] trans_4_io_pipe_phv_in_header_2; // @[ipsa.scala 79:25]
  wire [15:0] trans_4_io_pipe_phv_in_header_3; // @[ipsa.scala 79:25]
  wire [15:0] trans_4_io_pipe_phv_in_header_4; // @[ipsa.scala 79:25]
  wire [15:0] trans_4_io_pipe_phv_in_header_5; // @[ipsa.scala 79:25]
  wire [15:0] trans_4_io_pipe_phv_in_header_6; // @[ipsa.scala 79:25]
  wire [15:0] trans_4_io_pipe_phv_in_header_7; // @[ipsa.scala 79:25]
  wire [15:0] trans_4_io_pipe_phv_in_header_8; // @[ipsa.scala 79:25]
  wire [15:0] trans_4_io_pipe_phv_in_header_9; // @[ipsa.scala 79:25]
  wire [15:0] trans_4_io_pipe_phv_in_header_10; // @[ipsa.scala 79:25]
  wire [15:0] trans_4_io_pipe_phv_in_header_11; // @[ipsa.scala 79:25]
  wire [15:0] trans_4_io_pipe_phv_in_header_12; // @[ipsa.scala 79:25]
  wire [15:0] trans_4_io_pipe_phv_in_header_13; // @[ipsa.scala 79:25]
  wire [15:0] trans_4_io_pipe_phv_in_header_14; // @[ipsa.scala 79:25]
  wire [15:0] trans_4_io_pipe_phv_in_header_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_parse_current_state; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_in_parse_current_offset; // @[ipsa.scala 79:25]
  wire [15:0] trans_4_io_pipe_phv_in_parse_transition_field; // @[ipsa.scala 79:25]
  wire [3:0] trans_4_io_pipe_phv_in_next_processor_id; // @[ipsa.scala 79:25]
  wire  trans_4_io_pipe_phv_in_next_config_id; // @[ipsa.scala 79:25]
  wire  trans_4_io_pipe_phv_in_valid; // @[ipsa.scala 79:25]
  wire  trans_4_io_pipe_phv_in_last; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_0; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_1; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_2; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_3; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_4; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_5; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_6; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_7; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_8; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_9; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_10; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_11; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_12; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_13; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_14; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_16; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_17; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_18; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_19; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_20; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_21; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_22; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_23; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_24; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_25; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_26; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_27; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_28; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_29; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_30; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_31; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_32; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_33; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_34; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_35; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_36; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_37; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_38; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_39; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_40; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_41; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_42; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_43; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_44; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_45; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_46; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_47; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_48; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_49; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_50; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_51; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_52; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_53; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_54; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_55; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_56; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_57; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_58; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_59; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_60; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_61; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_62; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_63; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_64; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_65; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_66; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_67; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_68; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_69; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_70; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_71; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_72; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_73; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_74; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_75; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_76; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_77; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_78; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_79; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_80; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_81; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_82; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_83; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_84; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_85; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_86; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_87; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_88; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_89; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_90; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_91; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_92; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_93; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_94; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_95; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_96; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_97; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_98; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_99; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_100; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_101; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_102; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_103; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_104; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_105; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_106; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_107; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_108; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_109; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_110; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_111; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_112; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_113; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_114; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_115; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_116; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_117; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_118; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_119; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_120; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_121; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_122; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_123; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_124; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_125; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_126; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_127; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_128; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_129; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_130; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_131; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_132; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_133; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_134; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_135; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_136; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_137; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_138; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_139; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_140; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_141; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_142; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_143; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_144; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_145; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_146; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_147; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_148; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_149; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_150; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_151; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_152; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_153; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_154; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_155; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_156; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_157; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_158; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_data_159; // @[ipsa.scala 79:25]
  wire [15:0] trans_4_io_pipe_phv_out_header_0; // @[ipsa.scala 79:25]
  wire [15:0] trans_4_io_pipe_phv_out_header_1; // @[ipsa.scala 79:25]
  wire [15:0] trans_4_io_pipe_phv_out_header_2; // @[ipsa.scala 79:25]
  wire [15:0] trans_4_io_pipe_phv_out_header_3; // @[ipsa.scala 79:25]
  wire [15:0] trans_4_io_pipe_phv_out_header_4; // @[ipsa.scala 79:25]
  wire [15:0] trans_4_io_pipe_phv_out_header_5; // @[ipsa.scala 79:25]
  wire [15:0] trans_4_io_pipe_phv_out_header_6; // @[ipsa.scala 79:25]
  wire [15:0] trans_4_io_pipe_phv_out_header_7; // @[ipsa.scala 79:25]
  wire [15:0] trans_4_io_pipe_phv_out_header_8; // @[ipsa.scala 79:25]
  wire [15:0] trans_4_io_pipe_phv_out_header_9; // @[ipsa.scala 79:25]
  wire [15:0] trans_4_io_pipe_phv_out_header_10; // @[ipsa.scala 79:25]
  wire [15:0] trans_4_io_pipe_phv_out_header_11; // @[ipsa.scala 79:25]
  wire [15:0] trans_4_io_pipe_phv_out_header_12; // @[ipsa.scala 79:25]
  wire [15:0] trans_4_io_pipe_phv_out_header_13; // @[ipsa.scala 79:25]
  wire [15:0] trans_4_io_pipe_phv_out_header_14; // @[ipsa.scala 79:25]
  wire [15:0] trans_4_io_pipe_phv_out_header_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 79:25]
  wire [7:0] trans_4_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 79:25]
  wire [15:0] trans_4_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 79:25]
  wire [3:0] trans_4_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 79:25]
  wire  trans_4_io_pipe_phv_out_next_config_id; // @[ipsa.scala 79:25]
  wire  trans_4_io_pipe_phv_out_is_valid_processor; // @[ipsa.scala 79:25]
  wire  trans_4_io_pipe_phv_out_valid; // @[ipsa.scala 79:25]
  wire  trans_4_io_pipe_phv_out_last; // @[ipsa.scala 79:25]
  wire  trans_4_io_next_proc_exist; // @[ipsa.scala 79:25]
  wire  trans_5_clock; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_0; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_1; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_2; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_3; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_4; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_5; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_6; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_7; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_8; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_9; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_10; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_11; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_12; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_13; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_14; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_16; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_17; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_18; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_19; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_20; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_21; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_22; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_23; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_24; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_25; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_26; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_27; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_28; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_29; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_30; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_31; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_32; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_33; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_34; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_35; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_36; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_37; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_38; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_39; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_40; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_41; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_42; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_43; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_44; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_45; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_46; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_47; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_48; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_49; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_50; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_51; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_52; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_53; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_54; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_55; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_56; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_57; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_58; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_59; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_60; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_61; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_62; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_63; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_64; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_65; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_66; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_67; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_68; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_69; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_70; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_71; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_72; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_73; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_74; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_75; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_76; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_77; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_78; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_79; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_80; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_81; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_82; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_83; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_84; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_85; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_86; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_87; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_88; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_89; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_90; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_91; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_92; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_93; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_94; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_95; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_96; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_97; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_98; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_99; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_100; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_101; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_102; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_103; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_104; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_105; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_106; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_107; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_108; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_109; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_110; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_111; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_112; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_113; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_114; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_115; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_116; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_117; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_118; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_119; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_120; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_121; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_122; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_123; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_124; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_125; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_126; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_127; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_128; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_129; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_130; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_131; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_132; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_133; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_134; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_135; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_136; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_137; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_138; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_139; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_140; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_141; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_142; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_143; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_144; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_145; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_146; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_147; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_148; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_149; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_150; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_151; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_152; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_153; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_154; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_155; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_156; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_157; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_158; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_data_159; // @[ipsa.scala 79:25]
  wire [15:0] trans_5_io_pipe_phv_in_header_0; // @[ipsa.scala 79:25]
  wire [15:0] trans_5_io_pipe_phv_in_header_1; // @[ipsa.scala 79:25]
  wire [15:0] trans_5_io_pipe_phv_in_header_2; // @[ipsa.scala 79:25]
  wire [15:0] trans_5_io_pipe_phv_in_header_3; // @[ipsa.scala 79:25]
  wire [15:0] trans_5_io_pipe_phv_in_header_4; // @[ipsa.scala 79:25]
  wire [15:0] trans_5_io_pipe_phv_in_header_5; // @[ipsa.scala 79:25]
  wire [15:0] trans_5_io_pipe_phv_in_header_6; // @[ipsa.scala 79:25]
  wire [15:0] trans_5_io_pipe_phv_in_header_7; // @[ipsa.scala 79:25]
  wire [15:0] trans_5_io_pipe_phv_in_header_8; // @[ipsa.scala 79:25]
  wire [15:0] trans_5_io_pipe_phv_in_header_9; // @[ipsa.scala 79:25]
  wire [15:0] trans_5_io_pipe_phv_in_header_10; // @[ipsa.scala 79:25]
  wire [15:0] trans_5_io_pipe_phv_in_header_11; // @[ipsa.scala 79:25]
  wire [15:0] trans_5_io_pipe_phv_in_header_12; // @[ipsa.scala 79:25]
  wire [15:0] trans_5_io_pipe_phv_in_header_13; // @[ipsa.scala 79:25]
  wire [15:0] trans_5_io_pipe_phv_in_header_14; // @[ipsa.scala 79:25]
  wire [15:0] trans_5_io_pipe_phv_in_header_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_parse_current_state; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_in_parse_current_offset; // @[ipsa.scala 79:25]
  wire [15:0] trans_5_io_pipe_phv_in_parse_transition_field; // @[ipsa.scala 79:25]
  wire [3:0] trans_5_io_pipe_phv_in_next_processor_id; // @[ipsa.scala 79:25]
  wire  trans_5_io_pipe_phv_in_next_config_id; // @[ipsa.scala 79:25]
  wire  trans_5_io_pipe_phv_in_valid; // @[ipsa.scala 79:25]
  wire  trans_5_io_pipe_phv_in_last; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_0; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_1; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_2; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_3; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_4; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_5; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_6; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_7; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_8; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_9; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_10; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_11; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_12; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_13; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_14; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_16; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_17; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_18; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_19; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_20; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_21; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_22; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_23; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_24; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_25; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_26; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_27; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_28; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_29; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_30; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_31; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_32; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_33; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_34; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_35; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_36; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_37; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_38; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_39; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_40; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_41; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_42; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_43; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_44; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_45; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_46; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_47; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_48; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_49; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_50; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_51; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_52; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_53; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_54; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_55; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_56; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_57; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_58; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_59; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_60; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_61; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_62; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_63; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_64; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_65; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_66; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_67; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_68; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_69; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_70; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_71; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_72; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_73; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_74; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_75; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_76; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_77; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_78; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_79; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_80; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_81; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_82; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_83; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_84; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_85; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_86; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_87; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_88; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_89; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_90; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_91; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_92; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_93; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_94; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_95; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_96; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_97; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_98; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_99; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_100; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_101; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_102; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_103; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_104; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_105; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_106; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_107; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_108; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_109; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_110; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_111; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_112; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_113; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_114; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_115; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_116; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_117; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_118; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_119; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_120; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_121; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_122; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_123; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_124; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_125; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_126; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_127; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_128; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_129; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_130; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_131; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_132; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_133; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_134; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_135; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_136; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_137; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_138; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_139; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_140; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_141; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_142; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_143; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_144; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_145; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_146; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_147; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_148; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_149; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_150; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_151; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_152; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_153; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_154; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_155; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_156; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_157; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_158; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_data_159; // @[ipsa.scala 79:25]
  wire [15:0] trans_5_io_pipe_phv_out_header_0; // @[ipsa.scala 79:25]
  wire [15:0] trans_5_io_pipe_phv_out_header_1; // @[ipsa.scala 79:25]
  wire [15:0] trans_5_io_pipe_phv_out_header_2; // @[ipsa.scala 79:25]
  wire [15:0] trans_5_io_pipe_phv_out_header_3; // @[ipsa.scala 79:25]
  wire [15:0] trans_5_io_pipe_phv_out_header_4; // @[ipsa.scala 79:25]
  wire [15:0] trans_5_io_pipe_phv_out_header_5; // @[ipsa.scala 79:25]
  wire [15:0] trans_5_io_pipe_phv_out_header_6; // @[ipsa.scala 79:25]
  wire [15:0] trans_5_io_pipe_phv_out_header_7; // @[ipsa.scala 79:25]
  wire [15:0] trans_5_io_pipe_phv_out_header_8; // @[ipsa.scala 79:25]
  wire [15:0] trans_5_io_pipe_phv_out_header_9; // @[ipsa.scala 79:25]
  wire [15:0] trans_5_io_pipe_phv_out_header_10; // @[ipsa.scala 79:25]
  wire [15:0] trans_5_io_pipe_phv_out_header_11; // @[ipsa.scala 79:25]
  wire [15:0] trans_5_io_pipe_phv_out_header_12; // @[ipsa.scala 79:25]
  wire [15:0] trans_5_io_pipe_phv_out_header_13; // @[ipsa.scala 79:25]
  wire [15:0] trans_5_io_pipe_phv_out_header_14; // @[ipsa.scala 79:25]
  wire [15:0] trans_5_io_pipe_phv_out_header_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 79:25]
  wire [7:0] trans_5_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 79:25]
  wire [15:0] trans_5_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 79:25]
  wire [3:0] trans_5_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 79:25]
  wire  trans_5_io_pipe_phv_out_next_config_id; // @[ipsa.scala 79:25]
  wire  trans_5_io_pipe_phv_out_is_valid_processor; // @[ipsa.scala 79:25]
  wire  trans_5_io_pipe_phv_out_valid; // @[ipsa.scala 79:25]
  wire  trans_5_io_pipe_phv_out_last; // @[ipsa.scala 79:25]
  wire  trans_5_io_next_proc_exist; // @[ipsa.scala 79:25]
  wire  trans_6_clock; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_0; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_1; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_2; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_3; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_4; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_5; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_6; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_7; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_8; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_9; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_10; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_11; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_12; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_13; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_14; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_16; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_17; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_18; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_19; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_20; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_21; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_22; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_23; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_24; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_25; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_26; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_27; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_28; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_29; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_30; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_31; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_32; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_33; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_34; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_35; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_36; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_37; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_38; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_39; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_40; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_41; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_42; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_43; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_44; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_45; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_46; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_47; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_48; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_49; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_50; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_51; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_52; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_53; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_54; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_55; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_56; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_57; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_58; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_59; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_60; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_61; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_62; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_63; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_64; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_65; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_66; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_67; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_68; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_69; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_70; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_71; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_72; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_73; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_74; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_75; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_76; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_77; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_78; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_79; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_80; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_81; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_82; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_83; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_84; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_85; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_86; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_87; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_88; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_89; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_90; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_91; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_92; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_93; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_94; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_95; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_96; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_97; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_98; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_99; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_100; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_101; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_102; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_103; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_104; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_105; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_106; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_107; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_108; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_109; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_110; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_111; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_112; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_113; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_114; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_115; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_116; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_117; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_118; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_119; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_120; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_121; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_122; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_123; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_124; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_125; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_126; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_127; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_128; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_129; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_130; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_131; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_132; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_133; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_134; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_135; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_136; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_137; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_138; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_139; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_140; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_141; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_142; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_143; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_144; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_145; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_146; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_147; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_148; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_149; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_150; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_151; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_152; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_153; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_154; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_155; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_156; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_157; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_158; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_data_159; // @[ipsa.scala 79:25]
  wire [15:0] trans_6_io_pipe_phv_in_header_0; // @[ipsa.scala 79:25]
  wire [15:0] trans_6_io_pipe_phv_in_header_1; // @[ipsa.scala 79:25]
  wire [15:0] trans_6_io_pipe_phv_in_header_2; // @[ipsa.scala 79:25]
  wire [15:0] trans_6_io_pipe_phv_in_header_3; // @[ipsa.scala 79:25]
  wire [15:0] trans_6_io_pipe_phv_in_header_4; // @[ipsa.scala 79:25]
  wire [15:0] trans_6_io_pipe_phv_in_header_5; // @[ipsa.scala 79:25]
  wire [15:0] trans_6_io_pipe_phv_in_header_6; // @[ipsa.scala 79:25]
  wire [15:0] trans_6_io_pipe_phv_in_header_7; // @[ipsa.scala 79:25]
  wire [15:0] trans_6_io_pipe_phv_in_header_8; // @[ipsa.scala 79:25]
  wire [15:0] trans_6_io_pipe_phv_in_header_9; // @[ipsa.scala 79:25]
  wire [15:0] trans_6_io_pipe_phv_in_header_10; // @[ipsa.scala 79:25]
  wire [15:0] trans_6_io_pipe_phv_in_header_11; // @[ipsa.scala 79:25]
  wire [15:0] trans_6_io_pipe_phv_in_header_12; // @[ipsa.scala 79:25]
  wire [15:0] trans_6_io_pipe_phv_in_header_13; // @[ipsa.scala 79:25]
  wire [15:0] trans_6_io_pipe_phv_in_header_14; // @[ipsa.scala 79:25]
  wire [15:0] trans_6_io_pipe_phv_in_header_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_parse_current_state; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_in_parse_current_offset; // @[ipsa.scala 79:25]
  wire [15:0] trans_6_io_pipe_phv_in_parse_transition_field; // @[ipsa.scala 79:25]
  wire [3:0] trans_6_io_pipe_phv_in_next_processor_id; // @[ipsa.scala 79:25]
  wire  trans_6_io_pipe_phv_in_next_config_id; // @[ipsa.scala 79:25]
  wire  trans_6_io_pipe_phv_in_valid; // @[ipsa.scala 79:25]
  wire  trans_6_io_pipe_phv_in_last; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_0; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_1; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_2; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_3; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_4; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_5; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_6; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_7; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_8; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_9; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_10; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_11; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_12; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_13; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_14; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_16; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_17; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_18; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_19; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_20; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_21; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_22; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_23; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_24; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_25; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_26; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_27; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_28; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_29; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_30; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_31; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_32; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_33; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_34; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_35; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_36; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_37; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_38; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_39; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_40; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_41; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_42; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_43; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_44; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_45; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_46; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_47; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_48; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_49; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_50; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_51; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_52; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_53; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_54; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_55; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_56; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_57; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_58; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_59; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_60; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_61; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_62; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_63; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_64; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_65; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_66; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_67; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_68; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_69; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_70; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_71; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_72; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_73; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_74; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_75; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_76; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_77; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_78; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_79; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_80; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_81; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_82; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_83; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_84; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_85; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_86; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_87; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_88; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_89; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_90; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_91; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_92; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_93; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_94; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_95; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_96; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_97; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_98; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_99; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_100; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_101; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_102; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_103; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_104; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_105; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_106; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_107; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_108; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_109; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_110; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_111; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_112; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_113; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_114; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_115; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_116; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_117; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_118; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_119; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_120; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_121; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_122; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_123; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_124; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_125; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_126; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_127; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_128; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_129; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_130; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_131; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_132; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_133; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_134; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_135; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_136; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_137; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_138; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_139; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_140; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_141; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_142; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_143; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_144; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_145; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_146; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_147; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_148; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_149; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_150; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_151; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_152; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_153; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_154; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_155; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_156; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_157; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_158; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_data_159; // @[ipsa.scala 79:25]
  wire [15:0] trans_6_io_pipe_phv_out_header_0; // @[ipsa.scala 79:25]
  wire [15:0] trans_6_io_pipe_phv_out_header_1; // @[ipsa.scala 79:25]
  wire [15:0] trans_6_io_pipe_phv_out_header_2; // @[ipsa.scala 79:25]
  wire [15:0] trans_6_io_pipe_phv_out_header_3; // @[ipsa.scala 79:25]
  wire [15:0] trans_6_io_pipe_phv_out_header_4; // @[ipsa.scala 79:25]
  wire [15:0] trans_6_io_pipe_phv_out_header_5; // @[ipsa.scala 79:25]
  wire [15:0] trans_6_io_pipe_phv_out_header_6; // @[ipsa.scala 79:25]
  wire [15:0] trans_6_io_pipe_phv_out_header_7; // @[ipsa.scala 79:25]
  wire [15:0] trans_6_io_pipe_phv_out_header_8; // @[ipsa.scala 79:25]
  wire [15:0] trans_6_io_pipe_phv_out_header_9; // @[ipsa.scala 79:25]
  wire [15:0] trans_6_io_pipe_phv_out_header_10; // @[ipsa.scala 79:25]
  wire [15:0] trans_6_io_pipe_phv_out_header_11; // @[ipsa.scala 79:25]
  wire [15:0] trans_6_io_pipe_phv_out_header_12; // @[ipsa.scala 79:25]
  wire [15:0] trans_6_io_pipe_phv_out_header_13; // @[ipsa.scala 79:25]
  wire [15:0] trans_6_io_pipe_phv_out_header_14; // @[ipsa.scala 79:25]
  wire [15:0] trans_6_io_pipe_phv_out_header_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 79:25]
  wire [7:0] trans_6_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 79:25]
  wire [15:0] trans_6_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 79:25]
  wire [3:0] trans_6_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 79:25]
  wire  trans_6_io_pipe_phv_out_next_config_id; // @[ipsa.scala 79:25]
  wire  trans_6_io_pipe_phv_out_is_valid_processor; // @[ipsa.scala 79:25]
  wire  trans_6_io_pipe_phv_out_valid; // @[ipsa.scala 79:25]
  wire  trans_6_io_pipe_phv_out_last; // @[ipsa.scala 79:25]
  wire  trans_6_io_next_proc_exist; // @[ipsa.scala 79:25]
  wire  trans_7_clock; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_0; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_1; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_2; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_3; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_4; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_5; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_6; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_7; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_8; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_9; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_10; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_11; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_12; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_13; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_14; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_16; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_17; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_18; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_19; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_20; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_21; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_22; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_23; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_24; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_25; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_26; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_27; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_28; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_29; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_30; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_31; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_32; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_33; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_34; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_35; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_36; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_37; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_38; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_39; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_40; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_41; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_42; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_43; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_44; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_45; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_46; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_47; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_48; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_49; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_50; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_51; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_52; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_53; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_54; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_55; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_56; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_57; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_58; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_59; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_60; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_61; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_62; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_63; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_64; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_65; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_66; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_67; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_68; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_69; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_70; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_71; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_72; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_73; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_74; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_75; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_76; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_77; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_78; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_79; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_80; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_81; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_82; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_83; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_84; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_85; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_86; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_87; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_88; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_89; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_90; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_91; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_92; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_93; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_94; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_95; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_96; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_97; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_98; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_99; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_100; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_101; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_102; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_103; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_104; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_105; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_106; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_107; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_108; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_109; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_110; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_111; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_112; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_113; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_114; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_115; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_116; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_117; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_118; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_119; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_120; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_121; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_122; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_123; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_124; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_125; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_126; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_127; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_128; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_129; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_130; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_131; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_132; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_133; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_134; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_135; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_136; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_137; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_138; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_139; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_140; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_141; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_142; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_143; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_144; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_145; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_146; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_147; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_148; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_149; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_150; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_151; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_152; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_153; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_154; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_155; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_156; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_157; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_158; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_data_159; // @[ipsa.scala 79:25]
  wire [15:0] trans_7_io_pipe_phv_in_header_0; // @[ipsa.scala 79:25]
  wire [15:0] trans_7_io_pipe_phv_in_header_1; // @[ipsa.scala 79:25]
  wire [15:0] trans_7_io_pipe_phv_in_header_2; // @[ipsa.scala 79:25]
  wire [15:0] trans_7_io_pipe_phv_in_header_3; // @[ipsa.scala 79:25]
  wire [15:0] trans_7_io_pipe_phv_in_header_4; // @[ipsa.scala 79:25]
  wire [15:0] trans_7_io_pipe_phv_in_header_5; // @[ipsa.scala 79:25]
  wire [15:0] trans_7_io_pipe_phv_in_header_6; // @[ipsa.scala 79:25]
  wire [15:0] trans_7_io_pipe_phv_in_header_7; // @[ipsa.scala 79:25]
  wire [15:0] trans_7_io_pipe_phv_in_header_8; // @[ipsa.scala 79:25]
  wire [15:0] trans_7_io_pipe_phv_in_header_9; // @[ipsa.scala 79:25]
  wire [15:0] trans_7_io_pipe_phv_in_header_10; // @[ipsa.scala 79:25]
  wire [15:0] trans_7_io_pipe_phv_in_header_11; // @[ipsa.scala 79:25]
  wire [15:0] trans_7_io_pipe_phv_in_header_12; // @[ipsa.scala 79:25]
  wire [15:0] trans_7_io_pipe_phv_in_header_13; // @[ipsa.scala 79:25]
  wire [15:0] trans_7_io_pipe_phv_in_header_14; // @[ipsa.scala 79:25]
  wire [15:0] trans_7_io_pipe_phv_in_header_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_parse_current_state; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_in_parse_current_offset; // @[ipsa.scala 79:25]
  wire [15:0] trans_7_io_pipe_phv_in_parse_transition_field; // @[ipsa.scala 79:25]
  wire [3:0] trans_7_io_pipe_phv_in_next_processor_id; // @[ipsa.scala 79:25]
  wire  trans_7_io_pipe_phv_in_next_config_id; // @[ipsa.scala 79:25]
  wire  trans_7_io_pipe_phv_in_valid; // @[ipsa.scala 79:25]
  wire  trans_7_io_pipe_phv_in_last; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_0; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_1; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_2; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_3; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_4; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_5; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_6; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_7; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_8; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_9; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_10; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_11; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_12; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_13; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_14; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_16; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_17; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_18; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_19; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_20; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_21; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_22; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_23; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_24; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_25; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_26; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_27; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_28; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_29; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_30; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_31; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_32; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_33; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_34; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_35; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_36; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_37; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_38; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_39; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_40; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_41; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_42; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_43; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_44; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_45; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_46; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_47; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_48; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_49; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_50; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_51; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_52; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_53; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_54; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_55; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_56; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_57; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_58; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_59; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_60; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_61; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_62; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_63; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_64; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_65; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_66; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_67; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_68; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_69; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_70; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_71; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_72; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_73; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_74; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_75; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_76; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_77; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_78; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_79; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_80; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_81; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_82; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_83; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_84; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_85; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_86; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_87; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_88; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_89; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_90; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_91; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_92; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_93; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_94; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_95; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_96; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_97; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_98; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_99; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_100; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_101; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_102; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_103; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_104; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_105; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_106; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_107; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_108; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_109; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_110; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_111; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_112; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_113; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_114; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_115; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_116; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_117; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_118; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_119; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_120; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_121; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_122; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_123; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_124; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_125; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_126; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_127; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_128; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_129; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_130; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_131; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_132; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_133; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_134; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_135; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_136; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_137; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_138; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_139; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_140; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_141; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_142; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_143; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_144; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_145; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_146; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_147; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_148; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_149; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_150; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_151; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_152; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_153; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_154; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_155; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_156; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_157; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_158; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_data_159; // @[ipsa.scala 79:25]
  wire [15:0] trans_7_io_pipe_phv_out_header_0; // @[ipsa.scala 79:25]
  wire [15:0] trans_7_io_pipe_phv_out_header_1; // @[ipsa.scala 79:25]
  wire [15:0] trans_7_io_pipe_phv_out_header_2; // @[ipsa.scala 79:25]
  wire [15:0] trans_7_io_pipe_phv_out_header_3; // @[ipsa.scala 79:25]
  wire [15:0] trans_7_io_pipe_phv_out_header_4; // @[ipsa.scala 79:25]
  wire [15:0] trans_7_io_pipe_phv_out_header_5; // @[ipsa.scala 79:25]
  wire [15:0] trans_7_io_pipe_phv_out_header_6; // @[ipsa.scala 79:25]
  wire [15:0] trans_7_io_pipe_phv_out_header_7; // @[ipsa.scala 79:25]
  wire [15:0] trans_7_io_pipe_phv_out_header_8; // @[ipsa.scala 79:25]
  wire [15:0] trans_7_io_pipe_phv_out_header_9; // @[ipsa.scala 79:25]
  wire [15:0] trans_7_io_pipe_phv_out_header_10; // @[ipsa.scala 79:25]
  wire [15:0] trans_7_io_pipe_phv_out_header_11; // @[ipsa.scala 79:25]
  wire [15:0] trans_7_io_pipe_phv_out_header_12; // @[ipsa.scala 79:25]
  wire [15:0] trans_7_io_pipe_phv_out_header_13; // @[ipsa.scala 79:25]
  wire [15:0] trans_7_io_pipe_phv_out_header_14; // @[ipsa.scala 79:25]
  wire [15:0] trans_7_io_pipe_phv_out_header_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 79:25]
  wire [7:0] trans_7_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 79:25]
  wire [15:0] trans_7_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 79:25]
  wire [3:0] trans_7_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 79:25]
  wire  trans_7_io_pipe_phv_out_next_config_id; // @[ipsa.scala 79:25]
  wire  trans_7_io_pipe_phv_out_is_valid_processor; // @[ipsa.scala 79:25]
  wire  trans_7_io_pipe_phv_out_valid; // @[ipsa.scala 79:25]
  wire  trans_7_io_pipe_phv_out_last; // @[ipsa.scala 79:25]
  wire  trans_7_io_next_proc_exist; // @[ipsa.scala 79:25]
  wire  trans_8_clock; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_0; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_1; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_2; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_3; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_4; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_5; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_6; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_7; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_8; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_9; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_10; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_11; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_12; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_13; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_14; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_16; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_17; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_18; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_19; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_20; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_21; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_22; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_23; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_24; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_25; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_26; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_27; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_28; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_29; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_30; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_31; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_32; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_33; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_34; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_35; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_36; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_37; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_38; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_39; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_40; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_41; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_42; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_43; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_44; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_45; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_46; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_47; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_48; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_49; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_50; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_51; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_52; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_53; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_54; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_55; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_56; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_57; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_58; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_59; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_60; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_61; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_62; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_63; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_64; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_65; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_66; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_67; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_68; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_69; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_70; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_71; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_72; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_73; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_74; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_75; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_76; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_77; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_78; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_79; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_80; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_81; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_82; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_83; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_84; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_85; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_86; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_87; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_88; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_89; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_90; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_91; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_92; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_93; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_94; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_95; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_96; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_97; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_98; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_99; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_100; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_101; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_102; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_103; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_104; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_105; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_106; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_107; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_108; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_109; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_110; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_111; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_112; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_113; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_114; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_115; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_116; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_117; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_118; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_119; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_120; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_121; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_122; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_123; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_124; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_125; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_126; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_127; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_128; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_129; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_130; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_131; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_132; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_133; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_134; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_135; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_136; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_137; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_138; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_139; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_140; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_141; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_142; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_143; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_144; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_145; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_146; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_147; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_148; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_149; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_150; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_151; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_152; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_153; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_154; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_155; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_156; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_157; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_158; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_data_159; // @[ipsa.scala 79:25]
  wire [15:0] trans_8_io_pipe_phv_in_header_0; // @[ipsa.scala 79:25]
  wire [15:0] trans_8_io_pipe_phv_in_header_1; // @[ipsa.scala 79:25]
  wire [15:0] trans_8_io_pipe_phv_in_header_2; // @[ipsa.scala 79:25]
  wire [15:0] trans_8_io_pipe_phv_in_header_3; // @[ipsa.scala 79:25]
  wire [15:0] trans_8_io_pipe_phv_in_header_4; // @[ipsa.scala 79:25]
  wire [15:0] trans_8_io_pipe_phv_in_header_5; // @[ipsa.scala 79:25]
  wire [15:0] trans_8_io_pipe_phv_in_header_6; // @[ipsa.scala 79:25]
  wire [15:0] trans_8_io_pipe_phv_in_header_7; // @[ipsa.scala 79:25]
  wire [15:0] trans_8_io_pipe_phv_in_header_8; // @[ipsa.scala 79:25]
  wire [15:0] trans_8_io_pipe_phv_in_header_9; // @[ipsa.scala 79:25]
  wire [15:0] trans_8_io_pipe_phv_in_header_10; // @[ipsa.scala 79:25]
  wire [15:0] trans_8_io_pipe_phv_in_header_11; // @[ipsa.scala 79:25]
  wire [15:0] trans_8_io_pipe_phv_in_header_12; // @[ipsa.scala 79:25]
  wire [15:0] trans_8_io_pipe_phv_in_header_13; // @[ipsa.scala 79:25]
  wire [15:0] trans_8_io_pipe_phv_in_header_14; // @[ipsa.scala 79:25]
  wire [15:0] trans_8_io_pipe_phv_in_header_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_parse_current_state; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_in_parse_current_offset; // @[ipsa.scala 79:25]
  wire [15:0] trans_8_io_pipe_phv_in_parse_transition_field; // @[ipsa.scala 79:25]
  wire [3:0] trans_8_io_pipe_phv_in_next_processor_id; // @[ipsa.scala 79:25]
  wire  trans_8_io_pipe_phv_in_next_config_id; // @[ipsa.scala 79:25]
  wire  trans_8_io_pipe_phv_in_valid; // @[ipsa.scala 79:25]
  wire  trans_8_io_pipe_phv_in_last; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_0; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_1; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_2; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_3; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_4; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_5; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_6; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_7; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_8; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_9; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_10; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_11; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_12; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_13; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_14; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_16; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_17; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_18; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_19; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_20; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_21; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_22; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_23; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_24; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_25; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_26; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_27; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_28; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_29; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_30; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_31; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_32; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_33; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_34; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_35; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_36; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_37; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_38; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_39; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_40; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_41; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_42; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_43; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_44; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_45; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_46; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_47; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_48; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_49; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_50; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_51; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_52; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_53; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_54; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_55; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_56; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_57; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_58; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_59; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_60; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_61; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_62; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_63; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_64; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_65; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_66; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_67; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_68; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_69; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_70; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_71; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_72; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_73; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_74; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_75; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_76; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_77; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_78; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_79; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_80; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_81; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_82; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_83; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_84; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_85; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_86; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_87; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_88; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_89; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_90; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_91; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_92; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_93; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_94; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_95; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_96; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_97; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_98; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_99; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_100; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_101; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_102; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_103; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_104; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_105; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_106; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_107; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_108; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_109; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_110; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_111; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_112; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_113; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_114; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_115; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_116; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_117; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_118; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_119; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_120; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_121; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_122; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_123; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_124; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_125; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_126; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_127; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_128; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_129; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_130; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_131; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_132; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_133; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_134; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_135; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_136; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_137; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_138; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_139; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_140; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_141; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_142; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_143; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_144; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_145; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_146; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_147; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_148; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_149; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_150; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_151; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_152; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_153; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_154; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_155; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_156; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_157; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_158; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_data_159; // @[ipsa.scala 79:25]
  wire [15:0] trans_8_io_pipe_phv_out_header_0; // @[ipsa.scala 79:25]
  wire [15:0] trans_8_io_pipe_phv_out_header_1; // @[ipsa.scala 79:25]
  wire [15:0] trans_8_io_pipe_phv_out_header_2; // @[ipsa.scala 79:25]
  wire [15:0] trans_8_io_pipe_phv_out_header_3; // @[ipsa.scala 79:25]
  wire [15:0] trans_8_io_pipe_phv_out_header_4; // @[ipsa.scala 79:25]
  wire [15:0] trans_8_io_pipe_phv_out_header_5; // @[ipsa.scala 79:25]
  wire [15:0] trans_8_io_pipe_phv_out_header_6; // @[ipsa.scala 79:25]
  wire [15:0] trans_8_io_pipe_phv_out_header_7; // @[ipsa.scala 79:25]
  wire [15:0] trans_8_io_pipe_phv_out_header_8; // @[ipsa.scala 79:25]
  wire [15:0] trans_8_io_pipe_phv_out_header_9; // @[ipsa.scala 79:25]
  wire [15:0] trans_8_io_pipe_phv_out_header_10; // @[ipsa.scala 79:25]
  wire [15:0] trans_8_io_pipe_phv_out_header_11; // @[ipsa.scala 79:25]
  wire [15:0] trans_8_io_pipe_phv_out_header_12; // @[ipsa.scala 79:25]
  wire [15:0] trans_8_io_pipe_phv_out_header_13; // @[ipsa.scala 79:25]
  wire [15:0] trans_8_io_pipe_phv_out_header_14; // @[ipsa.scala 79:25]
  wire [15:0] trans_8_io_pipe_phv_out_header_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 79:25]
  wire [7:0] trans_8_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 79:25]
  wire [15:0] trans_8_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 79:25]
  wire [3:0] trans_8_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 79:25]
  wire  trans_8_io_pipe_phv_out_next_config_id; // @[ipsa.scala 79:25]
  wire  trans_8_io_pipe_phv_out_is_valid_processor; // @[ipsa.scala 79:25]
  wire  trans_8_io_pipe_phv_out_valid; // @[ipsa.scala 79:25]
  wire  trans_8_io_pipe_phv_out_last; // @[ipsa.scala 79:25]
  wire  trans_8_io_next_proc_exist; // @[ipsa.scala 79:25]
  wire  trans_9_clock; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_0; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_1; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_2; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_3; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_4; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_5; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_6; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_7; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_8; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_9; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_10; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_11; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_12; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_13; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_14; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_16; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_17; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_18; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_19; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_20; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_21; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_22; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_23; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_24; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_25; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_26; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_27; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_28; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_29; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_30; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_31; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_32; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_33; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_34; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_35; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_36; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_37; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_38; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_39; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_40; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_41; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_42; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_43; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_44; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_45; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_46; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_47; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_48; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_49; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_50; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_51; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_52; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_53; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_54; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_55; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_56; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_57; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_58; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_59; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_60; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_61; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_62; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_63; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_64; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_65; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_66; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_67; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_68; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_69; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_70; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_71; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_72; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_73; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_74; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_75; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_76; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_77; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_78; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_79; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_80; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_81; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_82; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_83; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_84; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_85; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_86; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_87; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_88; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_89; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_90; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_91; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_92; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_93; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_94; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_95; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_96; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_97; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_98; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_99; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_100; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_101; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_102; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_103; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_104; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_105; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_106; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_107; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_108; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_109; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_110; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_111; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_112; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_113; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_114; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_115; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_116; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_117; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_118; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_119; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_120; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_121; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_122; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_123; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_124; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_125; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_126; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_127; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_128; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_129; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_130; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_131; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_132; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_133; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_134; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_135; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_136; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_137; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_138; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_139; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_140; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_141; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_142; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_143; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_144; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_145; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_146; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_147; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_148; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_149; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_150; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_151; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_152; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_153; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_154; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_155; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_156; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_157; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_158; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_data_159; // @[ipsa.scala 79:25]
  wire [15:0] trans_9_io_pipe_phv_in_header_0; // @[ipsa.scala 79:25]
  wire [15:0] trans_9_io_pipe_phv_in_header_1; // @[ipsa.scala 79:25]
  wire [15:0] trans_9_io_pipe_phv_in_header_2; // @[ipsa.scala 79:25]
  wire [15:0] trans_9_io_pipe_phv_in_header_3; // @[ipsa.scala 79:25]
  wire [15:0] trans_9_io_pipe_phv_in_header_4; // @[ipsa.scala 79:25]
  wire [15:0] trans_9_io_pipe_phv_in_header_5; // @[ipsa.scala 79:25]
  wire [15:0] trans_9_io_pipe_phv_in_header_6; // @[ipsa.scala 79:25]
  wire [15:0] trans_9_io_pipe_phv_in_header_7; // @[ipsa.scala 79:25]
  wire [15:0] trans_9_io_pipe_phv_in_header_8; // @[ipsa.scala 79:25]
  wire [15:0] trans_9_io_pipe_phv_in_header_9; // @[ipsa.scala 79:25]
  wire [15:0] trans_9_io_pipe_phv_in_header_10; // @[ipsa.scala 79:25]
  wire [15:0] trans_9_io_pipe_phv_in_header_11; // @[ipsa.scala 79:25]
  wire [15:0] trans_9_io_pipe_phv_in_header_12; // @[ipsa.scala 79:25]
  wire [15:0] trans_9_io_pipe_phv_in_header_13; // @[ipsa.scala 79:25]
  wire [15:0] trans_9_io_pipe_phv_in_header_14; // @[ipsa.scala 79:25]
  wire [15:0] trans_9_io_pipe_phv_in_header_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_parse_current_state; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_in_parse_current_offset; // @[ipsa.scala 79:25]
  wire [15:0] trans_9_io_pipe_phv_in_parse_transition_field; // @[ipsa.scala 79:25]
  wire [3:0] trans_9_io_pipe_phv_in_next_processor_id; // @[ipsa.scala 79:25]
  wire  trans_9_io_pipe_phv_in_next_config_id; // @[ipsa.scala 79:25]
  wire  trans_9_io_pipe_phv_in_valid; // @[ipsa.scala 79:25]
  wire  trans_9_io_pipe_phv_in_last; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_0; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_1; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_2; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_3; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_4; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_5; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_6; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_7; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_8; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_9; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_10; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_11; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_12; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_13; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_14; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_16; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_17; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_18; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_19; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_20; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_21; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_22; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_23; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_24; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_25; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_26; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_27; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_28; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_29; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_30; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_31; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_32; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_33; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_34; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_35; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_36; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_37; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_38; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_39; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_40; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_41; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_42; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_43; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_44; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_45; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_46; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_47; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_48; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_49; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_50; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_51; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_52; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_53; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_54; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_55; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_56; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_57; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_58; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_59; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_60; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_61; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_62; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_63; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_64; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_65; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_66; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_67; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_68; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_69; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_70; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_71; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_72; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_73; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_74; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_75; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_76; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_77; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_78; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_79; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_80; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_81; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_82; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_83; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_84; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_85; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_86; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_87; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_88; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_89; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_90; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_91; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_92; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_93; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_94; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_95; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_96; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_97; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_98; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_99; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_100; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_101; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_102; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_103; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_104; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_105; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_106; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_107; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_108; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_109; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_110; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_111; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_112; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_113; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_114; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_115; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_116; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_117; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_118; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_119; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_120; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_121; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_122; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_123; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_124; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_125; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_126; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_127; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_128; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_129; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_130; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_131; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_132; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_133; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_134; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_135; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_136; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_137; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_138; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_139; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_140; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_141; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_142; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_143; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_144; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_145; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_146; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_147; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_148; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_149; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_150; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_151; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_152; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_153; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_154; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_155; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_156; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_157; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_158; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_data_159; // @[ipsa.scala 79:25]
  wire [15:0] trans_9_io_pipe_phv_out_header_0; // @[ipsa.scala 79:25]
  wire [15:0] trans_9_io_pipe_phv_out_header_1; // @[ipsa.scala 79:25]
  wire [15:0] trans_9_io_pipe_phv_out_header_2; // @[ipsa.scala 79:25]
  wire [15:0] trans_9_io_pipe_phv_out_header_3; // @[ipsa.scala 79:25]
  wire [15:0] trans_9_io_pipe_phv_out_header_4; // @[ipsa.scala 79:25]
  wire [15:0] trans_9_io_pipe_phv_out_header_5; // @[ipsa.scala 79:25]
  wire [15:0] trans_9_io_pipe_phv_out_header_6; // @[ipsa.scala 79:25]
  wire [15:0] trans_9_io_pipe_phv_out_header_7; // @[ipsa.scala 79:25]
  wire [15:0] trans_9_io_pipe_phv_out_header_8; // @[ipsa.scala 79:25]
  wire [15:0] trans_9_io_pipe_phv_out_header_9; // @[ipsa.scala 79:25]
  wire [15:0] trans_9_io_pipe_phv_out_header_10; // @[ipsa.scala 79:25]
  wire [15:0] trans_9_io_pipe_phv_out_header_11; // @[ipsa.scala 79:25]
  wire [15:0] trans_9_io_pipe_phv_out_header_12; // @[ipsa.scala 79:25]
  wire [15:0] trans_9_io_pipe_phv_out_header_13; // @[ipsa.scala 79:25]
  wire [15:0] trans_9_io_pipe_phv_out_header_14; // @[ipsa.scala 79:25]
  wire [15:0] trans_9_io_pipe_phv_out_header_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 79:25]
  wire [7:0] trans_9_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 79:25]
  wire [15:0] trans_9_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 79:25]
  wire [3:0] trans_9_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 79:25]
  wire  trans_9_io_pipe_phv_out_next_config_id; // @[ipsa.scala 79:25]
  wire  trans_9_io_pipe_phv_out_is_valid_processor; // @[ipsa.scala 79:25]
  wire  trans_9_io_pipe_phv_out_valid; // @[ipsa.scala 79:25]
  wire  trans_9_io_pipe_phv_out_last; // @[ipsa.scala 79:25]
  wire  trans_9_io_next_proc_exist; // @[ipsa.scala 79:25]
  wire  trans_10_clock; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_0; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_1; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_2; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_3; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_4; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_5; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_6; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_7; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_8; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_9; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_10; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_11; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_12; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_13; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_14; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_16; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_17; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_18; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_19; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_20; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_21; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_22; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_23; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_24; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_25; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_26; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_27; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_28; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_29; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_30; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_31; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_32; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_33; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_34; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_35; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_36; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_37; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_38; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_39; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_40; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_41; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_42; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_43; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_44; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_45; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_46; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_47; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_48; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_49; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_50; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_51; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_52; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_53; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_54; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_55; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_56; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_57; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_58; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_59; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_60; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_61; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_62; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_63; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_64; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_65; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_66; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_67; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_68; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_69; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_70; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_71; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_72; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_73; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_74; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_75; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_76; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_77; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_78; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_79; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_80; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_81; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_82; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_83; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_84; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_85; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_86; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_87; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_88; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_89; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_90; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_91; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_92; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_93; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_94; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_95; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_96; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_97; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_98; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_99; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_100; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_101; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_102; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_103; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_104; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_105; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_106; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_107; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_108; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_109; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_110; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_111; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_112; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_113; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_114; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_115; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_116; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_117; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_118; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_119; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_120; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_121; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_122; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_123; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_124; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_125; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_126; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_127; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_128; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_129; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_130; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_131; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_132; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_133; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_134; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_135; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_136; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_137; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_138; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_139; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_140; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_141; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_142; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_143; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_144; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_145; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_146; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_147; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_148; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_149; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_150; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_151; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_152; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_153; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_154; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_155; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_156; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_157; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_158; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_data_159; // @[ipsa.scala 79:25]
  wire [15:0] trans_10_io_pipe_phv_in_header_0; // @[ipsa.scala 79:25]
  wire [15:0] trans_10_io_pipe_phv_in_header_1; // @[ipsa.scala 79:25]
  wire [15:0] trans_10_io_pipe_phv_in_header_2; // @[ipsa.scala 79:25]
  wire [15:0] trans_10_io_pipe_phv_in_header_3; // @[ipsa.scala 79:25]
  wire [15:0] trans_10_io_pipe_phv_in_header_4; // @[ipsa.scala 79:25]
  wire [15:0] trans_10_io_pipe_phv_in_header_5; // @[ipsa.scala 79:25]
  wire [15:0] trans_10_io_pipe_phv_in_header_6; // @[ipsa.scala 79:25]
  wire [15:0] trans_10_io_pipe_phv_in_header_7; // @[ipsa.scala 79:25]
  wire [15:0] trans_10_io_pipe_phv_in_header_8; // @[ipsa.scala 79:25]
  wire [15:0] trans_10_io_pipe_phv_in_header_9; // @[ipsa.scala 79:25]
  wire [15:0] trans_10_io_pipe_phv_in_header_10; // @[ipsa.scala 79:25]
  wire [15:0] trans_10_io_pipe_phv_in_header_11; // @[ipsa.scala 79:25]
  wire [15:0] trans_10_io_pipe_phv_in_header_12; // @[ipsa.scala 79:25]
  wire [15:0] trans_10_io_pipe_phv_in_header_13; // @[ipsa.scala 79:25]
  wire [15:0] trans_10_io_pipe_phv_in_header_14; // @[ipsa.scala 79:25]
  wire [15:0] trans_10_io_pipe_phv_in_header_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_parse_current_state; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_in_parse_current_offset; // @[ipsa.scala 79:25]
  wire [15:0] trans_10_io_pipe_phv_in_parse_transition_field; // @[ipsa.scala 79:25]
  wire [3:0] trans_10_io_pipe_phv_in_next_processor_id; // @[ipsa.scala 79:25]
  wire  trans_10_io_pipe_phv_in_next_config_id; // @[ipsa.scala 79:25]
  wire  trans_10_io_pipe_phv_in_valid; // @[ipsa.scala 79:25]
  wire  trans_10_io_pipe_phv_in_last; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_0; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_1; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_2; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_3; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_4; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_5; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_6; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_7; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_8; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_9; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_10; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_11; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_12; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_13; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_14; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_16; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_17; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_18; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_19; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_20; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_21; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_22; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_23; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_24; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_25; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_26; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_27; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_28; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_29; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_30; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_31; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_32; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_33; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_34; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_35; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_36; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_37; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_38; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_39; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_40; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_41; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_42; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_43; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_44; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_45; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_46; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_47; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_48; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_49; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_50; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_51; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_52; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_53; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_54; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_55; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_56; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_57; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_58; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_59; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_60; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_61; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_62; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_63; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_64; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_65; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_66; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_67; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_68; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_69; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_70; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_71; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_72; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_73; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_74; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_75; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_76; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_77; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_78; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_79; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_80; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_81; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_82; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_83; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_84; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_85; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_86; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_87; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_88; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_89; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_90; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_91; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_92; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_93; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_94; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_95; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_96; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_97; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_98; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_99; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_100; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_101; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_102; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_103; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_104; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_105; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_106; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_107; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_108; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_109; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_110; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_111; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_112; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_113; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_114; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_115; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_116; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_117; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_118; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_119; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_120; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_121; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_122; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_123; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_124; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_125; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_126; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_127; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_128; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_129; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_130; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_131; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_132; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_133; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_134; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_135; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_136; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_137; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_138; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_139; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_140; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_141; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_142; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_143; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_144; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_145; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_146; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_147; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_148; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_149; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_150; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_151; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_152; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_153; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_154; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_155; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_156; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_157; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_158; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_data_159; // @[ipsa.scala 79:25]
  wire [15:0] trans_10_io_pipe_phv_out_header_0; // @[ipsa.scala 79:25]
  wire [15:0] trans_10_io_pipe_phv_out_header_1; // @[ipsa.scala 79:25]
  wire [15:0] trans_10_io_pipe_phv_out_header_2; // @[ipsa.scala 79:25]
  wire [15:0] trans_10_io_pipe_phv_out_header_3; // @[ipsa.scala 79:25]
  wire [15:0] trans_10_io_pipe_phv_out_header_4; // @[ipsa.scala 79:25]
  wire [15:0] trans_10_io_pipe_phv_out_header_5; // @[ipsa.scala 79:25]
  wire [15:0] trans_10_io_pipe_phv_out_header_6; // @[ipsa.scala 79:25]
  wire [15:0] trans_10_io_pipe_phv_out_header_7; // @[ipsa.scala 79:25]
  wire [15:0] trans_10_io_pipe_phv_out_header_8; // @[ipsa.scala 79:25]
  wire [15:0] trans_10_io_pipe_phv_out_header_9; // @[ipsa.scala 79:25]
  wire [15:0] trans_10_io_pipe_phv_out_header_10; // @[ipsa.scala 79:25]
  wire [15:0] trans_10_io_pipe_phv_out_header_11; // @[ipsa.scala 79:25]
  wire [15:0] trans_10_io_pipe_phv_out_header_12; // @[ipsa.scala 79:25]
  wire [15:0] trans_10_io_pipe_phv_out_header_13; // @[ipsa.scala 79:25]
  wire [15:0] trans_10_io_pipe_phv_out_header_14; // @[ipsa.scala 79:25]
  wire [15:0] trans_10_io_pipe_phv_out_header_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 79:25]
  wire [7:0] trans_10_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 79:25]
  wire [15:0] trans_10_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 79:25]
  wire [3:0] trans_10_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 79:25]
  wire  trans_10_io_pipe_phv_out_next_config_id; // @[ipsa.scala 79:25]
  wire  trans_10_io_pipe_phv_out_is_valid_processor; // @[ipsa.scala 79:25]
  wire  trans_10_io_pipe_phv_out_valid; // @[ipsa.scala 79:25]
  wire  trans_10_io_pipe_phv_out_last; // @[ipsa.scala 79:25]
  wire  trans_10_io_next_proc_exist; // @[ipsa.scala 79:25]
  wire  trans_11_clock; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_0; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_1; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_2; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_3; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_4; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_5; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_6; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_7; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_8; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_9; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_10; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_11; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_12; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_13; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_14; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_16; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_17; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_18; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_19; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_20; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_21; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_22; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_23; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_24; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_25; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_26; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_27; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_28; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_29; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_30; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_31; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_32; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_33; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_34; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_35; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_36; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_37; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_38; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_39; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_40; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_41; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_42; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_43; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_44; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_45; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_46; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_47; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_48; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_49; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_50; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_51; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_52; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_53; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_54; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_55; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_56; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_57; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_58; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_59; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_60; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_61; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_62; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_63; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_64; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_65; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_66; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_67; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_68; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_69; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_70; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_71; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_72; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_73; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_74; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_75; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_76; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_77; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_78; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_79; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_80; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_81; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_82; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_83; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_84; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_85; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_86; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_87; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_88; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_89; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_90; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_91; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_92; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_93; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_94; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_95; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_96; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_97; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_98; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_99; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_100; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_101; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_102; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_103; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_104; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_105; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_106; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_107; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_108; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_109; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_110; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_111; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_112; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_113; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_114; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_115; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_116; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_117; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_118; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_119; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_120; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_121; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_122; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_123; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_124; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_125; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_126; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_127; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_128; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_129; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_130; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_131; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_132; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_133; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_134; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_135; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_136; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_137; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_138; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_139; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_140; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_141; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_142; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_143; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_144; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_145; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_146; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_147; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_148; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_149; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_150; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_151; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_152; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_153; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_154; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_155; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_156; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_157; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_158; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_data_159; // @[ipsa.scala 79:25]
  wire [15:0] trans_11_io_pipe_phv_in_header_0; // @[ipsa.scala 79:25]
  wire [15:0] trans_11_io_pipe_phv_in_header_1; // @[ipsa.scala 79:25]
  wire [15:0] trans_11_io_pipe_phv_in_header_2; // @[ipsa.scala 79:25]
  wire [15:0] trans_11_io_pipe_phv_in_header_3; // @[ipsa.scala 79:25]
  wire [15:0] trans_11_io_pipe_phv_in_header_4; // @[ipsa.scala 79:25]
  wire [15:0] trans_11_io_pipe_phv_in_header_5; // @[ipsa.scala 79:25]
  wire [15:0] trans_11_io_pipe_phv_in_header_6; // @[ipsa.scala 79:25]
  wire [15:0] trans_11_io_pipe_phv_in_header_7; // @[ipsa.scala 79:25]
  wire [15:0] trans_11_io_pipe_phv_in_header_8; // @[ipsa.scala 79:25]
  wire [15:0] trans_11_io_pipe_phv_in_header_9; // @[ipsa.scala 79:25]
  wire [15:0] trans_11_io_pipe_phv_in_header_10; // @[ipsa.scala 79:25]
  wire [15:0] trans_11_io_pipe_phv_in_header_11; // @[ipsa.scala 79:25]
  wire [15:0] trans_11_io_pipe_phv_in_header_12; // @[ipsa.scala 79:25]
  wire [15:0] trans_11_io_pipe_phv_in_header_13; // @[ipsa.scala 79:25]
  wire [15:0] trans_11_io_pipe_phv_in_header_14; // @[ipsa.scala 79:25]
  wire [15:0] trans_11_io_pipe_phv_in_header_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_parse_current_state; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_in_parse_current_offset; // @[ipsa.scala 79:25]
  wire [15:0] trans_11_io_pipe_phv_in_parse_transition_field; // @[ipsa.scala 79:25]
  wire [3:0] trans_11_io_pipe_phv_in_next_processor_id; // @[ipsa.scala 79:25]
  wire  trans_11_io_pipe_phv_in_next_config_id; // @[ipsa.scala 79:25]
  wire  trans_11_io_pipe_phv_in_valid; // @[ipsa.scala 79:25]
  wire  trans_11_io_pipe_phv_in_last; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_0; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_1; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_2; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_3; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_4; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_5; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_6; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_7; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_8; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_9; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_10; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_11; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_12; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_13; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_14; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_16; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_17; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_18; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_19; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_20; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_21; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_22; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_23; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_24; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_25; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_26; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_27; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_28; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_29; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_30; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_31; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_32; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_33; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_34; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_35; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_36; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_37; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_38; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_39; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_40; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_41; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_42; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_43; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_44; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_45; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_46; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_47; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_48; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_49; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_50; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_51; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_52; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_53; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_54; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_55; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_56; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_57; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_58; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_59; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_60; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_61; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_62; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_63; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_64; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_65; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_66; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_67; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_68; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_69; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_70; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_71; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_72; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_73; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_74; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_75; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_76; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_77; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_78; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_79; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_80; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_81; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_82; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_83; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_84; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_85; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_86; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_87; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_88; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_89; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_90; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_91; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_92; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_93; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_94; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_95; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_96; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_97; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_98; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_99; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_100; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_101; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_102; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_103; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_104; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_105; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_106; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_107; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_108; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_109; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_110; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_111; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_112; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_113; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_114; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_115; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_116; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_117; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_118; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_119; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_120; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_121; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_122; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_123; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_124; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_125; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_126; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_127; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_128; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_129; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_130; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_131; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_132; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_133; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_134; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_135; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_136; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_137; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_138; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_139; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_140; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_141; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_142; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_143; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_144; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_145; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_146; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_147; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_148; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_149; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_150; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_151; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_152; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_153; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_154; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_155; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_156; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_157; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_158; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_data_159; // @[ipsa.scala 79:25]
  wire [15:0] trans_11_io_pipe_phv_out_header_0; // @[ipsa.scala 79:25]
  wire [15:0] trans_11_io_pipe_phv_out_header_1; // @[ipsa.scala 79:25]
  wire [15:0] trans_11_io_pipe_phv_out_header_2; // @[ipsa.scala 79:25]
  wire [15:0] trans_11_io_pipe_phv_out_header_3; // @[ipsa.scala 79:25]
  wire [15:0] trans_11_io_pipe_phv_out_header_4; // @[ipsa.scala 79:25]
  wire [15:0] trans_11_io_pipe_phv_out_header_5; // @[ipsa.scala 79:25]
  wire [15:0] trans_11_io_pipe_phv_out_header_6; // @[ipsa.scala 79:25]
  wire [15:0] trans_11_io_pipe_phv_out_header_7; // @[ipsa.scala 79:25]
  wire [15:0] trans_11_io_pipe_phv_out_header_8; // @[ipsa.scala 79:25]
  wire [15:0] trans_11_io_pipe_phv_out_header_9; // @[ipsa.scala 79:25]
  wire [15:0] trans_11_io_pipe_phv_out_header_10; // @[ipsa.scala 79:25]
  wire [15:0] trans_11_io_pipe_phv_out_header_11; // @[ipsa.scala 79:25]
  wire [15:0] trans_11_io_pipe_phv_out_header_12; // @[ipsa.scala 79:25]
  wire [15:0] trans_11_io_pipe_phv_out_header_13; // @[ipsa.scala 79:25]
  wire [15:0] trans_11_io_pipe_phv_out_header_14; // @[ipsa.scala 79:25]
  wire [15:0] trans_11_io_pipe_phv_out_header_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 79:25]
  wire [7:0] trans_11_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 79:25]
  wire [15:0] trans_11_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 79:25]
  wire [3:0] trans_11_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 79:25]
  wire  trans_11_io_pipe_phv_out_next_config_id; // @[ipsa.scala 79:25]
  wire  trans_11_io_pipe_phv_out_is_valid_processor; // @[ipsa.scala 79:25]
  wire  trans_11_io_pipe_phv_out_valid; // @[ipsa.scala 79:25]
  wire  trans_11_io_pipe_phv_out_last; // @[ipsa.scala 79:25]
  wire  trans_11_io_next_proc_exist; // @[ipsa.scala 79:25]
  wire  trans_12_clock; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_0; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_1; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_2; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_3; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_4; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_5; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_6; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_7; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_8; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_9; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_10; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_11; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_12; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_13; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_14; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_16; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_17; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_18; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_19; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_20; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_21; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_22; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_23; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_24; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_25; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_26; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_27; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_28; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_29; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_30; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_31; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_32; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_33; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_34; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_35; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_36; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_37; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_38; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_39; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_40; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_41; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_42; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_43; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_44; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_45; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_46; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_47; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_48; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_49; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_50; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_51; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_52; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_53; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_54; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_55; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_56; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_57; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_58; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_59; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_60; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_61; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_62; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_63; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_64; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_65; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_66; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_67; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_68; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_69; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_70; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_71; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_72; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_73; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_74; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_75; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_76; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_77; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_78; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_79; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_80; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_81; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_82; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_83; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_84; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_85; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_86; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_87; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_88; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_89; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_90; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_91; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_92; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_93; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_94; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_95; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_96; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_97; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_98; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_99; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_100; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_101; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_102; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_103; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_104; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_105; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_106; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_107; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_108; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_109; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_110; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_111; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_112; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_113; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_114; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_115; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_116; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_117; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_118; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_119; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_120; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_121; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_122; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_123; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_124; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_125; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_126; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_127; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_128; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_129; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_130; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_131; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_132; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_133; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_134; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_135; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_136; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_137; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_138; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_139; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_140; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_141; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_142; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_143; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_144; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_145; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_146; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_147; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_148; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_149; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_150; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_151; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_152; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_153; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_154; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_155; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_156; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_157; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_158; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_data_159; // @[ipsa.scala 79:25]
  wire [15:0] trans_12_io_pipe_phv_in_header_0; // @[ipsa.scala 79:25]
  wire [15:0] trans_12_io_pipe_phv_in_header_1; // @[ipsa.scala 79:25]
  wire [15:0] trans_12_io_pipe_phv_in_header_2; // @[ipsa.scala 79:25]
  wire [15:0] trans_12_io_pipe_phv_in_header_3; // @[ipsa.scala 79:25]
  wire [15:0] trans_12_io_pipe_phv_in_header_4; // @[ipsa.scala 79:25]
  wire [15:0] trans_12_io_pipe_phv_in_header_5; // @[ipsa.scala 79:25]
  wire [15:0] trans_12_io_pipe_phv_in_header_6; // @[ipsa.scala 79:25]
  wire [15:0] trans_12_io_pipe_phv_in_header_7; // @[ipsa.scala 79:25]
  wire [15:0] trans_12_io_pipe_phv_in_header_8; // @[ipsa.scala 79:25]
  wire [15:0] trans_12_io_pipe_phv_in_header_9; // @[ipsa.scala 79:25]
  wire [15:0] trans_12_io_pipe_phv_in_header_10; // @[ipsa.scala 79:25]
  wire [15:0] trans_12_io_pipe_phv_in_header_11; // @[ipsa.scala 79:25]
  wire [15:0] trans_12_io_pipe_phv_in_header_12; // @[ipsa.scala 79:25]
  wire [15:0] trans_12_io_pipe_phv_in_header_13; // @[ipsa.scala 79:25]
  wire [15:0] trans_12_io_pipe_phv_in_header_14; // @[ipsa.scala 79:25]
  wire [15:0] trans_12_io_pipe_phv_in_header_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_parse_current_state; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_in_parse_current_offset; // @[ipsa.scala 79:25]
  wire [15:0] trans_12_io_pipe_phv_in_parse_transition_field; // @[ipsa.scala 79:25]
  wire [3:0] trans_12_io_pipe_phv_in_next_processor_id; // @[ipsa.scala 79:25]
  wire  trans_12_io_pipe_phv_in_next_config_id; // @[ipsa.scala 79:25]
  wire  trans_12_io_pipe_phv_in_valid; // @[ipsa.scala 79:25]
  wire  trans_12_io_pipe_phv_in_last; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_0; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_1; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_2; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_3; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_4; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_5; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_6; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_7; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_8; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_9; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_10; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_11; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_12; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_13; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_14; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_16; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_17; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_18; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_19; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_20; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_21; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_22; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_23; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_24; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_25; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_26; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_27; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_28; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_29; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_30; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_31; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_32; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_33; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_34; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_35; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_36; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_37; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_38; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_39; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_40; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_41; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_42; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_43; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_44; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_45; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_46; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_47; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_48; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_49; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_50; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_51; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_52; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_53; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_54; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_55; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_56; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_57; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_58; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_59; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_60; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_61; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_62; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_63; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_64; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_65; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_66; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_67; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_68; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_69; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_70; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_71; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_72; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_73; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_74; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_75; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_76; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_77; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_78; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_79; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_80; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_81; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_82; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_83; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_84; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_85; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_86; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_87; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_88; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_89; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_90; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_91; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_92; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_93; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_94; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_95; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_96; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_97; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_98; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_99; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_100; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_101; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_102; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_103; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_104; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_105; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_106; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_107; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_108; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_109; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_110; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_111; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_112; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_113; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_114; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_115; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_116; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_117; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_118; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_119; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_120; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_121; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_122; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_123; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_124; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_125; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_126; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_127; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_128; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_129; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_130; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_131; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_132; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_133; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_134; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_135; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_136; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_137; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_138; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_139; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_140; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_141; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_142; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_143; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_144; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_145; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_146; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_147; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_148; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_149; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_150; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_151; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_152; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_153; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_154; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_155; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_156; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_157; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_158; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_data_159; // @[ipsa.scala 79:25]
  wire [15:0] trans_12_io_pipe_phv_out_header_0; // @[ipsa.scala 79:25]
  wire [15:0] trans_12_io_pipe_phv_out_header_1; // @[ipsa.scala 79:25]
  wire [15:0] trans_12_io_pipe_phv_out_header_2; // @[ipsa.scala 79:25]
  wire [15:0] trans_12_io_pipe_phv_out_header_3; // @[ipsa.scala 79:25]
  wire [15:0] trans_12_io_pipe_phv_out_header_4; // @[ipsa.scala 79:25]
  wire [15:0] trans_12_io_pipe_phv_out_header_5; // @[ipsa.scala 79:25]
  wire [15:0] trans_12_io_pipe_phv_out_header_6; // @[ipsa.scala 79:25]
  wire [15:0] trans_12_io_pipe_phv_out_header_7; // @[ipsa.scala 79:25]
  wire [15:0] trans_12_io_pipe_phv_out_header_8; // @[ipsa.scala 79:25]
  wire [15:0] trans_12_io_pipe_phv_out_header_9; // @[ipsa.scala 79:25]
  wire [15:0] trans_12_io_pipe_phv_out_header_10; // @[ipsa.scala 79:25]
  wire [15:0] trans_12_io_pipe_phv_out_header_11; // @[ipsa.scala 79:25]
  wire [15:0] trans_12_io_pipe_phv_out_header_12; // @[ipsa.scala 79:25]
  wire [15:0] trans_12_io_pipe_phv_out_header_13; // @[ipsa.scala 79:25]
  wire [15:0] trans_12_io_pipe_phv_out_header_14; // @[ipsa.scala 79:25]
  wire [15:0] trans_12_io_pipe_phv_out_header_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 79:25]
  wire [7:0] trans_12_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 79:25]
  wire [15:0] trans_12_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 79:25]
  wire [3:0] trans_12_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 79:25]
  wire  trans_12_io_pipe_phv_out_next_config_id; // @[ipsa.scala 79:25]
  wire  trans_12_io_pipe_phv_out_is_valid_processor; // @[ipsa.scala 79:25]
  wire  trans_12_io_pipe_phv_out_valid; // @[ipsa.scala 79:25]
  wire  trans_12_io_pipe_phv_out_last; // @[ipsa.scala 79:25]
  wire  trans_12_io_next_proc_exist; // @[ipsa.scala 79:25]
  wire  trans_13_clock; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_0; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_1; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_2; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_3; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_4; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_5; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_6; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_7; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_8; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_9; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_10; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_11; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_12; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_13; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_14; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_16; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_17; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_18; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_19; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_20; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_21; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_22; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_23; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_24; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_25; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_26; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_27; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_28; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_29; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_30; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_31; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_32; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_33; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_34; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_35; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_36; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_37; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_38; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_39; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_40; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_41; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_42; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_43; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_44; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_45; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_46; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_47; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_48; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_49; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_50; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_51; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_52; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_53; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_54; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_55; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_56; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_57; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_58; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_59; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_60; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_61; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_62; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_63; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_64; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_65; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_66; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_67; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_68; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_69; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_70; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_71; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_72; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_73; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_74; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_75; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_76; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_77; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_78; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_79; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_80; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_81; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_82; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_83; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_84; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_85; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_86; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_87; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_88; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_89; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_90; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_91; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_92; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_93; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_94; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_95; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_96; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_97; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_98; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_99; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_100; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_101; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_102; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_103; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_104; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_105; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_106; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_107; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_108; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_109; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_110; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_111; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_112; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_113; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_114; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_115; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_116; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_117; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_118; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_119; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_120; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_121; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_122; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_123; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_124; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_125; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_126; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_127; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_128; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_129; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_130; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_131; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_132; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_133; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_134; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_135; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_136; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_137; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_138; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_139; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_140; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_141; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_142; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_143; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_144; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_145; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_146; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_147; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_148; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_149; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_150; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_151; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_152; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_153; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_154; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_155; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_156; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_157; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_158; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_data_159; // @[ipsa.scala 79:25]
  wire [15:0] trans_13_io_pipe_phv_in_header_0; // @[ipsa.scala 79:25]
  wire [15:0] trans_13_io_pipe_phv_in_header_1; // @[ipsa.scala 79:25]
  wire [15:0] trans_13_io_pipe_phv_in_header_2; // @[ipsa.scala 79:25]
  wire [15:0] trans_13_io_pipe_phv_in_header_3; // @[ipsa.scala 79:25]
  wire [15:0] trans_13_io_pipe_phv_in_header_4; // @[ipsa.scala 79:25]
  wire [15:0] trans_13_io_pipe_phv_in_header_5; // @[ipsa.scala 79:25]
  wire [15:0] trans_13_io_pipe_phv_in_header_6; // @[ipsa.scala 79:25]
  wire [15:0] trans_13_io_pipe_phv_in_header_7; // @[ipsa.scala 79:25]
  wire [15:0] trans_13_io_pipe_phv_in_header_8; // @[ipsa.scala 79:25]
  wire [15:0] trans_13_io_pipe_phv_in_header_9; // @[ipsa.scala 79:25]
  wire [15:0] trans_13_io_pipe_phv_in_header_10; // @[ipsa.scala 79:25]
  wire [15:0] trans_13_io_pipe_phv_in_header_11; // @[ipsa.scala 79:25]
  wire [15:0] trans_13_io_pipe_phv_in_header_12; // @[ipsa.scala 79:25]
  wire [15:0] trans_13_io_pipe_phv_in_header_13; // @[ipsa.scala 79:25]
  wire [15:0] trans_13_io_pipe_phv_in_header_14; // @[ipsa.scala 79:25]
  wire [15:0] trans_13_io_pipe_phv_in_header_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_parse_current_state; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_in_parse_current_offset; // @[ipsa.scala 79:25]
  wire [15:0] trans_13_io_pipe_phv_in_parse_transition_field; // @[ipsa.scala 79:25]
  wire [3:0] trans_13_io_pipe_phv_in_next_processor_id; // @[ipsa.scala 79:25]
  wire  trans_13_io_pipe_phv_in_next_config_id; // @[ipsa.scala 79:25]
  wire  trans_13_io_pipe_phv_in_valid; // @[ipsa.scala 79:25]
  wire  trans_13_io_pipe_phv_in_last; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_0; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_1; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_2; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_3; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_4; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_5; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_6; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_7; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_8; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_9; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_10; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_11; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_12; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_13; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_14; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_16; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_17; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_18; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_19; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_20; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_21; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_22; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_23; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_24; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_25; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_26; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_27; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_28; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_29; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_30; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_31; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_32; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_33; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_34; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_35; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_36; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_37; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_38; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_39; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_40; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_41; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_42; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_43; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_44; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_45; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_46; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_47; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_48; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_49; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_50; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_51; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_52; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_53; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_54; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_55; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_56; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_57; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_58; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_59; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_60; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_61; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_62; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_63; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_64; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_65; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_66; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_67; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_68; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_69; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_70; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_71; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_72; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_73; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_74; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_75; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_76; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_77; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_78; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_79; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_80; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_81; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_82; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_83; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_84; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_85; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_86; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_87; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_88; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_89; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_90; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_91; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_92; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_93; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_94; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_95; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_96; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_97; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_98; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_99; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_100; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_101; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_102; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_103; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_104; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_105; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_106; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_107; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_108; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_109; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_110; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_111; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_112; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_113; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_114; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_115; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_116; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_117; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_118; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_119; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_120; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_121; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_122; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_123; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_124; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_125; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_126; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_127; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_128; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_129; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_130; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_131; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_132; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_133; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_134; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_135; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_136; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_137; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_138; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_139; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_140; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_141; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_142; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_143; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_144; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_145; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_146; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_147; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_148; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_149; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_150; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_151; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_152; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_153; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_154; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_155; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_156; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_157; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_158; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_data_159; // @[ipsa.scala 79:25]
  wire [15:0] trans_13_io_pipe_phv_out_header_0; // @[ipsa.scala 79:25]
  wire [15:0] trans_13_io_pipe_phv_out_header_1; // @[ipsa.scala 79:25]
  wire [15:0] trans_13_io_pipe_phv_out_header_2; // @[ipsa.scala 79:25]
  wire [15:0] trans_13_io_pipe_phv_out_header_3; // @[ipsa.scala 79:25]
  wire [15:0] trans_13_io_pipe_phv_out_header_4; // @[ipsa.scala 79:25]
  wire [15:0] trans_13_io_pipe_phv_out_header_5; // @[ipsa.scala 79:25]
  wire [15:0] trans_13_io_pipe_phv_out_header_6; // @[ipsa.scala 79:25]
  wire [15:0] trans_13_io_pipe_phv_out_header_7; // @[ipsa.scala 79:25]
  wire [15:0] trans_13_io_pipe_phv_out_header_8; // @[ipsa.scala 79:25]
  wire [15:0] trans_13_io_pipe_phv_out_header_9; // @[ipsa.scala 79:25]
  wire [15:0] trans_13_io_pipe_phv_out_header_10; // @[ipsa.scala 79:25]
  wire [15:0] trans_13_io_pipe_phv_out_header_11; // @[ipsa.scala 79:25]
  wire [15:0] trans_13_io_pipe_phv_out_header_12; // @[ipsa.scala 79:25]
  wire [15:0] trans_13_io_pipe_phv_out_header_13; // @[ipsa.scala 79:25]
  wire [15:0] trans_13_io_pipe_phv_out_header_14; // @[ipsa.scala 79:25]
  wire [15:0] trans_13_io_pipe_phv_out_header_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 79:25]
  wire [7:0] trans_13_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 79:25]
  wire [15:0] trans_13_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 79:25]
  wire [3:0] trans_13_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 79:25]
  wire  trans_13_io_pipe_phv_out_next_config_id; // @[ipsa.scala 79:25]
  wire  trans_13_io_pipe_phv_out_is_valid_processor; // @[ipsa.scala 79:25]
  wire  trans_13_io_pipe_phv_out_valid; // @[ipsa.scala 79:25]
  wire  trans_13_io_pipe_phv_out_last; // @[ipsa.scala 79:25]
  wire  trans_13_io_next_proc_exist; // @[ipsa.scala 79:25]
  wire  trans_14_clock; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_0; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_1; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_2; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_3; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_4; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_5; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_6; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_7; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_8; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_9; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_10; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_11; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_12; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_13; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_14; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_16; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_17; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_18; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_19; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_20; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_21; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_22; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_23; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_24; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_25; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_26; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_27; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_28; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_29; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_30; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_31; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_32; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_33; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_34; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_35; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_36; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_37; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_38; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_39; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_40; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_41; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_42; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_43; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_44; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_45; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_46; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_47; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_48; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_49; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_50; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_51; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_52; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_53; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_54; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_55; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_56; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_57; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_58; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_59; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_60; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_61; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_62; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_63; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_64; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_65; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_66; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_67; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_68; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_69; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_70; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_71; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_72; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_73; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_74; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_75; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_76; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_77; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_78; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_79; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_80; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_81; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_82; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_83; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_84; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_85; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_86; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_87; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_88; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_89; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_90; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_91; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_92; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_93; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_94; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_95; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_96; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_97; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_98; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_99; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_100; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_101; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_102; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_103; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_104; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_105; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_106; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_107; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_108; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_109; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_110; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_111; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_112; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_113; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_114; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_115; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_116; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_117; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_118; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_119; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_120; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_121; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_122; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_123; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_124; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_125; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_126; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_127; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_128; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_129; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_130; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_131; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_132; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_133; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_134; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_135; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_136; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_137; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_138; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_139; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_140; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_141; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_142; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_143; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_144; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_145; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_146; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_147; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_148; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_149; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_150; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_151; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_152; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_153; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_154; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_155; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_156; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_157; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_158; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_data_159; // @[ipsa.scala 79:25]
  wire [15:0] trans_14_io_pipe_phv_in_header_0; // @[ipsa.scala 79:25]
  wire [15:0] trans_14_io_pipe_phv_in_header_1; // @[ipsa.scala 79:25]
  wire [15:0] trans_14_io_pipe_phv_in_header_2; // @[ipsa.scala 79:25]
  wire [15:0] trans_14_io_pipe_phv_in_header_3; // @[ipsa.scala 79:25]
  wire [15:0] trans_14_io_pipe_phv_in_header_4; // @[ipsa.scala 79:25]
  wire [15:0] trans_14_io_pipe_phv_in_header_5; // @[ipsa.scala 79:25]
  wire [15:0] trans_14_io_pipe_phv_in_header_6; // @[ipsa.scala 79:25]
  wire [15:0] trans_14_io_pipe_phv_in_header_7; // @[ipsa.scala 79:25]
  wire [15:0] trans_14_io_pipe_phv_in_header_8; // @[ipsa.scala 79:25]
  wire [15:0] trans_14_io_pipe_phv_in_header_9; // @[ipsa.scala 79:25]
  wire [15:0] trans_14_io_pipe_phv_in_header_10; // @[ipsa.scala 79:25]
  wire [15:0] trans_14_io_pipe_phv_in_header_11; // @[ipsa.scala 79:25]
  wire [15:0] trans_14_io_pipe_phv_in_header_12; // @[ipsa.scala 79:25]
  wire [15:0] trans_14_io_pipe_phv_in_header_13; // @[ipsa.scala 79:25]
  wire [15:0] trans_14_io_pipe_phv_in_header_14; // @[ipsa.scala 79:25]
  wire [15:0] trans_14_io_pipe_phv_in_header_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_parse_current_state; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_in_parse_current_offset; // @[ipsa.scala 79:25]
  wire [15:0] trans_14_io_pipe_phv_in_parse_transition_field; // @[ipsa.scala 79:25]
  wire [3:0] trans_14_io_pipe_phv_in_next_processor_id; // @[ipsa.scala 79:25]
  wire  trans_14_io_pipe_phv_in_next_config_id; // @[ipsa.scala 79:25]
  wire  trans_14_io_pipe_phv_in_valid; // @[ipsa.scala 79:25]
  wire  trans_14_io_pipe_phv_in_last; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_0; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_1; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_2; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_3; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_4; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_5; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_6; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_7; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_8; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_9; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_10; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_11; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_12; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_13; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_14; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_16; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_17; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_18; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_19; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_20; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_21; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_22; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_23; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_24; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_25; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_26; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_27; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_28; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_29; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_30; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_31; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_32; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_33; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_34; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_35; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_36; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_37; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_38; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_39; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_40; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_41; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_42; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_43; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_44; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_45; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_46; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_47; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_48; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_49; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_50; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_51; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_52; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_53; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_54; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_55; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_56; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_57; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_58; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_59; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_60; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_61; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_62; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_63; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_64; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_65; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_66; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_67; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_68; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_69; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_70; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_71; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_72; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_73; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_74; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_75; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_76; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_77; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_78; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_79; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_80; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_81; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_82; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_83; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_84; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_85; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_86; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_87; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_88; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_89; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_90; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_91; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_92; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_93; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_94; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_95; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_96; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_97; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_98; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_99; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_100; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_101; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_102; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_103; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_104; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_105; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_106; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_107; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_108; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_109; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_110; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_111; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_112; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_113; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_114; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_115; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_116; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_117; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_118; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_119; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_120; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_121; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_122; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_123; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_124; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_125; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_126; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_127; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_128; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_129; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_130; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_131; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_132; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_133; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_134; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_135; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_136; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_137; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_138; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_139; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_140; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_141; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_142; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_143; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_144; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_145; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_146; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_147; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_148; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_149; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_150; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_151; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_152; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_153; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_154; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_155; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_156; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_157; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_158; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_data_159; // @[ipsa.scala 79:25]
  wire [15:0] trans_14_io_pipe_phv_out_header_0; // @[ipsa.scala 79:25]
  wire [15:0] trans_14_io_pipe_phv_out_header_1; // @[ipsa.scala 79:25]
  wire [15:0] trans_14_io_pipe_phv_out_header_2; // @[ipsa.scala 79:25]
  wire [15:0] trans_14_io_pipe_phv_out_header_3; // @[ipsa.scala 79:25]
  wire [15:0] trans_14_io_pipe_phv_out_header_4; // @[ipsa.scala 79:25]
  wire [15:0] trans_14_io_pipe_phv_out_header_5; // @[ipsa.scala 79:25]
  wire [15:0] trans_14_io_pipe_phv_out_header_6; // @[ipsa.scala 79:25]
  wire [15:0] trans_14_io_pipe_phv_out_header_7; // @[ipsa.scala 79:25]
  wire [15:0] trans_14_io_pipe_phv_out_header_8; // @[ipsa.scala 79:25]
  wire [15:0] trans_14_io_pipe_phv_out_header_9; // @[ipsa.scala 79:25]
  wire [15:0] trans_14_io_pipe_phv_out_header_10; // @[ipsa.scala 79:25]
  wire [15:0] trans_14_io_pipe_phv_out_header_11; // @[ipsa.scala 79:25]
  wire [15:0] trans_14_io_pipe_phv_out_header_12; // @[ipsa.scala 79:25]
  wire [15:0] trans_14_io_pipe_phv_out_header_13; // @[ipsa.scala 79:25]
  wire [15:0] trans_14_io_pipe_phv_out_header_14; // @[ipsa.scala 79:25]
  wire [15:0] trans_14_io_pipe_phv_out_header_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 79:25]
  wire [7:0] trans_14_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 79:25]
  wire [15:0] trans_14_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 79:25]
  wire [3:0] trans_14_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 79:25]
  wire  trans_14_io_pipe_phv_out_next_config_id; // @[ipsa.scala 79:25]
  wire  trans_14_io_pipe_phv_out_is_valid_processor; // @[ipsa.scala 79:25]
  wire  trans_14_io_pipe_phv_out_valid; // @[ipsa.scala 79:25]
  wire  trans_14_io_pipe_phv_out_last; // @[ipsa.scala 79:25]
  wire  trans_14_io_next_proc_exist; // @[ipsa.scala 79:25]
  wire  trans_15_clock; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_0; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_1; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_2; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_3; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_4; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_5; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_6; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_7; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_8; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_9; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_10; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_11; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_12; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_13; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_14; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_16; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_17; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_18; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_19; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_20; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_21; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_22; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_23; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_24; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_25; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_26; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_27; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_28; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_29; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_30; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_31; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_32; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_33; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_34; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_35; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_36; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_37; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_38; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_39; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_40; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_41; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_42; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_43; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_44; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_45; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_46; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_47; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_48; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_49; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_50; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_51; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_52; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_53; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_54; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_55; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_56; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_57; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_58; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_59; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_60; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_61; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_62; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_63; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_64; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_65; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_66; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_67; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_68; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_69; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_70; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_71; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_72; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_73; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_74; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_75; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_76; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_77; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_78; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_79; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_80; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_81; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_82; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_83; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_84; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_85; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_86; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_87; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_88; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_89; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_90; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_91; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_92; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_93; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_94; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_95; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_96; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_97; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_98; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_99; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_100; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_101; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_102; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_103; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_104; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_105; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_106; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_107; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_108; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_109; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_110; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_111; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_112; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_113; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_114; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_115; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_116; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_117; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_118; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_119; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_120; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_121; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_122; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_123; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_124; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_125; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_126; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_127; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_128; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_129; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_130; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_131; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_132; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_133; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_134; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_135; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_136; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_137; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_138; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_139; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_140; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_141; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_142; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_143; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_144; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_145; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_146; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_147; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_148; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_149; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_150; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_151; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_152; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_153; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_154; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_155; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_156; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_157; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_158; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_data_159; // @[ipsa.scala 79:25]
  wire [15:0] trans_15_io_pipe_phv_in_header_0; // @[ipsa.scala 79:25]
  wire [15:0] trans_15_io_pipe_phv_in_header_1; // @[ipsa.scala 79:25]
  wire [15:0] trans_15_io_pipe_phv_in_header_2; // @[ipsa.scala 79:25]
  wire [15:0] trans_15_io_pipe_phv_in_header_3; // @[ipsa.scala 79:25]
  wire [15:0] trans_15_io_pipe_phv_in_header_4; // @[ipsa.scala 79:25]
  wire [15:0] trans_15_io_pipe_phv_in_header_5; // @[ipsa.scala 79:25]
  wire [15:0] trans_15_io_pipe_phv_in_header_6; // @[ipsa.scala 79:25]
  wire [15:0] trans_15_io_pipe_phv_in_header_7; // @[ipsa.scala 79:25]
  wire [15:0] trans_15_io_pipe_phv_in_header_8; // @[ipsa.scala 79:25]
  wire [15:0] trans_15_io_pipe_phv_in_header_9; // @[ipsa.scala 79:25]
  wire [15:0] trans_15_io_pipe_phv_in_header_10; // @[ipsa.scala 79:25]
  wire [15:0] trans_15_io_pipe_phv_in_header_11; // @[ipsa.scala 79:25]
  wire [15:0] trans_15_io_pipe_phv_in_header_12; // @[ipsa.scala 79:25]
  wire [15:0] trans_15_io_pipe_phv_in_header_13; // @[ipsa.scala 79:25]
  wire [15:0] trans_15_io_pipe_phv_in_header_14; // @[ipsa.scala 79:25]
  wire [15:0] trans_15_io_pipe_phv_in_header_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_parse_current_state; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_in_parse_current_offset; // @[ipsa.scala 79:25]
  wire [15:0] trans_15_io_pipe_phv_in_parse_transition_field; // @[ipsa.scala 79:25]
  wire [3:0] trans_15_io_pipe_phv_in_next_processor_id; // @[ipsa.scala 79:25]
  wire  trans_15_io_pipe_phv_in_next_config_id; // @[ipsa.scala 79:25]
  wire  trans_15_io_pipe_phv_in_valid; // @[ipsa.scala 79:25]
  wire  trans_15_io_pipe_phv_in_last; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_0; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_1; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_2; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_3; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_4; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_5; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_6; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_7; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_8; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_9; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_10; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_11; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_12; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_13; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_14; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_16; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_17; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_18; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_19; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_20; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_21; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_22; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_23; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_24; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_25; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_26; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_27; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_28; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_29; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_30; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_31; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_32; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_33; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_34; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_35; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_36; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_37; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_38; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_39; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_40; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_41; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_42; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_43; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_44; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_45; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_46; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_47; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_48; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_49; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_50; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_51; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_52; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_53; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_54; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_55; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_56; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_57; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_58; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_59; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_60; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_61; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_62; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_63; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_64; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_65; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_66; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_67; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_68; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_69; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_70; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_71; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_72; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_73; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_74; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_75; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_76; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_77; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_78; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_79; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_80; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_81; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_82; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_83; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_84; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_85; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_86; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_87; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_88; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_89; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_90; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_91; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_92; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_93; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_94; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_95; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_96; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_97; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_98; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_99; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_100; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_101; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_102; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_103; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_104; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_105; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_106; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_107; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_108; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_109; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_110; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_111; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_112; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_113; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_114; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_115; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_116; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_117; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_118; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_119; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_120; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_121; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_122; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_123; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_124; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_125; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_126; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_127; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_128; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_129; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_130; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_131; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_132; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_133; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_134; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_135; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_136; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_137; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_138; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_139; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_140; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_141; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_142; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_143; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_144; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_145; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_146; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_147; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_148; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_149; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_150; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_151; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_152; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_153; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_154; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_155; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_156; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_157; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_158; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_data_159; // @[ipsa.scala 79:25]
  wire [15:0] trans_15_io_pipe_phv_out_header_0; // @[ipsa.scala 79:25]
  wire [15:0] trans_15_io_pipe_phv_out_header_1; // @[ipsa.scala 79:25]
  wire [15:0] trans_15_io_pipe_phv_out_header_2; // @[ipsa.scala 79:25]
  wire [15:0] trans_15_io_pipe_phv_out_header_3; // @[ipsa.scala 79:25]
  wire [15:0] trans_15_io_pipe_phv_out_header_4; // @[ipsa.scala 79:25]
  wire [15:0] trans_15_io_pipe_phv_out_header_5; // @[ipsa.scala 79:25]
  wire [15:0] trans_15_io_pipe_phv_out_header_6; // @[ipsa.scala 79:25]
  wire [15:0] trans_15_io_pipe_phv_out_header_7; // @[ipsa.scala 79:25]
  wire [15:0] trans_15_io_pipe_phv_out_header_8; // @[ipsa.scala 79:25]
  wire [15:0] trans_15_io_pipe_phv_out_header_9; // @[ipsa.scala 79:25]
  wire [15:0] trans_15_io_pipe_phv_out_header_10; // @[ipsa.scala 79:25]
  wire [15:0] trans_15_io_pipe_phv_out_header_11; // @[ipsa.scala 79:25]
  wire [15:0] trans_15_io_pipe_phv_out_header_12; // @[ipsa.scala 79:25]
  wire [15:0] trans_15_io_pipe_phv_out_header_13; // @[ipsa.scala 79:25]
  wire [15:0] trans_15_io_pipe_phv_out_header_14; // @[ipsa.scala 79:25]
  wire [15:0] trans_15_io_pipe_phv_out_header_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 79:25]
  wire [7:0] trans_15_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 79:25]
  wire [15:0] trans_15_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 79:25]
  wire [3:0] trans_15_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 79:25]
  wire  trans_15_io_pipe_phv_out_next_config_id; // @[ipsa.scala 79:25]
  wire  trans_15_io_pipe_phv_out_is_valid_processor; // @[ipsa.scala 79:25]
  wire  trans_15_io_pipe_phv_out_valid; // @[ipsa.scala 79:25]
  wire  trans_15_io_pipe_phv_out_last; // @[ipsa.scala 79:25]
  wire  trans_15_io_next_proc_exist; // @[ipsa.scala 79:25]
  Processor proc_0 ( // @[ipsa.scala 56:25]
    .clock(proc_0_clock),
    .io_pipe_phv_in_data_0(proc_0_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(proc_0_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(proc_0_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(proc_0_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(proc_0_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(proc_0_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(proc_0_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(proc_0_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(proc_0_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(proc_0_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(proc_0_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(proc_0_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(proc_0_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(proc_0_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(proc_0_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(proc_0_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(proc_0_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(proc_0_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(proc_0_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(proc_0_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(proc_0_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(proc_0_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(proc_0_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(proc_0_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(proc_0_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(proc_0_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(proc_0_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(proc_0_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(proc_0_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(proc_0_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(proc_0_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(proc_0_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(proc_0_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(proc_0_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(proc_0_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(proc_0_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(proc_0_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(proc_0_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(proc_0_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(proc_0_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(proc_0_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(proc_0_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(proc_0_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(proc_0_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(proc_0_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(proc_0_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(proc_0_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(proc_0_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(proc_0_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(proc_0_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(proc_0_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(proc_0_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(proc_0_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(proc_0_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(proc_0_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(proc_0_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(proc_0_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(proc_0_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(proc_0_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(proc_0_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(proc_0_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(proc_0_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(proc_0_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(proc_0_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(proc_0_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(proc_0_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(proc_0_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(proc_0_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(proc_0_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(proc_0_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(proc_0_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(proc_0_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(proc_0_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(proc_0_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(proc_0_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(proc_0_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(proc_0_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(proc_0_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(proc_0_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(proc_0_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(proc_0_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(proc_0_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(proc_0_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(proc_0_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(proc_0_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(proc_0_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(proc_0_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(proc_0_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(proc_0_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(proc_0_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(proc_0_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(proc_0_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(proc_0_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(proc_0_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(proc_0_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(proc_0_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(proc_0_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(proc_0_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(proc_0_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(proc_0_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(proc_0_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(proc_0_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(proc_0_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(proc_0_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(proc_0_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(proc_0_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(proc_0_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(proc_0_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(proc_0_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(proc_0_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(proc_0_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(proc_0_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(proc_0_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(proc_0_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(proc_0_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(proc_0_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(proc_0_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(proc_0_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(proc_0_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(proc_0_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(proc_0_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(proc_0_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(proc_0_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(proc_0_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(proc_0_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(proc_0_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(proc_0_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(proc_0_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(proc_0_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(proc_0_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(proc_0_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(proc_0_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(proc_0_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(proc_0_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(proc_0_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(proc_0_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(proc_0_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(proc_0_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(proc_0_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(proc_0_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(proc_0_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(proc_0_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(proc_0_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(proc_0_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(proc_0_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(proc_0_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(proc_0_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(proc_0_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(proc_0_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(proc_0_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(proc_0_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(proc_0_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(proc_0_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(proc_0_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(proc_0_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(proc_0_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(proc_0_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(proc_0_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(proc_0_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(proc_0_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_header_0(proc_0_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(proc_0_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(proc_0_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(proc_0_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(proc_0_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(proc_0_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(proc_0_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(proc_0_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(proc_0_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(proc_0_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(proc_0_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(proc_0_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(proc_0_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(proc_0_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(proc_0_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(proc_0_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(proc_0_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(proc_0_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(proc_0_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(proc_0_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(proc_0_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(proc_0_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_in_valid(proc_0_io_pipe_phv_in_valid),
    .io_pipe_phv_in_last(proc_0_io_pipe_phv_in_last),
    .io_pipe_phv_out_data_0(proc_0_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(proc_0_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(proc_0_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(proc_0_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(proc_0_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(proc_0_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(proc_0_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(proc_0_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(proc_0_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(proc_0_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(proc_0_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(proc_0_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(proc_0_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(proc_0_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(proc_0_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(proc_0_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(proc_0_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(proc_0_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(proc_0_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(proc_0_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(proc_0_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(proc_0_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(proc_0_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(proc_0_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(proc_0_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(proc_0_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(proc_0_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(proc_0_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(proc_0_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(proc_0_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(proc_0_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(proc_0_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(proc_0_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(proc_0_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(proc_0_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(proc_0_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(proc_0_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(proc_0_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(proc_0_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(proc_0_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(proc_0_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(proc_0_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(proc_0_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(proc_0_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(proc_0_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(proc_0_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(proc_0_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(proc_0_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(proc_0_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(proc_0_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(proc_0_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(proc_0_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(proc_0_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(proc_0_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(proc_0_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(proc_0_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(proc_0_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(proc_0_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(proc_0_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(proc_0_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(proc_0_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(proc_0_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(proc_0_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(proc_0_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(proc_0_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(proc_0_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(proc_0_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(proc_0_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(proc_0_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(proc_0_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(proc_0_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(proc_0_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(proc_0_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(proc_0_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(proc_0_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(proc_0_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(proc_0_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(proc_0_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(proc_0_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(proc_0_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(proc_0_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(proc_0_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(proc_0_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(proc_0_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(proc_0_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(proc_0_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(proc_0_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(proc_0_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(proc_0_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(proc_0_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(proc_0_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(proc_0_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(proc_0_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(proc_0_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(proc_0_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(proc_0_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(proc_0_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(proc_0_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(proc_0_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(proc_0_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(proc_0_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(proc_0_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(proc_0_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(proc_0_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(proc_0_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(proc_0_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(proc_0_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(proc_0_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(proc_0_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(proc_0_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(proc_0_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(proc_0_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(proc_0_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(proc_0_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(proc_0_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(proc_0_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(proc_0_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(proc_0_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(proc_0_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(proc_0_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(proc_0_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(proc_0_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(proc_0_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(proc_0_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(proc_0_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(proc_0_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(proc_0_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(proc_0_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(proc_0_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(proc_0_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(proc_0_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(proc_0_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(proc_0_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(proc_0_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(proc_0_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(proc_0_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(proc_0_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(proc_0_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(proc_0_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(proc_0_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(proc_0_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(proc_0_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(proc_0_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(proc_0_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(proc_0_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(proc_0_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(proc_0_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(proc_0_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(proc_0_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(proc_0_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(proc_0_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(proc_0_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(proc_0_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(proc_0_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(proc_0_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(proc_0_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(proc_0_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(proc_0_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(proc_0_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(proc_0_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_header_0(proc_0_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(proc_0_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(proc_0_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(proc_0_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(proc_0_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(proc_0_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(proc_0_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(proc_0_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(proc_0_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(proc_0_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(proc_0_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(proc_0_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(proc_0_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(proc_0_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(proc_0_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(proc_0_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(proc_0_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(proc_0_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(proc_0_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(proc_0_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(proc_0_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_valid(proc_0_io_pipe_phv_out_valid),
    .io_pipe_phv_out_last(proc_0_io_pipe_phv_out_last)
  );
  Processor proc_1 ( // @[ipsa.scala 56:25]
    .clock(proc_1_clock),
    .io_pipe_phv_in_data_0(proc_1_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(proc_1_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(proc_1_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(proc_1_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(proc_1_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(proc_1_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(proc_1_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(proc_1_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(proc_1_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(proc_1_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(proc_1_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(proc_1_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(proc_1_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(proc_1_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(proc_1_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(proc_1_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(proc_1_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(proc_1_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(proc_1_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(proc_1_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(proc_1_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(proc_1_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(proc_1_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(proc_1_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(proc_1_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(proc_1_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(proc_1_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(proc_1_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(proc_1_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(proc_1_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(proc_1_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(proc_1_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(proc_1_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(proc_1_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(proc_1_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(proc_1_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(proc_1_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(proc_1_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(proc_1_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(proc_1_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(proc_1_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(proc_1_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(proc_1_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(proc_1_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(proc_1_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(proc_1_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(proc_1_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(proc_1_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(proc_1_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(proc_1_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(proc_1_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(proc_1_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(proc_1_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(proc_1_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(proc_1_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(proc_1_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(proc_1_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(proc_1_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(proc_1_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(proc_1_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(proc_1_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(proc_1_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(proc_1_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(proc_1_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(proc_1_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(proc_1_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(proc_1_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(proc_1_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(proc_1_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(proc_1_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(proc_1_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(proc_1_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(proc_1_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(proc_1_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(proc_1_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(proc_1_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(proc_1_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(proc_1_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(proc_1_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(proc_1_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(proc_1_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(proc_1_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(proc_1_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(proc_1_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(proc_1_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(proc_1_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(proc_1_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(proc_1_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(proc_1_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(proc_1_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(proc_1_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(proc_1_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(proc_1_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(proc_1_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(proc_1_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(proc_1_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(proc_1_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(proc_1_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(proc_1_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(proc_1_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(proc_1_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(proc_1_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(proc_1_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(proc_1_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(proc_1_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(proc_1_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(proc_1_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(proc_1_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(proc_1_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(proc_1_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(proc_1_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(proc_1_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(proc_1_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(proc_1_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(proc_1_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(proc_1_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(proc_1_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(proc_1_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(proc_1_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(proc_1_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(proc_1_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(proc_1_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(proc_1_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(proc_1_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(proc_1_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(proc_1_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(proc_1_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(proc_1_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(proc_1_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(proc_1_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(proc_1_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(proc_1_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(proc_1_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(proc_1_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(proc_1_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(proc_1_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(proc_1_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(proc_1_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(proc_1_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(proc_1_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(proc_1_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(proc_1_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(proc_1_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(proc_1_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(proc_1_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(proc_1_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(proc_1_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(proc_1_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(proc_1_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(proc_1_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(proc_1_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(proc_1_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(proc_1_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(proc_1_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(proc_1_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(proc_1_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(proc_1_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(proc_1_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(proc_1_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(proc_1_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_header_0(proc_1_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(proc_1_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(proc_1_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(proc_1_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(proc_1_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(proc_1_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(proc_1_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(proc_1_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(proc_1_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(proc_1_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(proc_1_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(proc_1_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(proc_1_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(proc_1_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(proc_1_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(proc_1_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(proc_1_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(proc_1_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(proc_1_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(proc_1_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(proc_1_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(proc_1_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_in_valid(proc_1_io_pipe_phv_in_valid),
    .io_pipe_phv_in_last(proc_1_io_pipe_phv_in_last),
    .io_pipe_phv_out_data_0(proc_1_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(proc_1_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(proc_1_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(proc_1_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(proc_1_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(proc_1_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(proc_1_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(proc_1_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(proc_1_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(proc_1_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(proc_1_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(proc_1_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(proc_1_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(proc_1_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(proc_1_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(proc_1_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(proc_1_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(proc_1_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(proc_1_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(proc_1_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(proc_1_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(proc_1_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(proc_1_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(proc_1_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(proc_1_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(proc_1_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(proc_1_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(proc_1_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(proc_1_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(proc_1_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(proc_1_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(proc_1_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(proc_1_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(proc_1_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(proc_1_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(proc_1_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(proc_1_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(proc_1_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(proc_1_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(proc_1_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(proc_1_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(proc_1_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(proc_1_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(proc_1_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(proc_1_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(proc_1_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(proc_1_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(proc_1_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(proc_1_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(proc_1_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(proc_1_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(proc_1_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(proc_1_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(proc_1_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(proc_1_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(proc_1_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(proc_1_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(proc_1_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(proc_1_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(proc_1_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(proc_1_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(proc_1_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(proc_1_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(proc_1_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(proc_1_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(proc_1_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(proc_1_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(proc_1_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(proc_1_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(proc_1_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(proc_1_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(proc_1_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(proc_1_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(proc_1_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(proc_1_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(proc_1_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(proc_1_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(proc_1_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(proc_1_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(proc_1_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(proc_1_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(proc_1_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(proc_1_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(proc_1_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(proc_1_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(proc_1_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(proc_1_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(proc_1_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(proc_1_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(proc_1_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(proc_1_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(proc_1_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(proc_1_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(proc_1_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(proc_1_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(proc_1_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(proc_1_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(proc_1_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(proc_1_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(proc_1_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(proc_1_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(proc_1_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(proc_1_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(proc_1_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(proc_1_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(proc_1_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(proc_1_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(proc_1_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(proc_1_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(proc_1_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(proc_1_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(proc_1_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(proc_1_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(proc_1_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(proc_1_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(proc_1_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(proc_1_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(proc_1_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(proc_1_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(proc_1_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(proc_1_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(proc_1_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(proc_1_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(proc_1_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(proc_1_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(proc_1_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(proc_1_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(proc_1_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(proc_1_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(proc_1_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(proc_1_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(proc_1_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(proc_1_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(proc_1_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(proc_1_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(proc_1_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(proc_1_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(proc_1_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(proc_1_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(proc_1_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(proc_1_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(proc_1_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(proc_1_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(proc_1_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(proc_1_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(proc_1_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(proc_1_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(proc_1_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(proc_1_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(proc_1_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(proc_1_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(proc_1_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(proc_1_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(proc_1_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(proc_1_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(proc_1_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(proc_1_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(proc_1_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(proc_1_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(proc_1_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_header_0(proc_1_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(proc_1_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(proc_1_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(proc_1_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(proc_1_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(proc_1_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(proc_1_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(proc_1_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(proc_1_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(proc_1_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(proc_1_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(proc_1_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(proc_1_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(proc_1_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(proc_1_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(proc_1_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(proc_1_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(proc_1_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(proc_1_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(proc_1_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(proc_1_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_valid(proc_1_io_pipe_phv_out_valid),
    .io_pipe_phv_out_last(proc_1_io_pipe_phv_out_last)
  );
  Processor proc_2 ( // @[ipsa.scala 56:25]
    .clock(proc_2_clock),
    .io_pipe_phv_in_data_0(proc_2_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(proc_2_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(proc_2_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(proc_2_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(proc_2_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(proc_2_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(proc_2_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(proc_2_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(proc_2_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(proc_2_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(proc_2_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(proc_2_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(proc_2_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(proc_2_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(proc_2_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(proc_2_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(proc_2_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(proc_2_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(proc_2_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(proc_2_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(proc_2_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(proc_2_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(proc_2_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(proc_2_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(proc_2_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(proc_2_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(proc_2_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(proc_2_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(proc_2_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(proc_2_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(proc_2_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(proc_2_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(proc_2_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(proc_2_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(proc_2_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(proc_2_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(proc_2_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(proc_2_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(proc_2_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(proc_2_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(proc_2_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(proc_2_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(proc_2_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(proc_2_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(proc_2_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(proc_2_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(proc_2_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(proc_2_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(proc_2_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(proc_2_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(proc_2_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(proc_2_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(proc_2_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(proc_2_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(proc_2_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(proc_2_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(proc_2_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(proc_2_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(proc_2_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(proc_2_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(proc_2_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(proc_2_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(proc_2_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(proc_2_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(proc_2_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(proc_2_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(proc_2_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(proc_2_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(proc_2_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(proc_2_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(proc_2_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(proc_2_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(proc_2_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(proc_2_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(proc_2_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(proc_2_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(proc_2_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(proc_2_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(proc_2_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(proc_2_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(proc_2_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(proc_2_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(proc_2_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(proc_2_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(proc_2_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(proc_2_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(proc_2_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(proc_2_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(proc_2_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(proc_2_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(proc_2_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(proc_2_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(proc_2_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(proc_2_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(proc_2_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(proc_2_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(proc_2_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(proc_2_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(proc_2_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(proc_2_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(proc_2_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(proc_2_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(proc_2_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(proc_2_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(proc_2_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(proc_2_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(proc_2_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(proc_2_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(proc_2_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(proc_2_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(proc_2_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(proc_2_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(proc_2_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(proc_2_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(proc_2_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(proc_2_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(proc_2_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(proc_2_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(proc_2_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(proc_2_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(proc_2_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(proc_2_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(proc_2_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(proc_2_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(proc_2_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(proc_2_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(proc_2_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(proc_2_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(proc_2_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(proc_2_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(proc_2_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(proc_2_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(proc_2_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(proc_2_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(proc_2_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(proc_2_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(proc_2_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(proc_2_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(proc_2_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(proc_2_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(proc_2_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(proc_2_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(proc_2_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(proc_2_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(proc_2_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(proc_2_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(proc_2_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(proc_2_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(proc_2_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(proc_2_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(proc_2_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(proc_2_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(proc_2_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(proc_2_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(proc_2_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(proc_2_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(proc_2_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(proc_2_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(proc_2_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(proc_2_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_header_0(proc_2_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(proc_2_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(proc_2_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(proc_2_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(proc_2_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(proc_2_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(proc_2_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(proc_2_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(proc_2_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(proc_2_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(proc_2_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(proc_2_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(proc_2_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(proc_2_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(proc_2_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(proc_2_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(proc_2_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(proc_2_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(proc_2_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(proc_2_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(proc_2_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(proc_2_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_in_valid(proc_2_io_pipe_phv_in_valid),
    .io_pipe_phv_in_last(proc_2_io_pipe_phv_in_last),
    .io_pipe_phv_out_data_0(proc_2_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(proc_2_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(proc_2_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(proc_2_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(proc_2_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(proc_2_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(proc_2_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(proc_2_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(proc_2_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(proc_2_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(proc_2_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(proc_2_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(proc_2_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(proc_2_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(proc_2_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(proc_2_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(proc_2_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(proc_2_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(proc_2_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(proc_2_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(proc_2_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(proc_2_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(proc_2_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(proc_2_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(proc_2_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(proc_2_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(proc_2_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(proc_2_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(proc_2_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(proc_2_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(proc_2_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(proc_2_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(proc_2_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(proc_2_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(proc_2_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(proc_2_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(proc_2_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(proc_2_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(proc_2_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(proc_2_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(proc_2_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(proc_2_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(proc_2_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(proc_2_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(proc_2_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(proc_2_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(proc_2_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(proc_2_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(proc_2_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(proc_2_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(proc_2_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(proc_2_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(proc_2_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(proc_2_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(proc_2_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(proc_2_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(proc_2_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(proc_2_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(proc_2_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(proc_2_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(proc_2_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(proc_2_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(proc_2_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(proc_2_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(proc_2_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(proc_2_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(proc_2_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(proc_2_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(proc_2_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(proc_2_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(proc_2_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(proc_2_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(proc_2_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(proc_2_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(proc_2_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(proc_2_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(proc_2_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(proc_2_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(proc_2_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(proc_2_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(proc_2_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(proc_2_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(proc_2_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(proc_2_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(proc_2_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(proc_2_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(proc_2_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(proc_2_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(proc_2_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(proc_2_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(proc_2_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(proc_2_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(proc_2_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(proc_2_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(proc_2_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(proc_2_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(proc_2_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(proc_2_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(proc_2_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(proc_2_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(proc_2_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(proc_2_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(proc_2_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(proc_2_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(proc_2_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(proc_2_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(proc_2_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(proc_2_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(proc_2_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(proc_2_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(proc_2_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(proc_2_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(proc_2_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(proc_2_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(proc_2_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(proc_2_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(proc_2_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(proc_2_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(proc_2_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(proc_2_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(proc_2_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(proc_2_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(proc_2_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(proc_2_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(proc_2_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(proc_2_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(proc_2_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(proc_2_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(proc_2_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(proc_2_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(proc_2_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(proc_2_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(proc_2_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(proc_2_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(proc_2_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(proc_2_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(proc_2_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(proc_2_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(proc_2_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(proc_2_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(proc_2_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(proc_2_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(proc_2_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(proc_2_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(proc_2_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(proc_2_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(proc_2_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(proc_2_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(proc_2_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(proc_2_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(proc_2_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(proc_2_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(proc_2_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(proc_2_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(proc_2_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(proc_2_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(proc_2_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(proc_2_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(proc_2_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(proc_2_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_header_0(proc_2_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(proc_2_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(proc_2_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(proc_2_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(proc_2_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(proc_2_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(proc_2_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(proc_2_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(proc_2_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(proc_2_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(proc_2_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(proc_2_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(proc_2_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(proc_2_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(proc_2_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(proc_2_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(proc_2_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(proc_2_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(proc_2_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(proc_2_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(proc_2_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_valid(proc_2_io_pipe_phv_out_valid),
    .io_pipe_phv_out_last(proc_2_io_pipe_phv_out_last)
  );
  Processor proc_3 ( // @[ipsa.scala 56:25]
    .clock(proc_3_clock),
    .io_pipe_phv_in_data_0(proc_3_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(proc_3_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(proc_3_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(proc_3_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(proc_3_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(proc_3_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(proc_3_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(proc_3_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(proc_3_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(proc_3_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(proc_3_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(proc_3_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(proc_3_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(proc_3_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(proc_3_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(proc_3_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(proc_3_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(proc_3_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(proc_3_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(proc_3_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(proc_3_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(proc_3_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(proc_3_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(proc_3_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(proc_3_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(proc_3_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(proc_3_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(proc_3_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(proc_3_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(proc_3_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(proc_3_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(proc_3_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(proc_3_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(proc_3_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(proc_3_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(proc_3_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(proc_3_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(proc_3_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(proc_3_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(proc_3_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(proc_3_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(proc_3_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(proc_3_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(proc_3_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(proc_3_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(proc_3_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(proc_3_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(proc_3_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(proc_3_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(proc_3_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(proc_3_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(proc_3_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(proc_3_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(proc_3_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(proc_3_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(proc_3_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(proc_3_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(proc_3_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(proc_3_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(proc_3_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(proc_3_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(proc_3_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(proc_3_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(proc_3_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(proc_3_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(proc_3_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(proc_3_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(proc_3_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(proc_3_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(proc_3_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(proc_3_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(proc_3_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(proc_3_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(proc_3_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(proc_3_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(proc_3_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(proc_3_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(proc_3_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(proc_3_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(proc_3_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(proc_3_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(proc_3_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(proc_3_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(proc_3_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(proc_3_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(proc_3_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(proc_3_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(proc_3_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(proc_3_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(proc_3_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(proc_3_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(proc_3_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(proc_3_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(proc_3_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(proc_3_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(proc_3_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(proc_3_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(proc_3_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(proc_3_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(proc_3_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(proc_3_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(proc_3_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(proc_3_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(proc_3_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(proc_3_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(proc_3_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(proc_3_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(proc_3_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(proc_3_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(proc_3_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(proc_3_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(proc_3_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(proc_3_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(proc_3_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(proc_3_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(proc_3_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(proc_3_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(proc_3_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(proc_3_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(proc_3_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(proc_3_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(proc_3_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(proc_3_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(proc_3_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(proc_3_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(proc_3_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(proc_3_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(proc_3_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(proc_3_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(proc_3_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(proc_3_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(proc_3_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(proc_3_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(proc_3_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(proc_3_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(proc_3_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(proc_3_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(proc_3_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(proc_3_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(proc_3_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(proc_3_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(proc_3_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(proc_3_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(proc_3_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(proc_3_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(proc_3_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(proc_3_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(proc_3_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(proc_3_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(proc_3_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(proc_3_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(proc_3_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(proc_3_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(proc_3_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(proc_3_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(proc_3_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(proc_3_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(proc_3_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(proc_3_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(proc_3_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_header_0(proc_3_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(proc_3_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(proc_3_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(proc_3_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(proc_3_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(proc_3_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(proc_3_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(proc_3_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(proc_3_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(proc_3_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(proc_3_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(proc_3_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(proc_3_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(proc_3_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(proc_3_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(proc_3_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(proc_3_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(proc_3_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(proc_3_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(proc_3_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(proc_3_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(proc_3_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_in_valid(proc_3_io_pipe_phv_in_valid),
    .io_pipe_phv_in_last(proc_3_io_pipe_phv_in_last),
    .io_pipe_phv_out_data_0(proc_3_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(proc_3_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(proc_3_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(proc_3_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(proc_3_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(proc_3_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(proc_3_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(proc_3_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(proc_3_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(proc_3_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(proc_3_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(proc_3_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(proc_3_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(proc_3_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(proc_3_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(proc_3_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(proc_3_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(proc_3_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(proc_3_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(proc_3_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(proc_3_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(proc_3_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(proc_3_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(proc_3_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(proc_3_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(proc_3_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(proc_3_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(proc_3_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(proc_3_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(proc_3_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(proc_3_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(proc_3_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(proc_3_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(proc_3_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(proc_3_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(proc_3_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(proc_3_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(proc_3_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(proc_3_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(proc_3_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(proc_3_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(proc_3_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(proc_3_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(proc_3_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(proc_3_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(proc_3_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(proc_3_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(proc_3_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(proc_3_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(proc_3_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(proc_3_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(proc_3_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(proc_3_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(proc_3_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(proc_3_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(proc_3_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(proc_3_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(proc_3_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(proc_3_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(proc_3_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(proc_3_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(proc_3_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(proc_3_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(proc_3_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(proc_3_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(proc_3_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(proc_3_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(proc_3_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(proc_3_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(proc_3_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(proc_3_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(proc_3_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(proc_3_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(proc_3_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(proc_3_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(proc_3_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(proc_3_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(proc_3_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(proc_3_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(proc_3_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(proc_3_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(proc_3_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(proc_3_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(proc_3_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(proc_3_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(proc_3_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(proc_3_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(proc_3_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(proc_3_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(proc_3_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(proc_3_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(proc_3_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(proc_3_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(proc_3_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(proc_3_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(proc_3_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(proc_3_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(proc_3_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(proc_3_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(proc_3_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(proc_3_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(proc_3_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(proc_3_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(proc_3_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(proc_3_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(proc_3_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(proc_3_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(proc_3_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(proc_3_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(proc_3_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(proc_3_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(proc_3_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(proc_3_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(proc_3_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(proc_3_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(proc_3_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(proc_3_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(proc_3_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(proc_3_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(proc_3_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(proc_3_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(proc_3_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(proc_3_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(proc_3_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(proc_3_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(proc_3_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(proc_3_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(proc_3_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(proc_3_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(proc_3_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(proc_3_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(proc_3_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(proc_3_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(proc_3_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(proc_3_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(proc_3_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(proc_3_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(proc_3_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(proc_3_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(proc_3_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(proc_3_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(proc_3_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(proc_3_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(proc_3_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(proc_3_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(proc_3_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(proc_3_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(proc_3_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(proc_3_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(proc_3_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(proc_3_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(proc_3_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(proc_3_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(proc_3_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(proc_3_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(proc_3_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(proc_3_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(proc_3_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(proc_3_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(proc_3_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_header_0(proc_3_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(proc_3_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(proc_3_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(proc_3_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(proc_3_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(proc_3_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(proc_3_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(proc_3_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(proc_3_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(proc_3_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(proc_3_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(proc_3_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(proc_3_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(proc_3_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(proc_3_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(proc_3_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(proc_3_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(proc_3_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(proc_3_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(proc_3_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(proc_3_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_valid(proc_3_io_pipe_phv_out_valid),
    .io_pipe_phv_out_last(proc_3_io_pipe_phv_out_last)
  );
  Processor proc_4 ( // @[ipsa.scala 56:25]
    .clock(proc_4_clock),
    .io_pipe_phv_in_data_0(proc_4_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(proc_4_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(proc_4_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(proc_4_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(proc_4_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(proc_4_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(proc_4_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(proc_4_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(proc_4_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(proc_4_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(proc_4_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(proc_4_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(proc_4_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(proc_4_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(proc_4_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(proc_4_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(proc_4_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(proc_4_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(proc_4_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(proc_4_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(proc_4_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(proc_4_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(proc_4_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(proc_4_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(proc_4_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(proc_4_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(proc_4_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(proc_4_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(proc_4_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(proc_4_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(proc_4_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(proc_4_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(proc_4_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(proc_4_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(proc_4_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(proc_4_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(proc_4_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(proc_4_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(proc_4_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(proc_4_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(proc_4_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(proc_4_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(proc_4_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(proc_4_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(proc_4_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(proc_4_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(proc_4_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(proc_4_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(proc_4_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(proc_4_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(proc_4_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(proc_4_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(proc_4_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(proc_4_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(proc_4_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(proc_4_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(proc_4_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(proc_4_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(proc_4_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(proc_4_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(proc_4_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(proc_4_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(proc_4_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(proc_4_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(proc_4_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(proc_4_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(proc_4_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(proc_4_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(proc_4_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(proc_4_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(proc_4_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(proc_4_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(proc_4_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(proc_4_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(proc_4_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(proc_4_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(proc_4_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(proc_4_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(proc_4_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(proc_4_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(proc_4_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(proc_4_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(proc_4_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(proc_4_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(proc_4_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(proc_4_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(proc_4_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(proc_4_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(proc_4_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(proc_4_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(proc_4_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(proc_4_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(proc_4_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(proc_4_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(proc_4_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(proc_4_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(proc_4_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(proc_4_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(proc_4_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(proc_4_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(proc_4_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(proc_4_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(proc_4_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(proc_4_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(proc_4_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(proc_4_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(proc_4_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(proc_4_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(proc_4_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(proc_4_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(proc_4_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(proc_4_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(proc_4_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(proc_4_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(proc_4_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(proc_4_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(proc_4_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(proc_4_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(proc_4_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(proc_4_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(proc_4_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(proc_4_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(proc_4_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(proc_4_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(proc_4_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(proc_4_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(proc_4_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(proc_4_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(proc_4_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(proc_4_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(proc_4_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(proc_4_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(proc_4_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(proc_4_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(proc_4_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(proc_4_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(proc_4_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(proc_4_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(proc_4_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(proc_4_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(proc_4_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(proc_4_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(proc_4_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(proc_4_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(proc_4_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(proc_4_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(proc_4_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(proc_4_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(proc_4_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(proc_4_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(proc_4_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(proc_4_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(proc_4_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(proc_4_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(proc_4_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(proc_4_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(proc_4_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(proc_4_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(proc_4_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(proc_4_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_header_0(proc_4_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(proc_4_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(proc_4_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(proc_4_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(proc_4_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(proc_4_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(proc_4_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(proc_4_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(proc_4_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(proc_4_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(proc_4_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(proc_4_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(proc_4_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(proc_4_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(proc_4_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(proc_4_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(proc_4_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(proc_4_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(proc_4_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(proc_4_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(proc_4_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(proc_4_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_in_valid(proc_4_io_pipe_phv_in_valid),
    .io_pipe_phv_in_last(proc_4_io_pipe_phv_in_last),
    .io_pipe_phv_out_data_0(proc_4_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(proc_4_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(proc_4_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(proc_4_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(proc_4_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(proc_4_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(proc_4_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(proc_4_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(proc_4_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(proc_4_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(proc_4_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(proc_4_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(proc_4_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(proc_4_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(proc_4_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(proc_4_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(proc_4_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(proc_4_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(proc_4_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(proc_4_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(proc_4_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(proc_4_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(proc_4_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(proc_4_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(proc_4_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(proc_4_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(proc_4_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(proc_4_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(proc_4_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(proc_4_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(proc_4_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(proc_4_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(proc_4_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(proc_4_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(proc_4_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(proc_4_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(proc_4_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(proc_4_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(proc_4_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(proc_4_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(proc_4_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(proc_4_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(proc_4_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(proc_4_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(proc_4_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(proc_4_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(proc_4_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(proc_4_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(proc_4_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(proc_4_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(proc_4_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(proc_4_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(proc_4_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(proc_4_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(proc_4_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(proc_4_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(proc_4_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(proc_4_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(proc_4_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(proc_4_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(proc_4_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(proc_4_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(proc_4_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(proc_4_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(proc_4_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(proc_4_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(proc_4_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(proc_4_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(proc_4_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(proc_4_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(proc_4_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(proc_4_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(proc_4_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(proc_4_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(proc_4_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(proc_4_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(proc_4_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(proc_4_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(proc_4_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(proc_4_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(proc_4_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(proc_4_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(proc_4_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(proc_4_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(proc_4_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(proc_4_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(proc_4_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(proc_4_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(proc_4_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(proc_4_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(proc_4_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(proc_4_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(proc_4_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(proc_4_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(proc_4_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(proc_4_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(proc_4_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(proc_4_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(proc_4_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(proc_4_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(proc_4_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(proc_4_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(proc_4_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(proc_4_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(proc_4_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(proc_4_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(proc_4_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(proc_4_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(proc_4_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(proc_4_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(proc_4_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(proc_4_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(proc_4_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(proc_4_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(proc_4_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(proc_4_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(proc_4_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(proc_4_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(proc_4_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(proc_4_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(proc_4_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(proc_4_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(proc_4_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(proc_4_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(proc_4_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(proc_4_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(proc_4_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(proc_4_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(proc_4_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(proc_4_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(proc_4_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(proc_4_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(proc_4_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(proc_4_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(proc_4_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(proc_4_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(proc_4_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(proc_4_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(proc_4_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(proc_4_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(proc_4_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(proc_4_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(proc_4_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(proc_4_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(proc_4_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(proc_4_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(proc_4_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(proc_4_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(proc_4_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(proc_4_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(proc_4_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(proc_4_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(proc_4_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(proc_4_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(proc_4_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(proc_4_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(proc_4_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(proc_4_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(proc_4_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(proc_4_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_header_0(proc_4_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(proc_4_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(proc_4_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(proc_4_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(proc_4_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(proc_4_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(proc_4_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(proc_4_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(proc_4_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(proc_4_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(proc_4_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(proc_4_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(proc_4_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(proc_4_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(proc_4_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(proc_4_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(proc_4_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(proc_4_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(proc_4_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(proc_4_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(proc_4_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_valid(proc_4_io_pipe_phv_out_valid),
    .io_pipe_phv_out_last(proc_4_io_pipe_phv_out_last)
  );
  Processor proc_5 ( // @[ipsa.scala 56:25]
    .clock(proc_5_clock),
    .io_pipe_phv_in_data_0(proc_5_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(proc_5_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(proc_5_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(proc_5_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(proc_5_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(proc_5_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(proc_5_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(proc_5_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(proc_5_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(proc_5_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(proc_5_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(proc_5_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(proc_5_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(proc_5_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(proc_5_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(proc_5_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(proc_5_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(proc_5_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(proc_5_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(proc_5_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(proc_5_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(proc_5_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(proc_5_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(proc_5_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(proc_5_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(proc_5_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(proc_5_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(proc_5_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(proc_5_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(proc_5_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(proc_5_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(proc_5_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(proc_5_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(proc_5_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(proc_5_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(proc_5_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(proc_5_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(proc_5_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(proc_5_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(proc_5_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(proc_5_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(proc_5_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(proc_5_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(proc_5_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(proc_5_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(proc_5_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(proc_5_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(proc_5_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(proc_5_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(proc_5_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(proc_5_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(proc_5_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(proc_5_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(proc_5_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(proc_5_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(proc_5_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(proc_5_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(proc_5_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(proc_5_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(proc_5_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(proc_5_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(proc_5_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(proc_5_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(proc_5_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(proc_5_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(proc_5_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(proc_5_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(proc_5_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(proc_5_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(proc_5_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(proc_5_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(proc_5_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(proc_5_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(proc_5_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(proc_5_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(proc_5_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(proc_5_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(proc_5_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(proc_5_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(proc_5_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(proc_5_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(proc_5_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(proc_5_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(proc_5_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(proc_5_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(proc_5_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(proc_5_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(proc_5_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(proc_5_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(proc_5_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(proc_5_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(proc_5_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(proc_5_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(proc_5_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(proc_5_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(proc_5_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(proc_5_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(proc_5_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(proc_5_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(proc_5_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(proc_5_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(proc_5_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(proc_5_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(proc_5_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(proc_5_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(proc_5_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(proc_5_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(proc_5_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(proc_5_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(proc_5_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(proc_5_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(proc_5_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(proc_5_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(proc_5_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(proc_5_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(proc_5_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(proc_5_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(proc_5_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(proc_5_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(proc_5_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(proc_5_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(proc_5_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(proc_5_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(proc_5_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(proc_5_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(proc_5_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(proc_5_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(proc_5_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(proc_5_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(proc_5_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(proc_5_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(proc_5_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(proc_5_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(proc_5_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(proc_5_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(proc_5_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(proc_5_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(proc_5_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(proc_5_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(proc_5_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(proc_5_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(proc_5_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(proc_5_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(proc_5_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(proc_5_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(proc_5_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(proc_5_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(proc_5_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(proc_5_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(proc_5_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(proc_5_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(proc_5_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(proc_5_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(proc_5_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(proc_5_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(proc_5_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(proc_5_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(proc_5_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(proc_5_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(proc_5_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_header_0(proc_5_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(proc_5_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(proc_5_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(proc_5_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(proc_5_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(proc_5_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(proc_5_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(proc_5_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(proc_5_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(proc_5_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(proc_5_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(proc_5_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(proc_5_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(proc_5_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(proc_5_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(proc_5_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(proc_5_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(proc_5_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(proc_5_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(proc_5_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(proc_5_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(proc_5_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_in_valid(proc_5_io_pipe_phv_in_valid),
    .io_pipe_phv_in_last(proc_5_io_pipe_phv_in_last),
    .io_pipe_phv_out_data_0(proc_5_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(proc_5_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(proc_5_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(proc_5_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(proc_5_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(proc_5_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(proc_5_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(proc_5_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(proc_5_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(proc_5_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(proc_5_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(proc_5_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(proc_5_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(proc_5_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(proc_5_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(proc_5_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(proc_5_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(proc_5_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(proc_5_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(proc_5_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(proc_5_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(proc_5_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(proc_5_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(proc_5_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(proc_5_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(proc_5_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(proc_5_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(proc_5_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(proc_5_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(proc_5_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(proc_5_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(proc_5_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(proc_5_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(proc_5_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(proc_5_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(proc_5_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(proc_5_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(proc_5_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(proc_5_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(proc_5_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(proc_5_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(proc_5_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(proc_5_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(proc_5_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(proc_5_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(proc_5_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(proc_5_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(proc_5_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(proc_5_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(proc_5_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(proc_5_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(proc_5_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(proc_5_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(proc_5_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(proc_5_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(proc_5_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(proc_5_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(proc_5_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(proc_5_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(proc_5_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(proc_5_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(proc_5_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(proc_5_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(proc_5_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(proc_5_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(proc_5_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(proc_5_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(proc_5_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(proc_5_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(proc_5_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(proc_5_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(proc_5_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(proc_5_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(proc_5_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(proc_5_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(proc_5_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(proc_5_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(proc_5_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(proc_5_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(proc_5_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(proc_5_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(proc_5_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(proc_5_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(proc_5_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(proc_5_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(proc_5_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(proc_5_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(proc_5_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(proc_5_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(proc_5_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(proc_5_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(proc_5_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(proc_5_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(proc_5_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(proc_5_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(proc_5_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(proc_5_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(proc_5_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(proc_5_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(proc_5_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(proc_5_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(proc_5_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(proc_5_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(proc_5_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(proc_5_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(proc_5_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(proc_5_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(proc_5_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(proc_5_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(proc_5_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(proc_5_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(proc_5_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(proc_5_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(proc_5_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(proc_5_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(proc_5_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(proc_5_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(proc_5_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(proc_5_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(proc_5_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(proc_5_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(proc_5_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(proc_5_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(proc_5_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(proc_5_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(proc_5_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(proc_5_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(proc_5_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(proc_5_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(proc_5_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(proc_5_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(proc_5_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(proc_5_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(proc_5_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(proc_5_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(proc_5_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(proc_5_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(proc_5_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(proc_5_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(proc_5_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(proc_5_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(proc_5_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(proc_5_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(proc_5_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(proc_5_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(proc_5_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(proc_5_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(proc_5_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(proc_5_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(proc_5_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(proc_5_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(proc_5_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(proc_5_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(proc_5_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(proc_5_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(proc_5_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(proc_5_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(proc_5_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(proc_5_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(proc_5_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_header_0(proc_5_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(proc_5_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(proc_5_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(proc_5_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(proc_5_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(proc_5_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(proc_5_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(proc_5_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(proc_5_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(proc_5_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(proc_5_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(proc_5_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(proc_5_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(proc_5_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(proc_5_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(proc_5_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(proc_5_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(proc_5_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(proc_5_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(proc_5_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(proc_5_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_valid(proc_5_io_pipe_phv_out_valid),
    .io_pipe_phv_out_last(proc_5_io_pipe_phv_out_last)
  );
  Processor proc_6 ( // @[ipsa.scala 56:25]
    .clock(proc_6_clock),
    .io_pipe_phv_in_data_0(proc_6_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(proc_6_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(proc_6_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(proc_6_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(proc_6_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(proc_6_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(proc_6_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(proc_6_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(proc_6_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(proc_6_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(proc_6_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(proc_6_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(proc_6_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(proc_6_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(proc_6_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(proc_6_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(proc_6_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(proc_6_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(proc_6_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(proc_6_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(proc_6_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(proc_6_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(proc_6_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(proc_6_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(proc_6_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(proc_6_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(proc_6_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(proc_6_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(proc_6_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(proc_6_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(proc_6_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(proc_6_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(proc_6_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(proc_6_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(proc_6_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(proc_6_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(proc_6_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(proc_6_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(proc_6_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(proc_6_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(proc_6_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(proc_6_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(proc_6_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(proc_6_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(proc_6_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(proc_6_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(proc_6_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(proc_6_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(proc_6_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(proc_6_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(proc_6_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(proc_6_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(proc_6_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(proc_6_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(proc_6_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(proc_6_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(proc_6_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(proc_6_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(proc_6_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(proc_6_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(proc_6_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(proc_6_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(proc_6_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(proc_6_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(proc_6_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(proc_6_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(proc_6_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(proc_6_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(proc_6_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(proc_6_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(proc_6_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(proc_6_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(proc_6_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(proc_6_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(proc_6_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(proc_6_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(proc_6_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(proc_6_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(proc_6_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(proc_6_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(proc_6_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(proc_6_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(proc_6_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(proc_6_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(proc_6_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(proc_6_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(proc_6_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(proc_6_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(proc_6_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(proc_6_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(proc_6_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(proc_6_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(proc_6_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(proc_6_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(proc_6_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(proc_6_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(proc_6_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(proc_6_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(proc_6_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(proc_6_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(proc_6_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(proc_6_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(proc_6_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(proc_6_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(proc_6_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(proc_6_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(proc_6_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(proc_6_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(proc_6_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(proc_6_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(proc_6_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(proc_6_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(proc_6_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(proc_6_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(proc_6_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(proc_6_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(proc_6_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(proc_6_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(proc_6_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(proc_6_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(proc_6_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(proc_6_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(proc_6_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(proc_6_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(proc_6_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(proc_6_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(proc_6_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(proc_6_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(proc_6_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(proc_6_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(proc_6_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(proc_6_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(proc_6_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(proc_6_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(proc_6_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(proc_6_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(proc_6_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(proc_6_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(proc_6_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(proc_6_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(proc_6_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(proc_6_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(proc_6_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(proc_6_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(proc_6_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(proc_6_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(proc_6_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(proc_6_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(proc_6_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(proc_6_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(proc_6_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(proc_6_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(proc_6_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(proc_6_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(proc_6_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(proc_6_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(proc_6_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(proc_6_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(proc_6_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(proc_6_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_header_0(proc_6_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(proc_6_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(proc_6_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(proc_6_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(proc_6_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(proc_6_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(proc_6_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(proc_6_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(proc_6_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(proc_6_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(proc_6_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(proc_6_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(proc_6_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(proc_6_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(proc_6_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(proc_6_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(proc_6_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(proc_6_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(proc_6_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(proc_6_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(proc_6_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(proc_6_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_in_valid(proc_6_io_pipe_phv_in_valid),
    .io_pipe_phv_in_last(proc_6_io_pipe_phv_in_last),
    .io_pipe_phv_out_data_0(proc_6_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(proc_6_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(proc_6_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(proc_6_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(proc_6_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(proc_6_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(proc_6_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(proc_6_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(proc_6_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(proc_6_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(proc_6_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(proc_6_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(proc_6_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(proc_6_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(proc_6_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(proc_6_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(proc_6_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(proc_6_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(proc_6_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(proc_6_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(proc_6_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(proc_6_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(proc_6_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(proc_6_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(proc_6_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(proc_6_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(proc_6_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(proc_6_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(proc_6_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(proc_6_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(proc_6_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(proc_6_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(proc_6_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(proc_6_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(proc_6_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(proc_6_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(proc_6_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(proc_6_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(proc_6_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(proc_6_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(proc_6_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(proc_6_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(proc_6_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(proc_6_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(proc_6_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(proc_6_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(proc_6_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(proc_6_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(proc_6_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(proc_6_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(proc_6_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(proc_6_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(proc_6_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(proc_6_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(proc_6_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(proc_6_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(proc_6_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(proc_6_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(proc_6_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(proc_6_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(proc_6_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(proc_6_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(proc_6_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(proc_6_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(proc_6_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(proc_6_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(proc_6_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(proc_6_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(proc_6_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(proc_6_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(proc_6_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(proc_6_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(proc_6_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(proc_6_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(proc_6_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(proc_6_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(proc_6_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(proc_6_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(proc_6_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(proc_6_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(proc_6_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(proc_6_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(proc_6_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(proc_6_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(proc_6_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(proc_6_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(proc_6_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(proc_6_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(proc_6_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(proc_6_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(proc_6_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(proc_6_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(proc_6_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(proc_6_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(proc_6_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(proc_6_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(proc_6_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(proc_6_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(proc_6_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(proc_6_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(proc_6_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(proc_6_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(proc_6_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(proc_6_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(proc_6_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(proc_6_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(proc_6_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(proc_6_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(proc_6_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(proc_6_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(proc_6_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(proc_6_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(proc_6_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(proc_6_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(proc_6_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(proc_6_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(proc_6_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(proc_6_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(proc_6_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(proc_6_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(proc_6_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(proc_6_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(proc_6_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(proc_6_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(proc_6_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(proc_6_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(proc_6_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(proc_6_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(proc_6_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(proc_6_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(proc_6_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(proc_6_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(proc_6_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(proc_6_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(proc_6_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(proc_6_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(proc_6_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(proc_6_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(proc_6_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(proc_6_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(proc_6_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(proc_6_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(proc_6_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(proc_6_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(proc_6_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(proc_6_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(proc_6_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(proc_6_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(proc_6_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(proc_6_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(proc_6_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(proc_6_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(proc_6_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(proc_6_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(proc_6_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(proc_6_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(proc_6_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(proc_6_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(proc_6_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(proc_6_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_header_0(proc_6_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(proc_6_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(proc_6_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(proc_6_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(proc_6_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(proc_6_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(proc_6_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(proc_6_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(proc_6_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(proc_6_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(proc_6_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(proc_6_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(proc_6_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(proc_6_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(proc_6_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(proc_6_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(proc_6_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(proc_6_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(proc_6_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(proc_6_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(proc_6_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_valid(proc_6_io_pipe_phv_out_valid),
    .io_pipe_phv_out_last(proc_6_io_pipe_phv_out_last)
  );
  Processor proc_7 ( // @[ipsa.scala 56:25]
    .clock(proc_7_clock),
    .io_pipe_phv_in_data_0(proc_7_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(proc_7_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(proc_7_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(proc_7_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(proc_7_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(proc_7_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(proc_7_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(proc_7_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(proc_7_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(proc_7_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(proc_7_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(proc_7_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(proc_7_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(proc_7_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(proc_7_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(proc_7_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(proc_7_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(proc_7_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(proc_7_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(proc_7_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(proc_7_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(proc_7_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(proc_7_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(proc_7_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(proc_7_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(proc_7_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(proc_7_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(proc_7_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(proc_7_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(proc_7_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(proc_7_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(proc_7_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(proc_7_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(proc_7_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(proc_7_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(proc_7_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(proc_7_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(proc_7_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(proc_7_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(proc_7_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(proc_7_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(proc_7_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(proc_7_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(proc_7_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(proc_7_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(proc_7_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(proc_7_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(proc_7_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(proc_7_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(proc_7_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(proc_7_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(proc_7_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(proc_7_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(proc_7_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(proc_7_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(proc_7_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(proc_7_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(proc_7_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(proc_7_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(proc_7_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(proc_7_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(proc_7_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(proc_7_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(proc_7_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(proc_7_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(proc_7_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(proc_7_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(proc_7_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(proc_7_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(proc_7_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(proc_7_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(proc_7_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(proc_7_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(proc_7_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(proc_7_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(proc_7_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(proc_7_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(proc_7_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(proc_7_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(proc_7_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(proc_7_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(proc_7_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(proc_7_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(proc_7_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(proc_7_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(proc_7_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(proc_7_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(proc_7_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(proc_7_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(proc_7_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(proc_7_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(proc_7_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(proc_7_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(proc_7_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(proc_7_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(proc_7_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(proc_7_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(proc_7_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(proc_7_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(proc_7_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(proc_7_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(proc_7_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(proc_7_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(proc_7_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(proc_7_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(proc_7_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(proc_7_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(proc_7_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(proc_7_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(proc_7_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(proc_7_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(proc_7_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(proc_7_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(proc_7_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(proc_7_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(proc_7_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(proc_7_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(proc_7_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(proc_7_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(proc_7_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(proc_7_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(proc_7_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(proc_7_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(proc_7_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(proc_7_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(proc_7_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(proc_7_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(proc_7_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(proc_7_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(proc_7_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(proc_7_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(proc_7_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(proc_7_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(proc_7_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(proc_7_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(proc_7_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(proc_7_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(proc_7_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(proc_7_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(proc_7_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(proc_7_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(proc_7_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(proc_7_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(proc_7_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(proc_7_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(proc_7_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(proc_7_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(proc_7_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(proc_7_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(proc_7_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(proc_7_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(proc_7_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(proc_7_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(proc_7_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(proc_7_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(proc_7_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(proc_7_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(proc_7_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(proc_7_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(proc_7_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_header_0(proc_7_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(proc_7_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(proc_7_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(proc_7_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(proc_7_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(proc_7_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(proc_7_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(proc_7_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(proc_7_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(proc_7_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(proc_7_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(proc_7_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(proc_7_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(proc_7_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(proc_7_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(proc_7_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(proc_7_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(proc_7_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(proc_7_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(proc_7_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(proc_7_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(proc_7_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_in_valid(proc_7_io_pipe_phv_in_valid),
    .io_pipe_phv_in_last(proc_7_io_pipe_phv_in_last),
    .io_pipe_phv_out_data_0(proc_7_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(proc_7_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(proc_7_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(proc_7_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(proc_7_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(proc_7_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(proc_7_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(proc_7_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(proc_7_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(proc_7_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(proc_7_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(proc_7_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(proc_7_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(proc_7_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(proc_7_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(proc_7_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(proc_7_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(proc_7_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(proc_7_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(proc_7_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(proc_7_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(proc_7_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(proc_7_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(proc_7_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(proc_7_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(proc_7_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(proc_7_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(proc_7_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(proc_7_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(proc_7_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(proc_7_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(proc_7_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(proc_7_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(proc_7_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(proc_7_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(proc_7_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(proc_7_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(proc_7_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(proc_7_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(proc_7_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(proc_7_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(proc_7_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(proc_7_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(proc_7_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(proc_7_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(proc_7_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(proc_7_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(proc_7_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(proc_7_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(proc_7_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(proc_7_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(proc_7_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(proc_7_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(proc_7_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(proc_7_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(proc_7_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(proc_7_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(proc_7_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(proc_7_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(proc_7_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(proc_7_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(proc_7_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(proc_7_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(proc_7_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(proc_7_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(proc_7_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(proc_7_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(proc_7_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(proc_7_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(proc_7_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(proc_7_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(proc_7_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(proc_7_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(proc_7_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(proc_7_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(proc_7_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(proc_7_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(proc_7_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(proc_7_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(proc_7_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(proc_7_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(proc_7_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(proc_7_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(proc_7_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(proc_7_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(proc_7_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(proc_7_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(proc_7_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(proc_7_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(proc_7_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(proc_7_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(proc_7_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(proc_7_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(proc_7_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(proc_7_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(proc_7_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(proc_7_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(proc_7_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(proc_7_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(proc_7_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(proc_7_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(proc_7_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(proc_7_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(proc_7_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(proc_7_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(proc_7_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(proc_7_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(proc_7_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(proc_7_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(proc_7_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(proc_7_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(proc_7_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(proc_7_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(proc_7_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(proc_7_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(proc_7_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(proc_7_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(proc_7_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(proc_7_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(proc_7_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(proc_7_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(proc_7_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(proc_7_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(proc_7_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(proc_7_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(proc_7_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(proc_7_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(proc_7_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(proc_7_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(proc_7_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(proc_7_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(proc_7_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(proc_7_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(proc_7_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(proc_7_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(proc_7_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(proc_7_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(proc_7_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(proc_7_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(proc_7_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(proc_7_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(proc_7_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(proc_7_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(proc_7_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(proc_7_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(proc_7_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(proc_7_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(proc_7_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(proc_7_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(proc_7_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(proc_7_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(proc_7_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(proc_7_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(proc_7_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(proc_7_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(proc_7_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(proc_7_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(proc_7_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(proc_7_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(proc_7_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_header_0(proc_7_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(proc_7_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(proc_7_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(proc_7_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(proc_7_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(proc_7_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(proc_7_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(proc_7_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(proc_7_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(proc_7_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(proc_7_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(proc_7_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(proc_7_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(proc_7_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(proc_7_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(proc_7_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(proc_7_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(proc_7_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(proc_7_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(proc_7_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(proc_7_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_valid(proc_7_io_pipe_phv_out_valid),
    .io_pipe_phv_out_last(proc_7_io_pipe_phv_out_last)
  );
  Processor proc_8 ( // @[ipsa.scala 56:25]
    .clock(proc_8_clock),
    .io_pipe_phv_in_data_0(proc_8_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(proc_8_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(proc_8_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(proc_8_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(proc_8_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(proc_8_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(proc_8_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(proc_8_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(proc_8_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(proc_8_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(proc_8_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(proc_8_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(proc_8_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(proc_8_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(proc_8_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(proc_8_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(proc_8_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(proc_8_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(proc_8_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(proc_8_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(proc_8_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(proc_8_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(proc_8_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(proc_8_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(proc_8_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(proc_8_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(proc_8_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(proc_8_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(proc_8_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(proc_8_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(proc_8_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(proc_8_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(proc_8_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(proc_8_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(proc_8_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(proc_8_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(proc_8_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(proc_8_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(proc_8_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(proc_8_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(proc_8_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(proc_8_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(proc_8_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(proc_8_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(proc_8_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(proc_8_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(proc_8_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(proc_8_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(proc_8_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(proc_8_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(proc_8_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(proc_8_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(proc_8_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(proc_8_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(proc_8_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(proc_8_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(proc_8_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(proc_8_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(proc_8_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(proc_8_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(proc_8_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(proc_8_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(proc_8_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(proc_8_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(proc_8_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(proc_8_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(proc_8_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(proc_8_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(proc_8_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(proc_8_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(proc_8_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(proc_8_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(proc_8_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(proc_8_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(proc_8_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(proc_8_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(proc_8_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(proc_8_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(proc_8_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(proc_8_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(proc_8_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(proc_8_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(proc_8_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(proc_8_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(proc_8_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(proc_8_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(proc_8_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(proc_8_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(proc_8_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(proc_8_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(proc_8_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(proc_8_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(proc_8_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(proc_8_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(proc_8_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(proc_8_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(proc_8_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(proc_8_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(proc_8_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(proc_8_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(proc_8_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(proc_8_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(proc_8_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(proc_8_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(proc_8_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(proc_8_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(proc_8_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(proc_8_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(proc_8_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(proc_8_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(proc_8_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(proc_8_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(proc_8_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(proc_8_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(proc_8_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(proc_8_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(proc_8_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(proc_8_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(proc_8_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(proc_8_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(proc_8_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(proc_8_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(proc_8_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(proc_8_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(proc_8_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(proc_8_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(proc_8_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(proc_8_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(proc_8_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(proc_8_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(proc_8_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(proc_8_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(proc_8_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(proc_8_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(proc_8_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(proc_8_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(proc_8_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(proc_8_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(proc_8_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(proc_8_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(proc_8_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(proc_8_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(proc_8_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(proc_8_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(proc_8_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(proc_8_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(proc_8_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(proc_8_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(proc_8_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(proc_8_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(proc_8_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(proc_8_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(proc_8_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(proc_8_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(proc_8_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(proc_8_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(proc_8_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(proc_8_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(proc_8_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(proc_8_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_header_0(proc_8_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(proc_8_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(proc_8_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(proc_8_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(proc_8_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(proc_8_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(proc_8_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(proc_8_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(proc_8_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(proc_8_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(proc_8_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(proc_8_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(proc_8_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(proc_8_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(proc_8_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(proc_8_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(proc_8_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(proc_8_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(proc_8_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(proc_8_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(proc_8_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(proc_8_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_in_valid(proc_8_io_pipe_phv_in_valid),
    .io_pipe_phv_in_last(proc_8_io_pipe_phv_in_last),
    .io_pipe_phv_out_data_0(proc_8_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(proc_8_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(proc_8_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(proc_8_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(proc_8_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(proc_8_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(proc_8_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(proc_8_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(proc_8_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(proc_8_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(proc_8_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(proc_8_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(proc_8_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(proc_8_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(proc_8_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(proc_8_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(proc_8_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(proc_8_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(proc_8_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(proc_8_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(proc_8_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(proc_8_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(proc_8_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(proc_8_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(proc_8_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(proc_8_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(proc_8_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(proc_8_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(proc_8_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(proc_8_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(proc_8_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(proc_8_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(proc_8_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(proc_8_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(proc_8_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(proc_8_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(proc_8_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(proc_8_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(proc_8_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(proc_8_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(proc_8_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(proc_8_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(proc_8_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(proc_8_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(proc_8_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(proc_8_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(proc_8_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(proc_8_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(proc_8_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(proc_8_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(proc_8_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(proc_8_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(proc_8_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(proc_8_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(proc_8_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(proc_8_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(proc_8_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(proc_8_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(proc_8_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(proc_8_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(proc_8_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(proc_8_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(proc_8_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(proc_8_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(proc_8_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(proc_8_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(proc_8_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(proc_8_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(proc_8_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(proc_8_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(proc_8_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(proc_8_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(proc_8_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(proc_8_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(proc_8_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(proc_8_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(proc_8_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(proc_8_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(proc_8_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(proc_8_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(proc_8_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(proc_8_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(proc_8_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(proc_8_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(proc_8_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(proc_8_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(proc_8_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(proc_8_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(proc_8_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(proc_8_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(proc_8_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(proc_8_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(proc_8_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(proc_8_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(proc_8_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(proc_8_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(proc_8_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(proc_8_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(proc_8_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(proc_8_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(proc_8_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(proc_8_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(proc_8_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(proc_8_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(proc_8_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(proc_8_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(proc_8_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(proc_8_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(proc_8_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(proc_8_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(proc_8_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(proc_8_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(proc_8_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(proc_8_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(proc_8_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(proc_8_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(proc_8_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(proc_8_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(proc_8_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(proc_8_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(proc_8_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(proc_8_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(proc_8_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(proc_8_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(proc_8_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(proc_8_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(proc_8_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(proc_8_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(proc_8_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(proc_8_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(proc_8_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(proc_8_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(proc_8_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(proc_8_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(proc_8_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(proc_8_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(proc_8_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(proc_8_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(proc_8_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(proc_8_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(proc_8_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(proc_8_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(proc_8_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(proc_8_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(proc_8_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(proc_8_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(proc_8_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(proc_8_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(proc_8_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(proc_8_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(proc_8_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(proc_8_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(proc_8_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(proc_8_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(proc_8_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(proc_8_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(proc_8_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(proc_8_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(proc_8_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(proc_8_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_header_0(proc_8_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(proc_8_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(proc_8_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(proc_8_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(proc_8_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(proc_8_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(proc_8_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(proc_8_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(proc_8_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(proc_8_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(proc_8_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(proc_8_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(proc_8_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(proc_8_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(proc_8_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(proc_8_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(proc_8_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(proc_8_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(proc_8_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(proc_8_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(proc_8_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_valid(proc_8_io_pipe_phv_out_valid),
    .io_pipe_phv_out_last(proc_8_io_pipe_phv_out_last)
  );
  Processor proc_9 ( // @[ipsa.scala 56:25]
    .clock(proc_9_clock),
    .io_pipe_phv_in_data_0(proc_9_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(proc_9_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(proc_9_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(proc_9_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(proc_9_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(proc_9_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(proc_9_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(proc_9_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(proc_9_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(proc_9_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(proc_9_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(proc_9_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(proc_9_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(proc_9_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(proc_9_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(proc_9_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(proc_9_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(proc_9_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(proc_9_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(proc_9_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(proc_9_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(proc_9_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(proc_9_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(proc_9_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(proc_9_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(proc_9_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(proc_9_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(proc_9_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(proc_9_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(proc_9_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(proc_9_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(proc_9_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(proc_9_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(proc_9_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(proc_9_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(proc_9_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(proc_9_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(proc_9_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(proc_9_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(proc_9_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(proc_9_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(proc_9_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(proc_9_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(proc_9_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(proc_9_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(proc_9_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(proc_9_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(proc_9_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(proc_9_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(proc_9_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(proc_9_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(proc_9_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(proc_9_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(proc_9_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(proc_9_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(proc_9_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(proc_9_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(proc_9_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(proc_9_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(proc_9_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(proc_9_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(proc_9_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(proc_9_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(proc_9_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(proc_9_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(proc_9_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(proc_9_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(proc_9_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(proc_9_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(proc_9_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(proc_9_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(proc_9_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(proc_9_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(proc_9_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(proc_9_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(proc_9_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(proc_9_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(proc_9_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(proc_9_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(proc_9_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(proc_9_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(proc_9_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(proc_9_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(proc_9_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(proc_9_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(proc_9_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(proc_9_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(proc_9_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(proc_9_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(proc_9_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(proc_9_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(proc_9_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(proc_9_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(proc_9_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(proc_9_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(proc_9_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(proc_9_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(proc_9_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(proc_9_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(proc_9_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(proc_9_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(proc_9_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(proc_9_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(proc_9_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(proc_9_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(proc_9_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(proc_9_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(proc_9_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(proc_9_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(proc_9_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(proc_9_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(proc_9_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(proc_9_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(proc_9_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(proc_9_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(proc_9_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(proc_9_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(proc_9_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(proc_9_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(proc_9_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(proc_9_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(proc_9_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(proc_9_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(proc_9_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(proc_9_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(proc_9_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(proc_9_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(proc_9_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(proc_9_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(proc_9_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(proc_9_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(proc_9_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(proc_9_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(proc_9_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(proc_9_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(proc_9_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(proc_9_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(proc_9_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(proc_9_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(proc_9_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(proc_9_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(proc_9_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(proc_9_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(proc_9_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(proc_9_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(proc_9_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(proc_9_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(proc_9_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(proc_9_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(proc_9_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(proc_9_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(proc_9_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(proc_9_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(proc_9_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(proc_9_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(proc_9_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(proc_9_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(proc_9_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(proc_9_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(proc_9_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_header_0(proc_9_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(proc_9_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(proc_9_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(proc_9_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(proc_9_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(proc_9_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(proc_9_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(proc_9_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(proc_9_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(proc_9_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(proc_9_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(proc_9_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(proc_9_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(proc_9_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(proc_9_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(proc_9_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(proc_9_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(proc_9_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(proc_9_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(proc_9_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(proc_9_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(proc_9_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_in_valid(proc_9_io_pipe_phv_in_valid),
    .io_pipe_phv_in_last(proc_9_io_pipe_phv_in_last),
    .io_pipe_phv_out_data_0(proc_9_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(proc_9_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(proc_9_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(proc_9_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(proc_9_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(proc_9_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(proc_9_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(proc_9_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(proc_9_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(proc_9_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(proc_9_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(proc_9_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(proc_9_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(proc_9_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(proc_9_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(proc_9_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(proc_9_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(proc_9_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(proc_9_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(proc_9_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(proc_9_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(proc_9_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(proc_9_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(proc_9_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(proc_9_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(proc_9_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(proc_9_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(proc_9_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(proc_9_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(proc_9_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(proc_9_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(proc_9_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(proc_9_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(proc_9_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(proc_9_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(proc_9_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(proc_9_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(proc_9_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(proc_9_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(proc_9_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(proc_9_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(proc_9_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(proc_9_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(proc_9_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(proc_9_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(proc_9_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(proc_9_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(proc_9_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(proc_9_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(proc_9_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(proc_9_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(proc_9_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(proc_9_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(proc_9_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(proc_9_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(proc_9_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(proc_9_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(proc_9_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(proc_9_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(proc_9_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(proc_9_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(proc_9_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(proc_9_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(proc_9_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(proc_9_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(proc_9_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(proc_9_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(proc_9_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(proc_9_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(proc_9_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(proc_9_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(proc_9_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(proc_9_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(proc_9_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(proc_9_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(proc_9_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(proc_9_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(proc_9_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(proc_9_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(proc_9_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(proc_9_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(proc_9_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(proc_9_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(proc_9_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(proc_9_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(proc_9_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(proc_9_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(proc_9_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(proc_9_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(proc_9_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(proc_9_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(proc_9_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(proc_9_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(proc_9_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(proc_9_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(proc_9_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(proc_9_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(proc_9_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(proc_9_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(proc_9_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(proc_9_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(proc_9_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(proc_9_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(proc_9_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(proc_9_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(proc_9_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(proc_9_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(proc_9_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(proc_9_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(proc_9_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(proc_9_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(proc_9_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(proc_9_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(proc_9_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(proc_9_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(proc_9_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(proc_9_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(proc_9_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(proc_9_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(proc_9_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(proc_9_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(proc_9_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(proc_9_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(proc_9_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(proc_9_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(proc_9_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(proc_9_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(proc_9_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(proc_9_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(proc_9_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(proc_9_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(proc_9_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(proc_9_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(proc_9_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(proc_9_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(proc_9_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(proc_9_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(proc_9_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(proc_9_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(proc_9_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(proc_9_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(proc_9_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(proc_9_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(proc_9_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(proc_9_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(proc_9_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(proc_9_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(proc_9_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(proc_9_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(proc_9_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(proc_9_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(proc_9_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(proc_9_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(proc_9_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(proc_9_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(proc_9_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(proc_9_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(proc_9_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(proc_9_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(proc_9_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_header_0(proc_9_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(proc_9_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(proc_9_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(proc_9_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(proc_9_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(proc_9_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(proc_9_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(proc_9_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(proc_9_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(proc_9_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(proc_9_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(proc_9_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(proc_9_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(proc_9_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(proc_9_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(proc_9_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(proc_9_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(proc_9_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(proc_9_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(proc_9_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(proc_9_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_valid(proc_9_io_pipe_phv_out_valid),
    .io_pipe_phv_out_last(proc_9_io_pipe_phv_out_last)
  );
  Processor proc_10 ( // @[ipsa.scala 56:25]
    .clock(proc_10_clock),
    .io_pipe_phv_in_data_0(proc_10_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(proc_10_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(proc_10_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(proc_10_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(proc_10_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(proc_10_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(proc_10_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(proc_10_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(proc_10_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(proc_10_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(proc_10_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(proc_10_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(proc_10_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(proc_10_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(proc_10_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(proc_10_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(proc_10_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(proc_10_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(proc_10_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(proc_10_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(proc_10_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(proc_10_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(proc_10_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(proc_10_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(proc_10_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(proc_10_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(proc_10_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(proc_10_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(proc_10_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(proc_10_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(proc_10_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(proc_10_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(proc_10_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(proc_10_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(proc_10_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(proc_10_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(proc_10_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(proc_10_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(proc_10_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(proc_10_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(proc_10_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(proc_10_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(proc_10_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(proc_10_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(proc_10_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(proc_10_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(proc_10_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(proc_10_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(proc_10_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(proc_10_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(proc_10_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(proc_10_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(proc_10_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(proc_10_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(proc_10_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(proc_10_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(proc_10_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(proc_10_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(proc_10_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(proc_10_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(proc_10_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(proc_10_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(proc_10_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(proc_10_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(proc_10_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(proc_10_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(proc_10_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(proc_10_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(proc_10_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(proc_10_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(proc_10_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(proc_10_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(proc_10_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(proc_10_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(proc_10_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(proc_10_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(proc_10_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(proc_10_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(proc_10_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(proc_10_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(proc_10_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(proc_10_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(proc_10_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(proc_10_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(proc_10_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(proc_10_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(proc_10_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(proc_10_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(proc_10_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(proc_10_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(proc_10_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(proc_10_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(proc_10_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(proc_10_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(proc_10_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(proc_10_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(proc_10_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(proc_10_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(proc_10_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(proc_10_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(proc_10_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(proc_10_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(proc_10_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(proc_10_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(proc_10_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(proc_10_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(proc_10_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(proc_10_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(proc_10_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(proc_10_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(proc_10_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(proc_10_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(proc_10_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(proc_10_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(proc_10_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(proc_10_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(proc_10_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(proc_10_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(proc_10_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(proc_10_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(proc_10_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(proc_10_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(proc_10_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(proc_10_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(proc_10_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(proc_10_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(proc_10_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(proc_10_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(proc_10_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(proc_10_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(proc_10_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(proc_10_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(proc_10_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(proc_10_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(proc_10_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(proc_10_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(proc_10_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(proc_10_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(proc_10_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(proc_10_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(proc_10_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(proc_10_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(proc_10_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(proc_10_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(proc_10_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(proc_10_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(proc_10_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(proc_10_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(proc_10_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(proc_10_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(proc_10_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(proc_10_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(proc_10_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(proc_10_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(proc_10_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(proc_10_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(proc_10_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(proc_10_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(proc_10_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(proc_10_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_header_0(proc_10_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(proc_10_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(proc_10_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(proc_10_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(proc_10_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(proc_10_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(proc_10_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(proc_10_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(proc_10_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(proc_10_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(proc_10_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(proc_10_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(proc_10_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(proc_10_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(proc_10_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(proc_10_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(proc_10_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(proc_10_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(proc_10_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(proc_10_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(proc_10_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(proc_10_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_in_valid(proc_10_io_pipe_phv_in_valid),
    .io_pipe_phv_in_last(proc_10_io_pipe_phv_in_last),
    .io_pipe_phv_out_data_0(proc_10_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(proc_10_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(proc_10_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(proc_10_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(proc_10_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(proc_10_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(proc_10_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(proc_10_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(proc_10_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(proc_10_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(proc_10_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(proc_10_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(proc_10_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(proc_10_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(proc_10_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(proc_10_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(proc_10_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(proc_10_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(proc_10_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(proc_10_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(proc_10_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(proc_10_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(proc_10_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(proc_10_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(proc_10_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(proc_10_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(proc_10_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(proc_10_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(proc_10_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(proc_10_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(proc_10_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(proc_10_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(proc_10_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(proc_10_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(proc_10_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(proc_10_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(proc_10_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(proc_10_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(proc_10_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(proc_10_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(proc_10_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(proc_10_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(proc_10_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(proc_10_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(proc_10_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(proc_10_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(proc_10_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(proc_10_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(proc_10_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(proc_10_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(proc_10_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(proc_10_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(proc_10_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(proc_10_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(proc_10_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(proc_10_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(proc_10_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(proc_10_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(proc_10_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(proc_10_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(proc_10_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(proc_10_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(proc_10_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(proc_10_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(proc_10_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(proc_10_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(proc_10_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(proc_10_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(proc_10_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(proc_10_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(proc_10_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(proc_10_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(proc_10_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(proc_10_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(proc_10_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(proc_10_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(proc_10_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(proc_10_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(proc_10_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(proc_10_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(proc_10_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(proc_10_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(proc_10_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(proc_10_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(proc_10_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(proc_10_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(proc_10_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(proc_10_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(proc_10_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(proc_10_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(proc_10_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(proc_10_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(proc_10_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(proc_10_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(proc_10_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(proc_10_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(proc_10_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(proc_10_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(proc_10_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(proc_10_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(proc_10_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(proc_10_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(proc_10_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(proc_10_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(proc_10_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(proc_10_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(proc_10_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(proc_10_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(proc_10_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(proc_10_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(proc_10_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(proc_10_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(proc_10_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(proc_10_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(proc_10_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(proc_10_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(proc_10_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(proc_10_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(proc_10_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(proc_10_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(proc_10_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(proc_10_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(proc_10_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(proc_10_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(proc_10_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(proc_10_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(proc_10_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(proc_10_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(proc_10_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(proc_10_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(proc_10_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(proc_10_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(proc_10_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(proc_10_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(proc_10_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(proc_10_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(proc_10_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(proc_10_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(proc_10_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(proc_10_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(proc_10_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(proc_10_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(proc_10_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(proc_10_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(proc_10_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(proc_10_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(proc_10_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(proc_10_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(proc_10_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(proc_10_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(proc_10_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(proc_10_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(proc_10_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(proc_10_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(proc_10_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(proc_10_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(proc_10_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(proc_10_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(proc_10_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(proc_10_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_header_0(proc_10_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(proc_10_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(proc_10_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(proc_10_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(proc_10_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(proc_10_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(proc_10_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(proc_10_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(proc_10_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(proc_10_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(proc_10_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(proc_10_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(proc_10_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(proc_10_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(proc_10_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(proc_10_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(proc_10_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(proc_10_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(proc_10_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(proc_10_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(proc_10_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_valid(proc_10_io_pipe_phv_out_valid),
    .io_pipe_phv_out_last(proc_10_io_pipe_phv_out_last)
  );
  Processor proc_11 ( // @[ipsa.scala 56:25]
    .clock(proc_11_clock),
    .io_pipe_phv_in_data_0(proc_11_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(proc_11_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(proc_11_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(proc_11_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(proc_11_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(proc_11_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(proc_11_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(proc_11_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(proc_11_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(proc_11_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(proc_11_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(proc_11_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(proc_11_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(proc_11_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(proc_11_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(proc_11_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(proc_11_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(proc_11_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(proc_11_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(proc_11_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(proc_11_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(proc_11_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(proc_11_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(proc_11_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(proc_11_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(proc_11_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(proc_11_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(proc_11_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(proc_11_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(proc_11_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(proc_11_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(proc_11_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(proc_11_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(proc_11_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(proc_11_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(proc_11_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(proc_11_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(proc_11_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(proc_11_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(proc_11_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(proc_11_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(proc_11_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(proc_11_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(proc_11_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(proc_11_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(proc_11_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(proc_11_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(proc_11_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(proc_11_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(proc_11_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(proc_11_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(proc_11_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(proc_11_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(proc_11_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(proc_11_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(proc_11_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(proc_11_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(proc_11_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(proc_11_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(proc_11_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(proc_11_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(proc_11_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(proc_11_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(proc_11_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(proc_11_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(proc_11_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(proc_11_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(proc_11_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(proc_11_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(proc_11_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(proc_11_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(proc_11_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(proc_11_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(proc_11_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(proc_11_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(proc_11_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(proc_11_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(proc_11_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(proc_11_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(proc_11_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(proc_11_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(proc_11_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(proc_11_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(proc_11_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(proc_11_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(proc_11_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(proc_11_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(proc_11_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(proc_11_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(proc_11_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(proc_11_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(proc_11_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(proc_11_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(proc_11_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(proc_11_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(proc_11_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(proc_11_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(proc_11_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(proc_11_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(proc_11_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(proc_11_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(proc_11_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(proc_11_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(proc_11_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(proc_11_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(proc_11_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(proc_11_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(proc_11_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(proc_11_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(proc_11_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(proc_11_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(proc_11_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(proc_11_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(proc_11_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(proc_11_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(proc_11_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(proc_11_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(proc_11_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(proc_11_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(proc_11_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(proc_11_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(proc_11_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(proc_11_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(proc_11_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(proc_11_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(proc_11_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(proc_11_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(proc_11_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(proc_11_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(proc_11_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(proc_11_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(proc_11_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(proc_11_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(proc_11_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(proc_11_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(proc_11_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(proc_11_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(proc_11_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(proc_11_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(proc_11_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(proc_11_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(proc_11_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(proc_11_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(proc_11_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(proc_11_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(proc_11_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(proc_11_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(proc_11_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(proc_11_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(proc_11_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(proc_11_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(proc_11_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(proc_11_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(proc_11_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(proc_11_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(proc_11_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(proc_11_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(proc_11_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(proc_11_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(proc_11_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_header_0(proc_11_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(proc_11_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(proc_11_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(proc_11_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(proc_11_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(proc_11_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(proc_11_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(proc_11_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(proc_11_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(proc_11_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(proc_11_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(proc_11_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(proc_11_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(proc_11_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(proc_11_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(proc_11_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(proc_11_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(proc_11_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(proc_11_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(proc_11_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(proc_11_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(proc_11_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_in_valid(proc_11_io_pipe_phv_in_valid),
    .io_pipe_phv_in_last(proc_11_io_pipe_phv_in_last),
    .io_pipe_phv_out_data_0(proc_11_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(proc_11_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(proc_11_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(proc_11_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(proc_11_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(proc_11_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(proc_11_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(proc_11_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(proc_11_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(proc_11_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(proc_11_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(proc_11_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(proc_11_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(proc_11_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(proc_11_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(proc_11_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(proc_11_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(proc_11_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(proc_11_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(proc_11_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(proc_11_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(proc_11_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(proc_11_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(proc_11_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(proc_11_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(proc_11_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(proc_11_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(proc_11_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(proc_11_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(proc_11_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(proc_11_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(proc_11_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(proc_11_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(proc_11_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(proc_11_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(proc_11_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(proc_11_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(proc_11_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(proc_11_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(proc_11_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(proc_11_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(proc_11_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(proc_11_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(proc_11_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(proc_11_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(proc_11_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(proc_11_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(proc_11_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(proc_11_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(proc_11_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(proc_11_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(proc_11_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(proc_11_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(proc_11_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(proc_11_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(proc_11_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(proc_11_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(proc_11_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(proc_11_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(proc_11_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(proc_11_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(proc_11_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(proc_11_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(proc_11_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(proc_11_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(proc_11_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(proc_11_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(proc_11_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(proc_11_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(proc_11_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(proc_11_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(proc_11_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(proc_11_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(proc_11_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(proc_11_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(proc_11_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(proc_11_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(proc_11_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(proc_11_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(proc_11_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(proc_11_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(proc_11_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(proc_11_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(proc_11_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(proc_11_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(proc_11_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(proc_11_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(proc_11_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(proc_11_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(proc_11_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(proc_11_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(proc_11_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(proc_11_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(proc_11_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(proc_11_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(proc_11_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(proc_11_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(proc_11_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(proc_11_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(proc_11_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(proc_11_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(proc_11_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(proc_11_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(proc_11_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(proc_11_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(proc_11_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(proc_11_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(proc_11_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(proc_11_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(proc_11_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(proc_11_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(proc_11_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(proc_11_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(proc_11_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(proc_11_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(proc_11_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(proc_11_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(proc_11_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(proc_11_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(proc_11_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(proc_11_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(proc_11_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(proc_11_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(proc_11_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(proc_11_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(proc_11_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(proc_11_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(proc_11_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(proc_11_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(proc_11_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(proc_11_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(proc_11_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(proc_11_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(proc_11_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(proc_11_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(proc_11_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(proc_11_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(proc_11_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(proc_11_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(proc_11_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(proc_11_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(proc_11_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(proc_11_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(proc_11_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(proc_11_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(proc_11_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(proc_11_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(proc_11_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(proc_11_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(proc_11_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(proc_11_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(proc_11_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(proc_11_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(proc_11_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(proc_11_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(proc_11_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(proc_11_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(proc_11_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(proc_11_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(proc_11_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_header_0(proc_11_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(proc_11_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(proc_11_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(proc_11_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(proc_11_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(proc_11_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(proc_11_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(proc_11_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(proc_11_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(proc_11_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(proc_11_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(proc_11_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(proc_11_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(proc_11_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(proc_11_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(proc_11_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(proc_11_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(proc_11_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(proc_11_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(proc_11_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(proc_11_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_valid(proc_11_io_pipe_phv_out_valid),
    .io_pipe_phv_out_last(proc_11_io_pipe_phv_out_last)
  );
  Processor proc_12 ( // @[ipsa.scala 56:25]
    .clock(proc_12_clock),
    .io_pipe_phv_in_data_0(proc_12_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(proc_12_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(proc_12_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(proc_12_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(proc_12_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(proc_12_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(proc_12_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(proc_12_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(proc_12_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(proc_12_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(proc_12_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(proc_12_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(proc_12_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(proc_12_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(proc_12_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(proc_12_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(proc_12_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(proc_12_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(proc_12_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(proc_12_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(proc_12_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(proc_12_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(proc_12_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(proc_12_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(proc_12_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(proc_12_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(proc_12_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(proc_12_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(proc_12_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(proc_12_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(proc_12_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(proc_12_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(proc_12_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(proc_12_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(proc_12_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(proc_12_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(proc_12_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(proc_12_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(proc_12_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(proc_12_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(proc_12_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(proc_12_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(proc_12_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(proc_12_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(proc_12_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(proc_12_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(proc_12_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(proc_12_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(proc_12_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(proc_12_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(proc_12_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(proc_12_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(proc_12_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(proc_12_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(proc_12_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(proc_12_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(proc_12_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(proc_12_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(proc_12_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(proc_12_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(proc_12_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(proc_12_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(proc_12_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(proc_12_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(proc_12_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(proc_12_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(proc_12_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(proc_12_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(proc_12_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(proc_12_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(proc_12_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(proc_12_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(proc_12_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(proc_12_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(proc_12_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(proc_12_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(proc_12_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(proc_12_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(proc_12_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(proc_12_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(proc_12_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(proc_12_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(proc_12_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(proc_12_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(proc_12_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(proc_12_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(proc_12_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(proc_12_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(proc_12_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(proc_12_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(proc_12_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(proc_12_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(proc_12_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(proc_12_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(proc_12_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(proc_12_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(proc_12_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(proc_12_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(proc_12_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(proc_12_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(proc_12_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(proc_12_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(proc_12_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(proc_12_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(proc_12_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(proc_12_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(proc_12_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(proc_12_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(proc_12_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(proc_12_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(proc_12_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(proc_12_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(proc_12_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(proc_12_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(proc_12_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(proc_12_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(proc_12_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(proc_12_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(proc_12_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(proc_12_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(proc_12_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(proc_12_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(proc_12_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(proc_12_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(proc_12_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(proc_12_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(proc_12_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(proc_12_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(proc_12_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(proc_12_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(proc_12_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(proc_12_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(proc_12_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(proc_12_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(proc_12_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(proc_12_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(proc_12_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(proc_12_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(proc_12_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(proc_12_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(proc_12_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(proc_12_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(proc_12_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(proc_12_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(proc_12_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(proc_12_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(proc_12_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(proc_12_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(proc_12_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(proc_12_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(proc_12_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(proc_12_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(proc_12_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(proc_12_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(proc_12_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(proc_12_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(proc_12_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(proc_12_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(proc_12_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(proc_12_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_header_0(proc_12_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(proc_12_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(proc_12_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(proc_12_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(proc_12_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(proc_12_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(proc_12_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(proc_12_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(proc_12_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(proc_12_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(proc_12_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(proc_12_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(proc_12_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(proc_12_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(proc_12_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(proc_12_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(proc_12_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(proc_12_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(proc_12_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(proc_12_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(proc_12_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(proc_12_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_in_valid(proc_12_io_pipe_phv_in_valid),
    .io_pipe_phv_in_last(proc_12_io_pipe_phv_in_last),
    .io_pipe_phv_out_data_0(proc_12_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(proc_12_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(proc_12_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(proc_12_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(proc_12_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(proc_12_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(proc_12_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(proc_12_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(proc_12_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(proc_12_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(proc_12_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(proc_12_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(proc_12_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(proc_12_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(proc_12_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(proc_12_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(proc_12_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(proc_12_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(proc_12_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(proc_12_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(proc_12_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(proc_12_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(proc_12_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(proc_12_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(proc_12_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(proc_12_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(proc_12_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(proc_12_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(proc_12_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(proc_12_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(proc_12_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(proc_12_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(proc_12_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(proc_12_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(proc_12_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(proc_12_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(proc_12_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(proc_12_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(proc_12_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(proc_12_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(proc_12_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(proc_12_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(proc_12_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(proc_12_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(proc_12_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(proc_12_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(proc_12_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(proc_12_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(proc_12_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(proc_12_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(proc_12_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(proc_12_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(proc_12_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(proc_12_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(proc_12_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(proc_12_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(proc_12_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(proc_12_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(proc_12_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(proc_12_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(proc_12_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(proc_12_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(proc_12_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(proc_12_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(proc_12_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(proc_12_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(proc_12_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(proc_12_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(proc_12_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(proc_12_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(proc_12_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(proc_12_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(proc_12_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(proc_12_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(proc_12_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(proc_12_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(proc_12_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(proc_12_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(proc_12_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(proc_12_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(proc_12_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(proc_12_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(proc_12_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(proc_12_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(proc_12_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(proc_12_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(proc_12_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(proc_12_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(proc_12_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(proc_12_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(proc_12_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(proc_12_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(proc_12_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(proc_12_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(proc_12_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(proc_12_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(proc_12_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(proc_12_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(proc_12_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(proc_12_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(proc_12_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(proc_12_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(proc_12_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(proc_12_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(proc_12_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(proc_12_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(proc_12_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(proc_12_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(proc_12_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(proc_12_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(proc_12_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(proc_12_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(proc_12_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(proc_12_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(proc_12_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(proc_12_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(proc_12_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(proc_12_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(proc_12_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(proc_12_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(proc_12_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(proc_12_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(proc_12_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(proc_12_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(proc_12_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(proc_12_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(proc_12_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(proc_12_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(proc_12_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(proc_12_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(proc_12_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(proc_12_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(proc_12_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(proc_12_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(proc_12_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(proc_12_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(proc_12_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(proc_12_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(proc_12_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(proc_12_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(proc_12_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(proc_12_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(proc_12_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(proc_12_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(proc_12_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(proc_12_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(proc_12_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(proc_12_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(proc_12_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(proc_12_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(proc_12_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(proc_12_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(proc_12_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(proc_12_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(proc_12_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(proc_12_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(proc_12_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(proc_12_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(proc_12_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(proc_12_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_header_0(proc_12_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(proc_12_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(proc_12_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(proc_12_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(proc_12_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(proc_12_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(proc_12_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(proc_12_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(proc_12_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(proc_12_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(proc_12_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(proc_12_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(proc_12_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(proc_12_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(proc_12_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(proc_12_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(proc_12_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(proc_12_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(proc_12_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(proc_12_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(proc_12_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_valid(proc_12_io_pipe_phv_out_valid),
    .io_pipe_phv_out_last(proc_12_io_pipe_phv_out_last)
  );
  Processor proc_13 ( // @[ipsa.scala 56:25]
    .clock(proc_13_clock),
    .io_pipe_phv_in_data_0(proc_13_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(proc_13_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(proc_13_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(proc_13_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(proc_13_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(proc_13_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(proc_13_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(proc_13_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(proc_13_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(proc_13_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(proc_13_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(proc_13_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(proc_13_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(proc_13_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(proc_13_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(proc_13_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(proc_13_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(proc_13_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(proc_13_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(proc_13_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(proc_13_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(proc_13_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(proc_13_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(proc_13_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(proc_13_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(proc_13_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(proc_13_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(proc_13_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(proc_13_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(proc_13_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(proc_13_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(proc_13_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(proc_13_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(proc_13_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(proc_13_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(proc_13_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(proc_13_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(proc_13_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(proc_13_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(proc_13_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(proc_13_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(proc_13_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(proc_13_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(proc_13_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(proc_13_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(proc_13_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(proc_13_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(proc_13_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(proc_13_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(proc_13_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(proc_13_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(proc_13_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(proc_13_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(proc_13_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(proc_13_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(proc_13_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(proc_13_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(proc_13_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(proc_13_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(proc_13_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(proc_13_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(proc_13_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(proc_13_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(proc_13_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(proc_13_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(proc_13_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(proc_13_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(proc_13_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(proc_13_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(proc_13_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(proc_13_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(proc_13_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(proc_13_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(proc_13_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(proc_13_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(proc_13_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(proc_13_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(proc_13_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(proc_13_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(proc_13_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(proc_13_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(proc_13_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(proc_13_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(proc_13_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(proc_13_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(proc_13_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(proc_13_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(proc_13_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(proc_13_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(proc_13_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(proc_13_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(proc_13_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(proc_13_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(proc_13_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(proc_13_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(proc_13_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(proc_13_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(proc_13_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(proc_13_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(proc_13_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(proc_13_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(proc_13_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(proc_13_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(proc_13_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(proc_13_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(proc_13_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(proc_13_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(proc_13_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(proc_13_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(proc_13_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(proc_13_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(proc_13_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(proc_13_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(proc_13_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(proc_13_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(proc_13_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(proc_13_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(proc_13_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(proc_13_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(proc_13_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(proc_13_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(proc_13_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(proc_13_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(proc_13_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(proc_13_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(proc_13_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(proc_13_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(proc_13_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(proc_13_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(proc_13_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(proc_13_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(proc_13_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(proc_13_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(proc_13_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(proc_13_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(proc_13_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(proc_13_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(proc_13_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(proc_13_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(proc_13_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(proc_13_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(proc_13_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(proc_13_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(proc_13_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(proc_13_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(proc_13_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(proc_13_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(proc_13_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(proc_13_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(proc_13_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(proc_13_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(proc_13_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(proc_13_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(proc_13_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(proc_13_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(proc_13_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(proc_13_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(proc_13_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(proc_13_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(proc_13_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_header_0(proc_13_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(proc_13_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(proc_13_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(proc_13_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(proc_13_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(proc_13_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(proc_13_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(proc_13_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(proc_13_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(proc_13_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(proc_13_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(proc_13_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(proc_13_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(proc_13_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(proc_13_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(proc_13_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(proc_13_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(proc_13_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(proc_13_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(proc_13_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(proc_13_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(proc_13_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_in_valid(proc_13_io_pipe_phv_in_valid),
    .io_pipe_phv_in_last(proc_13_io_pipe_phv_in_last),
    .io_pipe_phv_out_data_0(proc_13_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(proc_13_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(proc_13_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(proc_13_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(proc_13_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(proc_13_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(proc_13_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(proc_13_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(proc_13_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(proc_13_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(proc_13_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(proc_13_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(proc_13_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(proc_13_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(proc_13_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(proc_13_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(proc_13_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(proc_13_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(proc_13_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(proc_13_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(proc_13_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(proc_13_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(proc_13_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(proc_13_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(proc_13_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(proc_13_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(proc_13_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(proc_13_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(proc_13_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(proc_13_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(proc_13_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(proc_13_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(proc_13_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(proc_13_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(proc_13_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(proc_13_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(proc_13_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(proc_13_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(proc_13_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(proc_13_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(proc_13_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(proc_13_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(proc_13_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(proc_13_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(proc_13_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(proc_13_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(proc_13_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(proc_13_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(proc_13_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(proc_13_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(proc_13_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(proc_13_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(proc_13_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(proc_13_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(proc_13_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(proc_13_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(proc_13_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(proc_13_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(proc_13_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(proc_13_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(proc_13_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(proc_13_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(proc_13_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(proc_13_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(proc_13_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(proc_13_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(proc_13_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(proc_13_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(proc_13_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(proc_13_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(proc_13_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(proc_13_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(proc_13_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(proc_13_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(proc_13_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(proc_13_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(proc_13_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(proc_13_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(proc_13_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(proc_13_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(proc_13_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(proc_13_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(proc_13_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(proc_13_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(proc_13_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(proc_13_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(proc_13_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(proc_13_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(proc_13_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(proc_13_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(proc_13_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(proc_13_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(proc_13_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(proc_13_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(proc_13_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(proc_13_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(proc_13_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(proc_13_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(proc_13_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(proc_13_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(proc_13_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(proc_13_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(proc_13_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(proc_13_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(proc_13_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(proc_13_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(proc_13_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(proc_13_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(proc_13_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(proc_13_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(proc_13_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(proc_13_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(proc_13_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(proc_13_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(proc_13_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(proc_13_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(proc_13_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(proc_13_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(proc_13_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(proc_13_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(proc_13_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(proc_13_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(proc_13_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(proc_13_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(proc_13_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(proc_13_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(proc_13_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(proc_13_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(proc_13_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(proc_13_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(proc_13_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(proc_13_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(proc_13_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(proc_13_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(proc_13_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(proc_13_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(proc_13_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(proc_13_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(proc_13_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(proc_13_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(proc_13_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(proc_13_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(proc_13_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(proc_13_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(proc_13_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(proc_13_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(proc_13_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(proc_13_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(proc_13_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(proc_13_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(proc_13_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(proc_13_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(proc_13_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(proc_13_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(proc_13_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(proc_13_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(proc_13_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(proc_13_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(proc_13_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(proc_13_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_header_0(proc_13_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(proc_13_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(proc_13_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(proc_13_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(proc_13_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(proc_13_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(proc_13_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(proc_13_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(proc_13_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(proc_13_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(proc_13_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(proc_13_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(proc_13_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(proc_13_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(proc_13_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(proc_13_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(proc_13_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(proc_13_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(proc_13_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(proc_13_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(proc_13_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_valid(proc_13_io_pipe_phv_out_valid),
    .io_pipe_phv_out_last(proc_13_io_pipe_phv_out_last)
  );
  Processor proc_14 ( // @[ipsa.scala 56:25]
    .clock(proc_14_clock),
    .io_pipe_phv_in_data_0(proc_14_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(proc_14_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(proc_14_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(proc_14_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(proc_14_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(proc_14_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(proc_14_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(proc_14_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(proc_14_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(proc_14_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(proc_14_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(proc_14_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(proc_14_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(proc_14_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(proc_14_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(proc_14_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(proc_14_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(proc_14_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(proc_14_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(proc_14_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(proc_14_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(proc_14_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(proc_14_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(proc_14_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(proc_14_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(proc_14_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(proc_14_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(proc_14_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(proc_14_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(proc_14_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(proc_14_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(proc_14_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(proc_14_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(proc_14_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(proc_14_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(proc_14_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(proc_14_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(proc_14_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(proc_14_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(proc_14_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(proc_14_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(proc_14_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(proc_14_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(proc_14_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(proc_14_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(proc_14_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(proc_14_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(proc_14_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(proc_14_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(proc_14_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(proc_14_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(proc_14_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(proc_14_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(proc_14_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(proc_14_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(proc_14_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(proc_14_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(proc_14_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(proc_14_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(proc_14_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(proc_14_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(proc_14_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(proc_14_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(proc_14_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(proc_14_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(proc_14_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(proc_14_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(proc_14_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(proc_14_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(proc_14_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(proc_14_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(proc_14_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(proc_14_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(proc_14_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(proc_14_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(proc_14_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(proc_14_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(proc_14_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(proc_14_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(proc_14_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(proc_14_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(proc_14_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(proc_14_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(proc_14_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(proc_14_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(proc_14_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(proc_14_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(proc_14_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(proc_14_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(proc_14_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(proc_14_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(proc_14_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(proc_14_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(proc_14_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(proc_14_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(proc_14_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(proc_14_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(proc_14_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(proc_14_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(proc_14_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(proc_14_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(proc_14_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(proc_14_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(proc_14_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(proc_14_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(proc_14_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(proc_14_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(proc_14_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(proc_14_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(proc_14_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(proc_14_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(proc_14_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(proc_14_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(proc_14_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(proc_14_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(proc_14_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(proc_14_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(proc_14_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(proc_14_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(proc_14_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(proc_14_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(proc_14_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(proc_14_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(proc_14_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(proc_14_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(proc_14_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(proc_14_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(proc_14_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(proc_14_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(proc_14_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(proc_14_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(proc_14_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(proc_14_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(proc_14_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(proc_14_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(proc_14_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(proc_14_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(proc_14_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(proc_14_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(proc_14_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(proc_14_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(proc_14_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(proc_14_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(proc_14_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(proc_14_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(proc_14_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(proc_14_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(proc_14_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(proc_14_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(proc_14_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(proc_14_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(proc_14_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(proc_14_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(proc_14_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(proc_14_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(proc_14_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(proc_14_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(proc_14_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(proc_14_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(proc_14_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_header_0(proc_14_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(proc_14_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(proc_14_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(proc_14_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(proc_14_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(proc_14_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(proc_14_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(proc_14_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(proc_14_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(proc_14_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(proc_14_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(proc_14_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(proc_14_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(proc_14_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(proc_14_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(proc_14_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(proc_14_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(proc_14_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(proc_14_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(proc_14_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(proc_14_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(proc_14_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_in_valid(proc_14_io_pipe_phv_in_valid),
    .io_pipe_phv_in_last(proc_14_io_pipe_phv_in_last),
    .io_pipe_phv_out_data_0(proc_14_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(proc_14_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(proc_14_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(proc_14_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(proc_14_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(proc_14_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(proc_14_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(proc_14_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(proc_14_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(proc_14_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(proc_14_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(proc_14_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(proc_14_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(proc_14_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(proc_14_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(proc_14_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(proc_14_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(proc_14_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(proc_14_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(proc_14_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(proc_14_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(proc_14_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(proc_14_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(proc_14_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(proc_14_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(proc_14_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(proc_14_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(proc_14_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(proc_14_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(proc_14_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(proc_14_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(proc_14_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(proc_14_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(proc_14_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(proc_14_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(proc_14_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(proc_14_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(proc_14_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(proc_14_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(proc_14_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(proc_14_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(proc_14_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(proc_14_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(proc_14_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(proc_14_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(proc_14_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(proc_14_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(proc_14_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(proc_14_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(proc_14_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(proc_14_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(proc_14_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(proc_14_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(proc_14_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(proc_14_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(proc_14_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(proc_14_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(proc_14_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(proc_14_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(proc_14_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(proc_14_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(proc_14_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(proc_14_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(proc_14_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(proc_14_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(proc_14_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(proc_14_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(proc_14_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(proc_14_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(proc_14_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(proc_14_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(proc_14_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(proc_14_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(proc_14_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(proc_14_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(proc_14_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(proc_14_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(proc_14_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(proc_14_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(proc_14_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(proc_14_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(proc_14_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(proc_14_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(proc_14_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(proc_14_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(proc_14_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(proc_14_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(proc_14_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(proc_14_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(proc_14_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(proc_14_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(proc_14_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(proc_14_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(proc_14_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(proc_14_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(proc_14_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(proc_14_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(proc_14_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(proc_14_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(proc_14_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(proc_14_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(proc_14_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(proc_14_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(proc_14_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(proc_14_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(proc_14_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(proc_14_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(proc_14_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(proc_14_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(proc_14_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(proc_14_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(proc_14_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(proc_14_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(proc_14_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(proc_14_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(proc_14_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(proc_14_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(proc_14_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(proc_14_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(proc_14_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(proc_14_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(proc_14_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(proc_14_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(proc_14_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(proc_14_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(proc_14_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(proc_14_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(proc_14_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(proc_14_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(proc_14_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(proc_14_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(proc_14_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(proc_14_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(proc_14_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(proc_14_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(proc_14_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(proc_14_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(proc_14_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(proc_14_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(proc_14_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(proc_14_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(proc_14_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(proc_14_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(proc_14_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(proc_14_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(proc_14_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(proc_14_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(proc_14_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(proc_14_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(proc_14_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(proc_14_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(proc_14_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(proc_14_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(proc_14_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(proc_14_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(proc_14_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(proc_14_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(proc_14_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(proc_14_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(proc_14_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_header_0(proc_14_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(proc_14_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(proc_14_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(proc_14_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(proc_14_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(proc_14_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(proc_14_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(proc_14_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(proc_14_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(proc_14_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(proc_14_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(proc_14_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(proc_14_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(proc_14_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(proc_14_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(proc_14_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(proc_14_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(proc_14_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(proc_14_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(proc_14_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(proc_14_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_valid(proc_14_io_pipe_phv_out_valid),
    .io_pipe_phv_out_last(proc_14_io_pipe_phv_out_last)
  );
  Processor proc_15 ( // @[ipsa.scala 56:25]
    .clock(proc_15_clock),
    .io_pipe_phv_in_data_0(proc_15_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(proc_15_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(proc_15_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(proc_15_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(proc_15_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(proc_15_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(proc_15_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(proc_15_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(proc_15_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(proc_15_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(proc_15_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(proc_15_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(proc_15_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(proc_15_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(proc_15_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(proc_15_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(proc_15_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(proc_15_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(proc_15_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(proc_15_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(proc_15_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(proc_15_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(proc_15_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(proc_15_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(proc_15_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(proc_15_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(proc_15_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(proc_15_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(proc_15_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(proc_15_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(proc_15_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(proc_15_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(proc_15_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(proc_15_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(proc_15_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(proc_15_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(proc_15_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(proc_15_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(proc_15_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(proc_15_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(proc_15_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(proc_15_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(proc_15_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(proc_15_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(proc_15_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(proc_15_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(proc_15_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(proc_15_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(proc_15_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(proc_15_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(proc_15_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(proc_15_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(proc_15_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(proc_15_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(proc_15_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(proc_15_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(proc_15_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(proc_15_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(proc_15_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(proc_15_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(proc_15_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(proc_15_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(proc_15_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(proc_15_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(proc_15_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(proc_15_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(proc_15_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(proc_15_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(proc_15_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(proc_15_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(proc_15_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(proc_15_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(proc_15_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(proc_15_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(proc_15_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(proc_15_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(proc_15_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(proc_15_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(proc_15_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(proc_15_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(proc_15_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(proc_15_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(proc_15_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(proc_15_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(proc_15_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(proc_15_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(proc_15_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(proc_15_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(proc_15_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(proc_15_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(proc_15_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(proc_15_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(proc_15_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(proc_15_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(proc_15_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(proc_15_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(proc_15_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(proc_15_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(proc_15_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(proc_15_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(proc_15_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(proc_15_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(proc_15_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(proc_15_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(proc_15_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(proc_15_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(proc_15_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(proc_15_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(proc_15_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(proc_15_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(proc_15_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(proc_15_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(proc_15_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(proc_15_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(proc_15_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(proc_15_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(proc_15_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(proc_15_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(proc_15_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(proc_15_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(proc_15_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(proc_15_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(proc_15_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(proc_15_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(proc_15_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(proc_15_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(proc_15_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(proc_15_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(proc_15_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(proc_15_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(proc_15_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(proc_15_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(proc_15_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(proc_15_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(proc_15_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(proc_15_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(proc_15_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(proc_15_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(proc_15_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(proc_15_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(proc_15_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(proc_15_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(proc_15_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(proc_15_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(proc_15_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(proc_15_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(proc_15_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(proc_15_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(proc_15_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(proc_15_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(proc_15_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(proc_15_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(proc_15_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(proc_15_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(proc_15_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(proc_15_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(proc_15_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(proc_15_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(proc_15_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(proc_15_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_header_0(proc_15_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(proc_15_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(proc_15_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(proc_15_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(proc_15_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(proc_15_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(proc_15_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(proc_15_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(proc_15_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(proc_15_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(proc_15_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(proc_15_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(proc_15_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(proc_15_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(proc_15_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(proc_15_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(proc_15_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(proc_15_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(proc_15_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(proc_15_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(proc_15_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(proc_15_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_in_valid(proc_15_io_pipe_phv_in_valid),
    .io_pipe_phv_in_last(proc_15_io_pipe_phv_in_last),
    .io_pipe_phv_out_data_0(proc_15_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(proc_15_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(proc_15_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(proc_15_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(proc_15_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(proc_15_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(proc_15_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(proc_15_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(proc_15_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(proc_15_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(proc_15_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(proc_15_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(proc_15_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(proc_15_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(proc_15_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(proc_15_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(proc_15_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(proc_15_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(proc_15_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(proc_15_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(proc_15_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(proc_15_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(proc_15_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(proc_15_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(proc_15_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(proc_15_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(proc_15_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(proc_15_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(proc_15_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(proc_15_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(proc_15_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(proc_15_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(proc_15_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(proc_15_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(proc_15_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(proc_15_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(proc_15_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(proc_15_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(proc_15_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(proc_15_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(proc_15_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(proc_15_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(proc_15_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(proc_15_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(proc_15_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(proc_15_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(proc_15_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(proc_15_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(proc_15_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(proc_15_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(proc_15_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(proc_15_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(proc_15_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(proc_15_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(proc_15_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(proc_15_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(proc_15_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(proc_15_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(proc_15_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(proc_15_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(proc_15_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(proc_15_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(proc_15_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(proc_15_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(proc_15_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(proc_15_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(proc_15_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(proc_15_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(proc_15_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(proc_15_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(proc_15_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(proc_15_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(proc_15_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(proc_15_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(proc_15_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(proc_15_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(proc_15_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(proc_15_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(proc_15_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(proc_15_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(proc_15_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(proc_15_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(proc_15_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(proc_15_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(proc_15_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(proc_15_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(proc_15_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(proc_15_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(proc_15_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(proc_15_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(proc_15_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(proc_15_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(proc_15_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(proc_15_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(proc_15_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(proc_15_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(proc_15_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(proc_15_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(proc_15_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(proc_15_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(proc_15_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(proc_15_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(proc_15_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(proc_15_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(proc_15_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(proc_15_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(proc_15_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(proc_15_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(proc_15_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(proc_15_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(proc_15_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(proc_15_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(proc_15_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(proc_15_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(proc_15_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(proc_15_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(proc_15_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(proc_15_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(proc_15_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(proc_15_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(proc_15_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(proc_15_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(proc_15_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(proc_15_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(proc_15_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(proc_15_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(proc_15_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(proc_15_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(proc_15_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(proc_15_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(proc_15_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(proc_15_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(proc_15_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(proc_15_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(proc_15_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(proc_15_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(proc_15_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(proc_15_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(proc_15_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(proc_15_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(proc_15_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(proc_15_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(proc_15_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(proc_15_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(proc_15_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(proc_15_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(proc_15_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(proc_15_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(proc_15_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(proc_15_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(proc_15_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(proc_15_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(proc_15_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(proc_15_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(proc_15_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(proc_15_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(proc_15_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(proc_15_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(proc_15_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(proc_15_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_header_0(proc_15_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(proc_15_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(proc_15_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(proc_15_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(proc_15_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(proc_15_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(proc_15_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(proc_15_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(proc_15_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(proc_15_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(proc_15_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(proc_15_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(proc_15_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(proc_15_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(proc_15_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(proc_15_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(proc_15_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(proc_15_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(proc_15_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(proc_15_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(proc_15_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_valid(proc_15_io_pipe_phv_out_valid),
    .io_pipe_phv_out_last(proc_15_io_pipe_phv_out_last)
  );
  SRAMCluster sram_cluster_0 ( // @[ipsa.scala 62:25]
    .clock(sram_cluster_0_clock)
  );
  SRAMCluster sram_cluster_1 ( // @[ipsa.scala 62:25]
    .clock(sram_cluster_1_clock)
  );
  SRAMCluster sram_cluster_2 ( // @[ipsa.scala 62:25]
    .clock(sram_cluster_2_clock)
  );
  SRAMCluster sram_cluster_3 ( // @[ipsa.scala 62:25]
    .clock(sram_cluster_3_clock)
  );
  SRAMCluster sram_cluster_4 ( // @[ipsa.scala 62:25]
    .clock(sram_cluster_4_clock)
  );
  SRAMCluster sram_cluster_5 ( // @[ipsa.scala 62:25]
    .clock(sram_cluster_5_clock)
  );
  SRAMCluster sram_cluster_6 ( // @[ipsa.scala 62:25]
    .clock(sram_cluster_6_clock)
  );
  SRAMCluster sram_cluster_7 ( // @[ipsa.scala 62:25]
    .clock(sram_cluster_7_clock)
  );
  Initializer init ( // @[ipsa.scala 74:22]
    .clock(init_clock),
    .io_pipe_phv_in_data_0(init_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(init_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(init_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(init_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(init_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(init_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(init_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(init_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(init_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(init_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(init_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(init_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(init_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(init_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(init_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(init_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(init_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(init_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(init_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(init_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(init_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(init_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(init_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(init_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(init_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(init_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(init_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(init_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(init_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(init_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(init_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(init_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(init_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(init_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(init_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(init_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(init_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(init_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(init_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(init_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(init_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(init_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(init_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(init_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(init_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(init_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(init_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(init_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(init_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(init_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(init_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(init_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(init_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(init_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(init_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(init_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(init_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(init_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(init_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(init_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(init_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(init_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(init_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(init_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(init_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(init_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(init_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(init_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(init_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(init_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(init_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(init_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(init_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(init_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(init_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(init_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(init_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(init_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(init_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(init_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(init_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(init_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(init_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(init_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(init_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(init_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(init_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(init_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(init_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(init_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(init_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(init_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(init_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(init_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(init_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(init_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(init_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(init_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(init_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(init_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(init_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(init_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(init_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(init_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(init_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(init_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(init_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(init_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(init_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(init_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(init_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(init_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(init_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(init_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(init_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(init_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(init_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(init_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(init_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(init_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(init_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(init_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(init_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(init_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(init_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(init_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(init_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(init_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_valid(init_io_pipe_phv_in_valid),
    .io_pipe_phv_in_last(init_io_pipe_phv_in_last),
    .io_pipe_phv_out_data_0(init_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(init_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(init_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(init_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(init_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(init_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(init_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(init_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(init_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(init_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(init_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(init_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(init_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(init_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(init_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(init_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(init_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(init_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(init_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(init_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(init_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(init_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(init_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(init_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(init_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(init_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(init_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(init_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(init_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(init_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(init_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(init_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(init_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(init_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(init_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(init_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(init_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(init_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(init_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(init_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(init_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(init_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(init_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(init_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(init_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(init_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(init_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(init_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(init_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(init_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(init_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(init_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(init_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(init_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(init_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(init_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(init_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(init_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(init_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(init_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(init_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(init_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(init_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(init_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(init_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(init_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(init_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(init_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(init_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(init_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(init_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(init_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(init_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(init_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(init_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(init_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(init_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(init_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(init_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(init_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(init_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(init_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(init_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(init_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(init_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(init_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(init_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(init_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(init_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(init_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(init_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(init_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(init_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(init_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(init_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(init_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(init_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(init_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(init_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(init_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(init_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(init_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(init_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(init_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(init_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(init_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(init_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(init_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(init_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(init_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(init_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(init_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(init_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(init_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(init_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(init_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(init_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(init_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(init_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(init_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(init_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(init_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(init_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(init_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(init_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(init_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(init_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(init_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_valid(init_io_pipe_phv_out_valid),
    .io_pipe_phv_out_last(init_io_pipe_phv_out_last)
  );
  InterProcessorTransfer trans_0 ( // @[ipsa.scala 79:25]
    .clock(trans_0_clock),
    .io_pipe_phv_in_data_0(trans_0_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(trans_0_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(trans_0_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(trans_0_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(trans_0_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(trans_0_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(trans_0_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(trans_0_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(trans_0_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(trans_0_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(trans_0_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(trans_0_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(trans_0_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(trans_0_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(trans_0_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(trans_0_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(trans_0_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(trans_0_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(trans_0_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(trans_0_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(trans_0_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(trans_0_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(trans_0_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(trans_0_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(trans_0_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(trans_0_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(trans_0_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(trans_0_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(trans_0_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(trans_0_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(trans_0_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(trans_0_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(trans_0_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(trans_0_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(trans_0_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(trans_0_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(trans_0_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(trans_0_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(trans_0_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(trans_0_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(trans_0_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(trans_0_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(trans_0_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(trans_0_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(trans_0_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(trans_0_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(trans_0_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(trans_0_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(trans_0_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(trans_0_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(trans_0_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(trans_0_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(trans_0_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(trans_0_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(trans_0_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(trans_0_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(trans_0_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(trans_0_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(trans_0_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(trans_0_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(trans_0_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(trans_0_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(trans_0_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(trans_0_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(trans_0_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(trans_0_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(trans_0_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(trans_0_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(trans_0_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(trans_0_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(trans_0_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(trans_0_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(trans_0_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(trans_0_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(trans_0_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(trans_0_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(trans_0_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(trans_0_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(trans_0_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(trans_0_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(trans_0_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(trans_0_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(trans_0_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(trans_0_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(trans_0_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(trans_0_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(trans_0_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(trans_0_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(trans_0_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(trans_0_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(trans_0_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(trans_0_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(trans_0_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(trans_0_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(trans_0_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(trans_0_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(trans_0_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(trans_0_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(trans_0_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(trans_0_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(trans_0_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(trans_0_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(trans_0_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(trans_0_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(trans_0_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(trans_0_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(trans_0_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(trans_0_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(trans_0_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(trans_0_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(trans_0_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(trans_0_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(trans_0_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(trans_0_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(trans_0_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(trans_0_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(trans_0_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(trans_0_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(trans_0_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(trans_0_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(trans_0_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(trans_0_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(trans_0_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(trans_0_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(trans_0_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(trans_0_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(trans_0_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(trans_0_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(trans_0_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(trans_0_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(trans_0_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(trans_0_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(trans_0_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(trans_0_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(trans_0_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(trans_0_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(trans_0_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(trans_0_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(trans_0_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(trans_0_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(trans_0_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(trans_0_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(trans_0_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(trans_0_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(trans_0_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(trans_0_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(trans_0_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(trans_0_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(trans_0_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(trans_0_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(trans_0_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(trans_0_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(trans_0_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(trans_0_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(trans_0_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(trans_0_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(trans_0_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(trans_0_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(trans_0_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(trans_0_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_header_0(trans_0_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(trans_0_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(trans_0_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(trans_0_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(trans_0_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(trans_0_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(trans_0_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(trans_0_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(trans_0_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(trans_0_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(trans_0_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(trans_0_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(trans_0_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(trans_0_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(trans_0_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(trans_0_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(trans_0_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(trans_0_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(trans_0_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(trans_0_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(trans_0_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_valid(trans_0_io_pipe_phv_in_valid),
    .io_pipe_phv_in_last(trans_0_io_pipe_phv_in_last),
    .io_pipe_phv_out_data_0(trans_0_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(trans_0_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(trans_0_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(trans_0_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(trans_0_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(trans_0_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(trans_0_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(trans_0_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(trans_0_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(trans_0_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(trans_0_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(trans_0_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(trans_0_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(trans_0_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(trans_0_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(trans_0_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(trans_0_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(trans_0_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(trans_0_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(trans_0_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(trans_0_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(trans_0_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(trans_0_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(trans_0_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(trans_0_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(trans_0_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(trans_0_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(trans_0_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(trans_0_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(trans_0_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(trans_0_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(trans_0_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(trans_0_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(trans_0_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(trans_0_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(trans_0_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(trans_0_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(trans_0_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(trans_0_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(trans_0_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(trans_0_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(trans_0_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(trans_0_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(trans_0_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(trans_0_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(trans_0_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(trans_0_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(trans_0_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(trans_0_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(trans_0_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(trans_0_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(trans_0_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(trans_0_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(trans_0_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(trans_0_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(trans_0_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(trans_0_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(trans_0_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(trans_0_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(trans_0_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(trans_0_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(trans_0_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(trans_0_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(trans_0_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(trans_0_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(trans_0_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(trans_0_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(trans_0_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(trans_0_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(trans_0_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(trans_0_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(trans_0_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(trans_0_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(trans_0_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(trans_0_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(trans_0_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(trans_0_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(trans_0_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(trans_0_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(trans_0_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(trans_0_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(trans_0_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(trans_0_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(trans_0_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(trans_0_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(trans_0_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(trans_0_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(trans_0_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(trans_0_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(trans_0_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(trans_0_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(trans_0_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(trans_0_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(trans_0_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(trans_0_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(trans_0_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(trans_0_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(trans_0_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(trans_0_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(trans_0_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(trans_0_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(trans_0_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(trans_0_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(trans_0_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(trans_0_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(trans_0_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(trans_0_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(trans_0_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(trans_0_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(trans_0_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(trans_0_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(trans_0_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(trans_0_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(trans_0_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(trans_0_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(trans_0_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(trans_0_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(trans_0_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(trans_0_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(trans_0_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(trans_0_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(trans_0_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(trans_0_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(trans_0_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(trans_0_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(trans_0_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(trans_0_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(trans_0_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(trans_0_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(trans_0_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(trans_0_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(trans_0_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(trans_0_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(trans_0_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(trans_0_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(trans_0_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(trans_0_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(trans_0_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(trans_0_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(trans_0_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(trans_0_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(trans_0_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(trans_0_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(trans_0_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(trans_0_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(trans_0_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(trans_0_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(trans_0_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(trans_0_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(trans_0_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(trans_0_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(trans_0_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(trans_0_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(trans_0_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(trans_0_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(trans_0_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(trans_0_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(trans_0_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(trans_0_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(trans_0_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_header_0(trans_0_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(trans_0_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(trans_0_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(trans_0_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(trans_0_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(trans_0_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(trans_0_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(trans_0_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(trans_0_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(trans_0_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(trans_0_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(trans_0_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(trans_0_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(trans_0_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(trans_0_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(trans_0_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(trans_0_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(trans_0_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(trans_0_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(trans_0_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(trans_0_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(trans_0_io_pipe_phv_out_is_valid_processor),
    .io_pipe_phv_out_valid(trans_0_io_pipe_phv_out_valid),
    .io_pipe_phv_out_last(trans_0_io_pipe_phv_out_last),
    .io_next_proc_exist(trans_0_io_next_proc_exist)
  );
  InterProcessorTransfer trans_1 ( // @[ipsa.scala 79:25]
    .clock(trans_1_clock),
    .io_pipe_phv_in_data_0(trans_1_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(trans_1_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(trans_1_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(trans_1_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(trans_1_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(trans_1_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(trans_1_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(trans_1_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(trans_1_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(trans_1_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(trans_1_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(trans_1_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(trans_1_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(trans_1_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(trans_1_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(trans_1_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(trans_1_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(trans_1_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(trans_1_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(trans_1_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(trans_1_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(trans_1_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(trans_1_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(trans_1_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(trans_1_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(trans_1_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(trans_1_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(trans_1_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(trans_1_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(trans_1_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(trans_1_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(trans_1_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(trans_1_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(trans_1_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(trans_1_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(trans_1_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(trans_1_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(trans_1_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(trans_1_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(trans_1_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(trans_1_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(trans_1_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(trans_1_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(trans_1_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(trans_1_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(trans_1_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(trans_1_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(trans_1_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(trans_1_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(trans_1_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(trans_1_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(trans_1_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(trans_1_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(trans_1_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(trans_1_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(trans_1_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(trans_1_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(trans_1_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(trans_1_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(trans_1_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(trans_1_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(trans_1_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(trans_1_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(trans_1_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(trans_1_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(trans_1_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(trans_1_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(trans_1_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(trans_1_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(trans_1_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(trans_1_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(trans_1_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(trans_1_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(trans_1_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(trans_1_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(trans_1_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(trans_1_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(trans_1_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(trans_1_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(trans_1_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(trans_1_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(trans_1_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(trans_1_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(trans_1_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(trans_1_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(trans_1_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(trans_1_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(trans_1_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(trans_1_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(trans_1_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(trans_1_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(trans_1_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(trans_1_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(trans_1_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(trans_1_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(trans_1_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(trans_1_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(trans_1_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(trans_1_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(trans_1_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(trans_1_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(trans_1_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(trans_1_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(trans_1_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(trans_1_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(trans_1_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(trans_1_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(trans_1_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(trans_1_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(trans_1_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(trans_1_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(trans_1_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(trans_1_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(trans_1_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(trans_1_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(trans_1_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(trans_1_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(trans_1_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(trans_1_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(trans_1_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(trans_1_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(trans_1_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(trans_1_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(trans_1_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(trans_1_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(trans_1_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(trans_1_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(trans_1_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(trans_1_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(trans_1_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(trans_1_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(trans_1_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(trans_1_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(trans_1_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(trans_1_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(trans_1_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(trans_1_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(trans_1_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(trans_1_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(trans_1_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(trans_1_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(trans_1_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(trans_1_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(trans_1_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(trans_1_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(trans_1_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(trans_1_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(trans_1_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(trans_1_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(trans_1_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(trans_1_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(trans_1_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(trans_1_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(trans_1_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(trans_1_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(trans_1_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(trans_1_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(trans_1_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(trans_1_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(trans_1_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_header_0(trans_1_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(trans_1_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(trans_1_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(trans_1_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(trans_1_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(trans_1_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(trans_1_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(trans_1_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(trans_1_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(trans_1_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(trans_1_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(trans_1_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(trans_1_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(trans_1_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(trans_1_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(trans_1_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(trans_1_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(trans_1_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(trans_1_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(trans_1_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(trans_1_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_valid(trans_1_io_pipe_phv_in_valid),
    .io_pipe_phv_in_last(trans_1_io_pipe_phv_in_last),
    .io_pipe_phv_out_data_0(trans_1_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(trans_1_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(trans_1_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(trans_1_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(trans_1_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(trans_1_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(trans_1_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(trans_1_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(trans_1_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(trans_1_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(trans_1_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(trans_1_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(trans_1_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(trans_1_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(trans_1_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(trans_1_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(trans_1_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(trans_1_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(trans_1_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(trans_1_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(trans_1_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(trans_1_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(trans_1_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(trans_1_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(trans_1_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(trans_1_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(trans_1_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(trans_1_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(trans_1_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(trans_1_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(trans_1_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(trans_1_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(trans_1_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(trans_1_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(trans_1_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(trans_1_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(trans_1_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(trans_1_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(trans_1_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(trans_1_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(trans_1_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(trans_1_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(trans_1_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(trans_1_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(trans_1_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(trans_1_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(trans_1_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(trans_1_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(trans_1_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(trans_1_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(trans_1_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(trans_1_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(trans_1_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(trans_1_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(trans_1_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(trans_1_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(trans_1_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(trans_1_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(trans_1_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(trans_1_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(trans_1_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(trans_1_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(trans_1_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(trans_1_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(trans_1_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(trans_1_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(trans_1_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(trans_1_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(trans_1_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(trans_1_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(trans_1_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(trans_1_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(trans_1_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(trans_1_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(trans_1_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(trans_1_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(trans_1_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(trans_1_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(trans_1_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(trans_1_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(trans_1_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(trans_1_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(trans_1_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(trans_1_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(trans_1_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(trans_1_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(trans_1_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(trans_1_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(trans_1_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(trans_1_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(trans_1_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(trans_1_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(trans_1_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(trans_1_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(trans_1_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(trans_1_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(trans_1_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(trans_1_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(trans_1_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(trans_1_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(trans_1_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(trans_1_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(trans_1_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(trans_1_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(trans_1_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(trans_1_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(trans_1_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(trans_1_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(trans_1_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(trans_1_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(trans_1_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(trans_1_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(trans_1_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(trans_1_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(trans_1_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(trans_1_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(trans_1_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(trans_1_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(trans_1_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(trans_1_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(trans_1_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(trans_1_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(trans_1_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(trans_1_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(trans_1_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(trans_1_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(trans_1_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(trans_1_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(trans_1_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(trans_1_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(trans_1_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(trans_1_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(trans_1_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(trans_1_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(trans_1_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(trans_1_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(trans_1_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(trans_1_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(trans_1_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(trans_1_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(trans_1_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(trans_1_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(trans_1_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(trans_1_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(trans_1_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(trans_1_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(trans_1_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(trans_1_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(trans_1_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(trans_1_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(trans_1_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(trans_1_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(trans_1_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(trans_1_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(trans_1_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(trans_1_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(trans_1_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(trans_1_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(trans_1_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(trans_1_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_header_0(trans_1_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(trans_1_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(trans_1_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(trans_1_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(trans_1_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(trans_1_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(trans_1_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(trans_1_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(trans_1_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(trans_1_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(trans_1_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(trans_1_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(trans_1_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(trans_1_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(trans_1_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(trans_1_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(trans_1_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(trans_1_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(trans_1_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(trans_1_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(trans_1_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(trans_1_io_pipe_phv_out_is_valid_processor),
    .io_pipe_phv_out_valid(trans_1_io_pipe_phv_out_valid),
    .io_pipe_phv_out_last(trans_1_io_pipe_phv_out_last),
    .io_next_proc_exist(trans_1_io_next_proc_exist)
  );
  InterProcessorTransfer trans_2 ( // @[ipsa.scala 79:25]
    .clock(trans_2_clock),
    .io_pipe_phv_in_data_0(trans_2_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(trans_2_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(trans_2_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(trans_2_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(trans_2_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(trans_2_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(trans_2_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(trans_2_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(trans_2_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(trans_2_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(trans_2_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(trans_2_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(trans_2_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(trans_2_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(trans_2_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(trans_2_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(trans_2_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(trans_2_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(trans_2_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(trans_2_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(trans_2_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(trans_2_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(trans_2_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(trans_2_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(trans_2_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(trans_2_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(trans_2_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(trans_2_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(trans_2_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(trans_2_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(trans_2_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(trans_2_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(trans_2_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(trans_2_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(trans_2_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(trans_2_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(trans_2_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(trans_2_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(trans_2_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(trans_2_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(trans_2_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(trans_2_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(trans_2_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(trans_2_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(trans_2_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(trans_2_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(trans_2_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(trans_2_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(trans_2_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(trans_2_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(trans_2_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(trans_2_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(trans_2_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(trans_2_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(trans_2_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(trans_2_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(trans_2_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(trans_2_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(trans_2_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(trans_2_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(trans_2_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(trans_2_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(trans_2_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(trans_2_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(trans_2_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(trans_2_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(trans_2_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(trans_2_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(trans_2_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(trans_2_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(trans_2_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(trans_2_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(trans_2_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(trans_2_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(trans_2_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(trans_2_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(trans_2_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(trans_2_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(trans_2_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(trans_2_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(trans_2_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(trans_2_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(trans_2_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(trans_2_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(trans_2_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(trans_2_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(trans_2_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(trans_2_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(trans_2_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(trans_2_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(trans_2_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(trans_2_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(trans_2_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(trans_2_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(trans_2_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(trans_2_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(trans_2_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(trans_2_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(trans_2_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(trans_2_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(trans_2_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(trans_2_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(trans_2_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(trans_2_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(trans_2_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(trans_2_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(trans_2_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(trans_2_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(trans_2_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(trans_2_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(trans_2_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(trans_2_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(trans_2_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(trans_2_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(trans_2_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(trans_2_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(trans_2_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(trans_2_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(trans_2_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(trans_2_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(trans_2_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(trans_2_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(trans_2_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(trans_2_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(trans_2_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(trans_2_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(trans_2_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(trans_2_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(trans_2_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(trans_2_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(trans_2_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(trans_2_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(trans_2_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(trans_2_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(trans_2_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(trans_2_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(trans_2_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(trans_2_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(trans_2_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(trans_2_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(trans_2_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(trans_2_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(trans_2_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(trans_2_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(trans_2_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(trans_2_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(trans_2_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(trans_2_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(trans_2_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(trans_2_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(trans_2_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(trans_2_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(trans_2_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(trans_2_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(trans_2_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(trans_2_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(trans_2_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(trans_2_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(trans_2_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(trans_2_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_header_0(trans_2_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(trans_2_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(trans_2_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(trans_2_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(trans_2_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(trans_2_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(trans_2_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(trans_2_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(trans_2_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(trans_2_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(trans_2_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(trans_2_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(trans_2_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(trans_2_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(trans_2_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(trans_2_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(trans_2_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(trans_2_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(trans_2_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(trans_2_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(trans_2_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_valid(trans_2_io_pipe_phv_in_valid),
    .io_pipe_phv_in_last(trans_2_io_pipe_phv_in_last),
    .io_pipe_phv_out_data_0(trans_2_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(trans_2_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(trans_2_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(trans_2_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(trans_2_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(trans_2_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(trans_2_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(trans_2_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(trans_2_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(trans_2_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(trans_2_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(trans_2_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(trans_2_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(trans_2_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(trans_2_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(trans_2_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(trans_2_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(trans_2_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(trans_2_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(trans_2_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(trans_2_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(trans_2_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(trans_2_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(trans_2_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(trans_2_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(trans_2_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(trans_2_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(trans_2_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(trans_2_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(trans_2_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(trans_2_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(trans_2_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(trans_2_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(trans_2_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(trans_2_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(trans_2_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(trans_2_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(trans_2_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(trans_2_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(trans_2_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(trans_2_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(trans_2_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(trans_2_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(trans_2_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(trans_2_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(trans_2_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(trans_2_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(trans_2_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(trans_2_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(trans_2_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(trans_2_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(trans_2_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(trans_2_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(trans_2_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(trans_2_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(trans_2_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(trans_2_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(trans_2_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(trans_2_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(trans_2_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(trans_2_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(trans_2_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(trans_2_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(trans_2_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(trans_2_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(trans_2_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(trans_2_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(trans_2_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(trans_2_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(trans_2_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(trans_2_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(trans_2_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(trans_2_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(trans_2_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(trans_2_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(trans_2_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(trans_2_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(trans_2_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(trans_2_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(trans_2_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(trans_2_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(trans_2_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(trans_2_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(trans_2_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(trans_2_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(trans_2_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(trans_2_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(trans_2_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(trans_2_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(trans_2_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(trans_2_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(trans_2_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(trans_2_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(trans_2_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(trans_2_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(trans_2_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(trans_2_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(trans_2_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(trans_2_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(trans_2_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(trans_2_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(trans_2_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(trans_2_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(trans_2_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(trans_2_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(trans_2_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(trans_2_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(trans_2_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(trans_2_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(trans_2_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(trans_2_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(trans_2_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(trans_2_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(trans_2_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(trans_2_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(trans_2_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(trans_2_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(trans_2_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(trans_2_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(trans_2_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(trans_2_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(trans_2_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(trans_2_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(trans_2_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(trans_2_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(trans_2_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(trans_2_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(trans_2_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(trans_2_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(trans_2_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(trans_2_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(trans_2_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(trans_2_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(trans_2_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(trans_2_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(trans_2_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(trans_2_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(trans_2_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(trans_2_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(trans_2_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(trans_2_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(trans_2_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(trans_2_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(trans_2_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(trans_2_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(trans_2_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(trans_2_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(trans_2_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(trans_2_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(trans_2_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(trans_2_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(trans_2_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(trans_2_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(trans_2_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(trans_2_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(trans_2_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(trans_2_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(trans_2_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(trans_2_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(trans_2_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_header_0(trans_2_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(trans_2_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(trans_2_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(trans_2_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(trans_2_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(trans_2_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(trans_2_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(trans_2_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(trans_2_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(trans_2_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(trans_2_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(trans_2_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(trans_2_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(trans_2_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(trans_2_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(trans_2_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(trans_2_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(trans_2_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(trans_2_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(trans_2_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(trans_2_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(trans_2_io_pipe_phv_out_is_valid_processor),
    .io_pipe_phv_out_valid(trans_2_io_pipe_phv_out_valid),
    .io_pipe_phv_out_last(trans_2_io_pipe_phv_out_last),
    .io_next_proc_exist(trans_2_io_next_proc_exist)
  );
  InterProcessorTransfer trans_3 ( // @[ipsa.scala 79:25]
    .clock(trans_3_clock),
    .io_pipe_phv_in_data_0(trans_3_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(trans_3_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(trans_3_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(trans_3_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(trans_3_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(trans_3_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(trans_3_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(trans_3_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(trans_3_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(trans_3_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(trans_3_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(trans_3_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(trans_3_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(trans_3_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(trans_3_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(trans_3_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(trans_3_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(trans_3_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(trans_3_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(trans_3_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(trans_3_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(trans_3_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(trans_3_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(trans_3_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(trans_3_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(trans_3_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(trans_3_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(trans_3_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(trans_3_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(trans_3_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(trans_3_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(trans_3_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(trans_3_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(trans_3_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(trans_3_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(trans_3_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(trans_3_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(trans_3_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(trans_3_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(trans_3_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(trans_3_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(trans_3_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(trans_3_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(trans_3_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(trans_3_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(trans_3_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(trans_3_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(trans_3_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(trans_3_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(trans_3_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(trans_3_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(trans_3_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(trans_3_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(trans_3_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(trans_3_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(trans_3_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(trans_3_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(trans_3_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(trans_3_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(trans_3_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(trans_3_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(trans_3_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(trans_3_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(trans_3_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(trans_3_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(trans_3_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(trans_3_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(trans_3_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(trans_3_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(trans_3_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(trans_3_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(trans_3_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(trans_3_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(trans_3_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(trans_3_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(trans_3_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(trans_3_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(trans_3_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(trans_3_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(trans_3_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(trans_3_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(trans_3_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(trans_3_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(trans_3_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(trans_3_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(trans_3_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(trans_3_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(trans_3_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(trans_3_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(trans_3_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(trans_3_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(trans_3_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(trans_3_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(trans_3_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(trans_3_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(trans_3_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(trans_3_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(trans_3_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(trans_3_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(trans_3_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(trans_3_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(trans_3_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(trans_3_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(trans_3_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(trans_3_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(trans_3_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(trans_3_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(trans_3_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(trans_3_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(trans_3_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(trans_3_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(trans_3_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(trans_3_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(trans_3_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(trans_3_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(trans_3_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(trans_3_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(trans_3_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(trans_3_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(trans_3_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(trans_3_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(trans_3_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(trans_3_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(trans_3_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(trans_3_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(trans_3_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(trans_3_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(trans_3_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(trans_3_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(trans_3_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(trans_3_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(trans_3_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(trans_3_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(trans_3_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(trans_3_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(trans_3_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(trans_3_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(trans_3_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(trans_3_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(trans_3_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(trans_3_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(trans_3_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(trans_3_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(trans_3_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(trans_3_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(trans_3_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(trans_3_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(trans_3_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(trans_3_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(trans_3_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(trans_3_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(trans_3_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(trans_3_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(trans_3_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(trans_3_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(trans_3_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(trans_3_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(trans_3_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(trans_3_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(trans_3_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_header_0(trans_3_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(trans_3_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(trans_3_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(trans_3_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(trans_3_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(trans_3_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(trans_3_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(trans_3_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(trans_3_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(trans_3_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(trans_3_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(trans_3_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(trans_3_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(trans_3_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(trans_3_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(trans_3_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(trans_3_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(trans_3_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(trans_3_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(trans_3_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(trans_3_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_valid(trans_3_io_pipe_phv_in_valid),
    .io_pipe_phv_in_last(trans_3_io_pipe_phv_in_last),
    .io_pipe_phv_out_data_0(trans_3_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(trans_3_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(trans_3_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(trans_3_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(trans_3_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(trans_3_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(trans_3_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(trans_3_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(trans_3_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(trans_3_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(trans_3_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(trans_3_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(trans_3_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(trans_3_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(trans_3_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(trans_3_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(trans_3_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(trans_3_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(trans_3_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(trans_3_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(trans_3_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(trans_3_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(trans_3_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(trans_3_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(trans_3_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(trans_3_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(trans_3_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(trans_3_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(trans_3_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(trans_3_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(trans_3_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(trans_3_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(trans_3_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(trans_3_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(trans_3_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(trans_3_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(trans_3_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(trans_3_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(trans_3_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(trans_3_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(trans_3_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(trans_3_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(trans_3_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(trans_3_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(trans_3_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(trans_3_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(trans_3_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(trans_3_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(trans_3_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(trans_3_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(trans_3_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(trans_3_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(trans_3_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(trans_3_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(trans_3_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(trans_3_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(trans_3_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(trans_3_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(trans_3_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(trans_3_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(trans_3_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(trans_3_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(trans_3_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(trans_3_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(trans_3_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(trans_3_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(trans_3_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(trans_3_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(trans_3_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(trans_3_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(trans_3_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(trans_3_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(trans_3_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(trans_3_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(trans_3_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(trans_3_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(trans_3_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(trans_3_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(trans_3_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(trans_3_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(trans_3_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(trans_3_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(trans_3_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(trans_3_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(trans_3_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(trans_3_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(trans_3_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(trans_3_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(trans_3_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(trans_3_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(trans_3_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(trans_3_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(trans_3_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(trans_3_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(trans_3_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(trans_3_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(trans_3_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(trans_3_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(trans_3_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(trans_3_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(trans_3_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(trans_3_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(trans_3_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(trans_3_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(trans_3_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(trans_3_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(trans_3_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(trans_3_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(trans_3_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(trans_3_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(trans_3_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(trans_3_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(trans_3_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(trans_3_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(trans_3_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(trans_3_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(trans_3_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(trans_3_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(trans_3_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(trans_3_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(trans_3_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(trans_3_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(trans_3_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(trans_3_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(trans_3_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(trans_3_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(trans_3_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(trans_3_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(trans_3_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(trans_3_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(trans_3_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(trans_3_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(trans_3_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(trans_3_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(trans_3_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(trans_3_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(trans_3_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(trans_3_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(trans_3_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(trans_3_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(trans_3_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(trans_3_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(trans_3_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(trans_3_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(trans_3_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(trans_3_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(trans_3_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(trans_3_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(trans_3_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(trans_3_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(trans_3_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(trans_3_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(trans_3_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(trans_3_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(trans_3_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(trans_3_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(trans_3_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(trans_3_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(trans_3_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(trans_3_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_header_0(trans_3_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(trans_3_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(trans_3_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(trans_3_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(trans_3_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(trans_3_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(trans_3_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(trans_3_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(trans_3_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(trans_3_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(trans_3_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(trans_3_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(trans_3_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(trans_3_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(trans_3_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(trans_3_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(trans_3_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(trans_3_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(trans_3_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(trans_3_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(trans_3_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(trans_3_io_pipe_phv_out_is_valid_processor),
    .io_pipe_phv_out_valid(trans_3_io_pipe_phv_out_valid),
    .io_pipe_phv_out_last(trans_3_io_pipe_phv_out_last),
    .io_next_proc_exist(trans_3_io_next_proc_exist)
  );
  InterProcessorTransfer trans_4 ( // @[ipsa.scala 79:25]
    .clock(trans_4_clock),
    .io_pipe_phv_in_data_0(trans_4_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(trans_4_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(trans_4_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(trans_4_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(trans_4_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(trans_4_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(trans_4_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(trans_4_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(trans_4_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(trans_4_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(trans_4_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(trans_4_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(trans_4_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(trans_4_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(trans_4_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(trans_4_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(trans_4_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(trans_4_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(trans_4_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(trans_4_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(trans_4_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(trans_4_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(trans_4_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(trans_4_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(trans_4_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(trans_4_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(trans_4_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(trans_4_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(trans_4_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(trans_4_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(trans_4_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(trans_4_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(trans_4_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(trans_4_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(trans_4_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(trans_4_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(trans_4_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(trans_4_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(trans_4_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(trans_4_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(trans_4_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(trans_4_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(trans_4_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(trans_4_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(trans_4_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(trans_4_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(trans_4_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(trans_4_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(trans_4_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(trans_4_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(trans_4_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(trans_4_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(trans_4_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(trans_4_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(trans_4_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(trans_4_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(trans_4_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(trans_4_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(trans_4_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(trans_4_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(trans_4_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(trans_4_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(trans_4_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(trans_4_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(trans_4_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(trans_4_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(trans_4_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(trans_4_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(trans_4_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(trans_4_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(trans_4_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(trans_4_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(trans_4_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(trans_4_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(trans_4_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(trans_4_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(trans_4_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(trans_4_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(trans_4_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(trans_4_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(trans_4_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(trans_4_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(trans_4_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(trans_4_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(trans_4_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(trans_4_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(trans_4_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(trans_4_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(trans_4_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(trans_4_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(trans_4_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(trans_4_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(trans_4_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(trans_4_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(trans_4_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(trans_4_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(trans_4_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(trans_4_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(trans_4_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(trans_4_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(trans_4_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(trans_4_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(trans_4_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(trans_4_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(trans_4_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(trans_4_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(trans_4_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(trans_4_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(trans_4_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(trans_4_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(trans_4_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(trans_4_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(trans_4_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(trans_4_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(trans_4_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(trans_4_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(trans_4_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(trans_4_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(trans_4_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(trans_4_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(trans_4_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(trans_4_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(trans_4_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(trans_4_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(trans_4_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(trans_4_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(trans_4_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(trans_4_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(trans_4_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(trans_4_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(trans_4_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(trans_4_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(trans_4_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(trans_4_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(trans_4_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(trans_4_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(trans_4_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(trans_4_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(trans_4_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(trans_4_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(trans_4_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(trans_4_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(trans_4_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(trans_4_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(trans_4_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(trans_4_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(trans_4_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(trans_4_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(trans_4_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(trans_4_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(trans_4_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(trans_4_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(trans_4_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(trans_4_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(trans_4_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(trans_4_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(trans_4_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(trans_4_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(trans_4_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(trans_4_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_header_0(trans_4_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(trans_4_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(trans_4_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(trans_4_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(trans_4_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(trans_4_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(trans_4_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(trans_4_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(trans_4_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(trans_4_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(trans_4_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(trans_4_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(trans_4_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(trans_4_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(trans_4_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(trans_4_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(trans_4_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(trans_4_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(trans_4_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(trans_4_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(trans_4_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_valid(trans_4_io_pipe_phv_in_valid),
    .io_pipe_phv_in_last(trans_4_io_pipe_phv_in_last),
    .io_pipe_phv_out_data_0(trans_4_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(trans_4_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(trans_4_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(trans_4_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(trans_4_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(trans_4_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(trans_4_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(trans_4_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(trans_4_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(trans_4_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(trans_4_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(trans_4_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(trans_4_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(trans_4_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(trans_4_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(trans_4_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(trans_4_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(trans_4_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(trans_4_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(trans_4_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(trans_4_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(trans_4_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(trans_4_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(trans_4_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(trans_4_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(trans_4_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(trans_4_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(trans_4_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(trans_4_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(trans_4_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(trans_4_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(trans_4_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(trans_4_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(trans_4_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(trans_4_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(trans_4_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(trans_4_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(trans_4_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(trans_4_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(trans_4_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(trans_4_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(trans_4_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(trans_4_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(trans_4_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(trans_4_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(trans_4_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(trans_4_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(trans_4_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(trans_4_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(trans_4_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(trans_4_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(trans_4_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(trans_4_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(trans_4_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(trans_4_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(trans_4_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(trans_4_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(trans_4_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(trans_4_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(trans_4_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(trans_4_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(trans_4_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(trans_4_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(trans_4_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(trans_4_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(trans_4_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(trans_4_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(trans_4_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(trans_4_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(trans_4_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(trans_4_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(trans_4_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(trans_4_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(trans_4_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(trans_4_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(trans_4_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(trans_4_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(trans_4_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(trans_4_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(trans_4_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(trans_4_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(trans_4_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(trans_4_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(trans_4_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(trans_4_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(trans_4_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(trans_4_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(trans_4_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(trans_4_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(trans_4_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(trans_4_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(trans_4_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(trans_4_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(trans_4_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(trans_4_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(trans_4_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(trans_4_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(trans_4_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(trans_4_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(trans_4_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(trans_4_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(trans_4_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(trans_4_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(trans_4_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(trans_4_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(trans_4_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(trans_4_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(trans_4_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(trans_4_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(trans_4_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(trans_4_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(trans_4_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(trans_4_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(trans_4_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(trans_4_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(trans_4_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(trans_4_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(trans_4_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(trans_4_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(trans_4_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(trans_4_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(trans_4_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(trans_4_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(trans_4_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(trans_4_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(trans_4_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(trans_4_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(trans_4_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(trans_4_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(trans_4_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(trans_4_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(trans_4_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(trans_4_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(trans_4_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(trans_4_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(trans_4_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(trans_4_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(trans_4_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(trans_4_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(trans_4_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(trans_4_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(trans_4_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(trans_4_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(trans_4_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(trans_4_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(trans_4_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(trans_4_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(trans_4_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(trans_4_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(trans_4_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(trans_4_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(trans_4_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(trans_4_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(trans_4_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(trans_4_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(trans_4_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(trans_4_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(trans_4_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(trans_4_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(trans_4_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_header_0(trans_4_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(trans_4_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(trans_4_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(trans_4_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(trans_4_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(trans_4_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(trans_4_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(trans_4_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(trans_4_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(trans_4_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(trans_4_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(trans_4_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(trans_4_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(trans_4_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(trans_4_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(trans_4_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(trans_4_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(trans_4_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(trans_4_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(trans_4_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(trans_4_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(trans_4_io_pipe_phv_out_is_valid_processor),
    .io_pipe_phv_out_valid(trans_4_io_pipe_phv_out_valid),
    .io_pipe_phv_out_last(trans_4_io_pipe_phv_out_last),
    .io_next_proc_exist(trans_4_io_next_proc_exist)
  );
  InterProcessorTransfer trans_5 ( // @[ipsa.scala 79:25]
    .clock(trans_5_clock),
    .io_pipe_phv_in_data_0(trans_5_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(trans_5_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(trans_5_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(trans_5_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(trans_5_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(trans_5_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(trans_5_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(trans_5_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(trans_5_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(trans_5_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(trans_5_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(trans_5_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(trans_5_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(trans_5_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(trans_5_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(trans_5_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(trans_5_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(trans_5_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(trans_5_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(trans_5_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(trans_5_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(trans_5_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(trans_5_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(trans_5_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(trans_5_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(trans_5_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(trans_5_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(trans_5_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(trans_5_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(trans_5_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(trans_5_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(trans_5_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(trans_5_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(trans_5_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(trans_5_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(trans_5_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(trans_5_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(trans_5_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(trans_5_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(trans_5_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(trans_5_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(trans_5_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(trans_5_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(trans_5_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(trans_5_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(trans_5_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(trans_5_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(trans_5_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(trans_5_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(trans_5_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(trans_5_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(trans_5_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(trans_5_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(trans_5_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(trans_5_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(trans_5_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(trans_5_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(trans_5_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(trans_5_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(trans_5_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(trans_5_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(trans_5_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(trans_5_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(trans_5_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(trans_5_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(trans_5_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(trans_5_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(trans_5_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(trans_5_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(trans_5_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(trans_5_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(trans_5_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(trans_5_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(trans_5_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(trans_5_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(trans_5_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(trans_5_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(trans_5_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(trans_5_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(trans_5_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(trans_5_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(trans_5_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(trans_5_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(trans_5_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(trans_5_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(trans_5_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(trans_5_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(trans_5_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(trans_5_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(trans_5_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(trans_5_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(trans_5_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(trans_5_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(trans_5_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(trans_5_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(trans_5_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(trans_5_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(trans_5_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(trans_5_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(trans_5_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(trans_5_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(trans_5_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(trans_5_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(trans_5_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(trans_5_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(trans_5_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(trans_5_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(trans_5_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(trans_5_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(trans_5_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(trans_5_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(trans_5_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(trans_5_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(trans_5_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(trans_5_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(trans_5_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(trans_5_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(trans_5_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(trans_5_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(trans_5_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(trans_5_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(trans_5_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(trans_5_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(trans_5_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(trans_5_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(trans_5_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(trans_5_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(trans_5_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(trans_5_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(trans_5_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(trans_5_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(trans_5_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(trans_5_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(trans_5_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(trans_5_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(trans_5_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(trans_5_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(trans_5_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(trans_5_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(trans_5_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(trans_5_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(trans_5_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(trans_5_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(trans_5_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(trans_5_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(trans_5_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(trans_5_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(trans_5_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(trans_5_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(trans_5_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(trans_5_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(trans_5_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(trans_5_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(trans_5_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(trans_5_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(trans_5_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(trans_5_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(trans_5_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(trans_5_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(trans_5_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_header_0(trans_5_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(trans_5_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(trans_5_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(trans_5_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(trans_5_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(trans_5_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(trans_5_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(trans_5_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(trans_5_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(trans_5_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(trans_5_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(trans_5_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(trans_5_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(trans_5_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(trans_5_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(trans_5_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(trans_5_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(trans_5_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(trans_5_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(trans_5_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(trans_5_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_valid(trans_5_io_pipe_phv_in_valid),
    .io_pipe_phv_in_last(trans_5_io_pipe_phv_in_last),
    .io_pipe_phv_out_data_0(trans_5_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(trans_5_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(trans_5_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(trans_5_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(trans_5_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(trans_5_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(trans_5_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(trans_5_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(trans_5_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(trans_5_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(trans_5_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(trans_5_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(trans_5_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(trans_5_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(trans_5_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(trans_5_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(trans_5_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(trans_5_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(trans_5_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(trans_5_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(trans_5_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(trans_5_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(trans_5_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(trans_5_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(trans_5_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(trans_5_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(trans_5_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(trans_5_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(trans_5_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(trans_5_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(trans_5_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(trans_5_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(trans_5_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(trans_5_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(trans_5_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(trans_5_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(trans_5_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(trans_5_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(trans_5_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(trans_5_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(trans_5_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(trans_5_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(trans_5_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(trans_5_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(trans_5_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(trans_5_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(trans_5_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(trans_5_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(trans_5_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(trans_5_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(trans_5_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(trans_5_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(trans_5_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(trans_5_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(trans_5_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(trans_5_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(trans_5_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(trans_5_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(trans_5_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(trans_5_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(trans_5_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(trans_5_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(trans_5_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(trans_5_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(trans_5_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(trans_5_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(trans_5_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(trans_5_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(trans_5_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(trans_5_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(trans_5_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(trans_5_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(trans_5_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(trans_5_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(trans_5_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(trans_5_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(trans_5_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(trans_5_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(trans_5_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(trans_5_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(trans_5_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(trans_5_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(trans_5_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(trans_5_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(trans_5_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(trans_5_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(trans_5_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(trans_5_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(trans_5_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(trans_5_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(trans_5_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(trans_5_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(trans_5_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(trans_5_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(trans_5_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(trans_5_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(trans_5_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(trans_5_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(trans_5_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(trans_5_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(trans_5_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(trans_5_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(trans_5_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(trans_5_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(trans_5_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(trans_5_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(trans_5_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(trans_5_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(trans_5_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(trans_5_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(trans_5_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(trans_5_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(trans_5_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(trans_5_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(trans_5_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(trans_5_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(trans_5_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(trans_5_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(trans_5_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(trans_5_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(trans_5_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(trans_5_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(trans_5_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(trans_5_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(trans_5_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(trans_5_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(trans_5_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(trans_5_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(trans_5_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(trans_5_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(trans_5_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(trans_5_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(trans_5_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(trans_5_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(trans_5_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(trans_5_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(trans_5_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(trans_5_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(trans_5_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(trans_5_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(trans_5_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(trans_5_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(trans_5_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(trans_5_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(trans_5_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(trans_5_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(trans_5_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(trans_5_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(trans_5_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(trans_5_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(trans_5_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(trans_5_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(trans_5_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(trans_5_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(trans_5_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(trans_5_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(trans_5_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(trans_5_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(trans_5_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(trans_5_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_header_0(trans_5_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(trans_5_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(trans_5_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(trans_5_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(trans_5_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(trans_5_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(trans_5_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(trans_5_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(trans_5_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(trans_5_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(trans_5_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(trans_5_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(trans_5_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(trans_5_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(trans_5_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(trans_5_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(trans_5_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(trans_5_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(trans_5_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(trans_5_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(trans_5_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(trans_5_io_pipe_phv_out_is_valid_processor),
    .io_pipe_phv_out_valid(trans_5_io_pipe_phv_out_valid),
    .io_pipe_phv_out_last(trans_5_io_pipe_phv_out_last),
    .io_next_proc_exist(trans_5_io_next_proc_exist)
  );
  InterProcessorTransfer trans_6 ( // @[ipsa.scala 79:25]
    .clock(trans_6_clock),
    .io_pipe_phv_in_data_0(trans_6_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(trans_6_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(trans_6_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(trans_6_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(trans_6_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(trans_6_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(trans_6_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(trans_6_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(trans_6_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(trans_6_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(trans_6_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(trans_6_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(trans_6_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(trans_6_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(trans_6_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(trans_6_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(trans_6_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(trans_6_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(trans_6_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(trans_6_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(trans_6_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(trans_6_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(trans_6_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(trans_6_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(trans_6_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(trans_6_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(trans_6_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(trans_6_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(trans_6_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(trans_6_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(trans_6_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(trans_6_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(trans_6_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(trans_6_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(trans_6_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(trans_6_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(trans_6_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(trans_6_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(trans_6_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(trans_6_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(trans_6_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(trans_6_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(trans_6_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(trans_6_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(trans_6_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(trans_6_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(trans_6_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(trans_6_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(trans_6_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(trans_6_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(trans_6_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(trans_6_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(trans_6_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(trans_6_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(trans_6_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(trans_6_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(trans_6_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(trans_6_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(trans_6_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(trans_6_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(trans_6_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(trans_6_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(trans_6_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(trans_6_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(trans_6_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(trans_6_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(trans_6_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(trans_6_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(trans_6_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(trans_6_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(trans_6_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(trans_6_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(trans_6_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(trans_6_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(trans_6_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(trans_6_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(trans_6_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(trans_6_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(trans_6_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(trans_6_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(trans_6_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(trans_6_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(trans_6_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(trans_6_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(trans_6_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(trans_6_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(trans_6_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(trans_6_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(trans_6_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(trans_6_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(trans_6_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(trans_6_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(trans_6_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(trans_6_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(trans_6_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(trans_6_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(trans_6_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(trans_6_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(trans_6_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(trans_6_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(trans_6_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(trans_6_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(trans_6_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(trans_6_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(trans_6_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(trans_6_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(trans_6_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(trans_6_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(trans_6_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(trans_6_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(trans_6_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(trans_6_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(trans_6_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(trans_6_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(trans_6_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(trans_6_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(trans_6_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(trans_6_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(trans_6_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(trans_6_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(trans_6_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(trans_6_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(trans_6_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(trans_6_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(trans_6_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(trans_6_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(trans_6_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(trans_6_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(trans_6_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(trans_6_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(trans_6_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(trans_6_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(trans_6_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(trans_6_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(trans_6_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(trans_6_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(trans_6_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(trans_6_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(trans_6_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(trans_6_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(trans_6_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(trans_6_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(trans_6_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(trans_6_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(trans_6_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(trans_6_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(trans_6_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(trans_6_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(trans_6_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(trans_6_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(trans_6_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(trans_6_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(trans_6_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(trans_6_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(trans_6_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(trans_6_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(trans_6_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(trans_6_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(trans_6_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(trans_6_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_header_0(trans_6_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(trans_6_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(trans_6_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(trans_6_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(trans_6_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(trans_6_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(trans_6_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(trans_6_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(trans_6_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(trans_6_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(trans_6_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(trans_6_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(trans_6_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(trans_6_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(trans_6_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(trans_6_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(trans_6_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(trans_6_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(trans_6_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(trans_6_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(trans_6_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_valid(trans_6_io_pipe_phv_in_valid),
    .io_pipe_phv_in_last(trans_6_io_pipe_phv_in_last),
    .io_pipe_phv_out_data_0(trans_6_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(trans_6_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(trans_6_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(trans_6_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(trans_6_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(trans_6_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(trans_6_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(trans_6_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(trans_6_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(trans_6_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(trans_6_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(trans_6_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(trans_6_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(trans_6_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(trans_6_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(trans_6_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(trans_6_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(trans_6_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(trans_6_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(trans_6_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(trans_6_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(trans_6_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(trans_6_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(trans_6_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(trans_6_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(trans_6_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(trans_6_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(trans_6_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(trans_6_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(trans_6_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(trans_6_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(trans_6_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(trans_6_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(trans_6_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(trans_6_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(trans_6_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(trans_6_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(trans_6_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(trans_6_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(trans_6_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(trans_6_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(trans_6_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(trans_6_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(trans_6_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(trans_6_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(trans_6_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(trans_6_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(trans_6_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(trans_6_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(trans_6_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(trans_6_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(trans_6_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(trans_6_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(trans_6_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(trans_6_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(trans_6_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(trans_6_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(trans_6_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(trans_6_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(trans_6_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(trans_6_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(trans_6_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(trans_6_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(trans_6_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(trans_6_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(trans_6_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(trans_6_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(trans_6_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(trans_6_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(trans_6_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(trans_6_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(trans_6_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(trans_6_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(trans_6_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(trans_6_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(trans_6_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(trans_6_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(trans_6_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(trans_6_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(trans_6_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(trans_6_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(trans_6_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(trans_6_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(trans_6_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(trans_6_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(trans_6_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(trans_6_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(trans_6_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(trans_6_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(trans_6_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(trans_6_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(trans_6_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(trans_6_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(trans_6_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(trans_6_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(trans_6_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(trans_6_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(trans_6_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(trans_6_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(trans_6_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(trans_6_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(trans_6_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(trans_6_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(trans_6_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(trans_6_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(trans_6_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(trans_6_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(trans_6_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(trans_6_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(trans_6_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(trans_6_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(trans_6_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(trans_6_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(trans_6_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(trans_6_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(trans_6_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(trans_6_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(trans_6_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(trans_6_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(trans_6_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(trans_6_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(trans_6_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(trans_6_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(trans_6_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(trans_6_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(trans_6_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(trans_6_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(trans_6_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(trans_6_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(trans_6_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(trans_6_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(trans_6_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(trans_6_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(trans_6_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(trans_6_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(trans_6_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(trans_6_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(trans_6_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(trans_6_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(trans_6_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(trans_6_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(trans_6_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(trans_6_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(trans_6_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(trans_6_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(trans_6_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(trans_6_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(trans_6_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(trans_6_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(trans_6_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(trans_6_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(trans_6_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(trans_6_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(trans_6_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(trans_6_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(trans_6_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(trans_6_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(trans_6_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(trans_6_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(trans_6_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_header_0(trans_6_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(trans_6_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(trans_6_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(trans_6_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(trans_6_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(trans_6_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(trans_6_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(trans_6_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(trans_6_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(trans_6_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(trans_6_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(trans_6_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(trans_6_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(trans_6_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(trans_6_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(trans_6_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(trans_6_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(trans_6_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(trans_6_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(trans_6_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(trans_6_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(trans_6_io_pipe_phv_out_is_valid_processor),
    .io_pipe_phv_out_valid(trans_6_io_pipe_phv_out_valid),
    .io_pipe_phv_out_last(trans_6_io_pipe_phv_out_last),
    .io_next_proc_exist(trans_6_io_next_proc_exist)
  );
  InterProcessorTransfer trans_7 ( // @[ipsa.scala 79:25]
    .clock(trans_7_clock),
    .io_pipe_phv_in_data_0(trans_7_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(trans_7_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(trans_7_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(trans_7_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(trans_7_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(trans_7_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(trans_7_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(trans_7_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(trans_7_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(trans_7_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(trans_7_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(trans_7_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(trans_7_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(trans_7_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(trans_7_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(trans_7_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(trans_7_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(trans_7_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(trans_7_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(trans_7_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(trans_7_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(trans_7_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(trans_7_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(trans_7_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(trans_7_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(trans_7_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(trans_7_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(trans_7_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(trans_7_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(trans_7_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(trans_7_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(trans_7_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(trans_7_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(trans_7_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(trans_7_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(trans_7_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(trans_7_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(trans_7_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(trans_7_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(trans_7_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(trans_7_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(trans_7_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(trans_7_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(trans_7_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(trans_7_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(trans_7_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(trans_7_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(trans_7_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(trans_7_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(trans_7_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(trans_7_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(trans_7_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(trans_7_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(trans_7_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(trans_7_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(trans_7_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(trans_7_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(trans_7_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(trans_7_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(trans_7_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(trans_7_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(trans_7_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(trans_7_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(trans_7_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(trans_7_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(trans_7_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(trans_7_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(trans_7_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(trans_7_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(trans_7_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(trans_7_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(trans_7_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(trans_7_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(trans_7_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(trans_7_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(trans_7_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(trans_7_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(trans_7_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(trans_7_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(trans_7_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(trans_7_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(trans_7_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(trans_7_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(trans_7_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(trans_7_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(trans_7_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(trans_7_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(trans_7_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(trans_7_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(trans_7_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(trans_7_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(trans_7_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(trans_7_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(trans_7_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(trans_7_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(trans_7_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(trans_7_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(trans_7_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(trans_7_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(trans_7_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(trans_7_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(trans_7_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(trans_7_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(trans_7_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(trans_7_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(trans_7_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(trans_7_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(trans_7_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(trans_7_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(trans_7_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(trans_7_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(trans_7_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(trans_7_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(trans_7_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(trans_7_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(trans_7_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(trans_7_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(trans_7_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(trans_7_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(trans_7_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(trans_7_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(trans_7_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(trans_7_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(trans_7_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(trans_7_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(trans_7_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(trans_7_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(trans_7_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(trans_7_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(trans_7_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(trans_7_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(trans_7_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(trans_7_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(trans_7_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(trans_7_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(trans_7_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(trans_7_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(trans_7_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(trans_7_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(trans_7_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(trans_7_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(trans_7_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(trans_7_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(trans_7_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(trans_7_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(trans_7_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(trans_7_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(trans_7_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(trans_7_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(trans_7_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(trans_7_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(trans_7_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(trans_7_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(trans_7_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(trans_7_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(trans_7_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(trans_7_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(trans_7_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(trans_7_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(trans_7_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_header_0(trans_7_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(trans_7_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(trans_7_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(trans_7_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(trans_7_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(trans_7_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(trans_7_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(trans_7_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(trans_7_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(trans_7_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(trans_7_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(trans_7_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(trans_7_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(trans_7_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(trans_7_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(trans_7_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(trans_7_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(trans_7_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(trans_7_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(trans_7_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(trans_7_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_valid(trans_7_io_pipe_phv_in_valid),
    .io_pipe_phv_in_last(trans_7_io_pipe_phv_in_last),
    .io_pipe_phv_out_data_0(trans_7_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(trans_7_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(trans_7_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(trans_7_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(trans_7_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(trans_7_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(trans_7_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(trans_7_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(trans_7_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(trans_7_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(trans_7_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(trans_7_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(trans_7_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(trans_7_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(trans_7_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(trans_7_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(trans_7_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(trans_7_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(trans_7_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(trans_7_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(trans_7_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(trans_7_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(trans_7_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(trans_7_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(trans_7_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(trans_7_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(trans_7_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(trans_7_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(trans_7_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(trans_7_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(trans_7_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(trans_7_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(trans_7_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(trans_7_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(trans_7_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(trans_7_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(trans_7_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(trans_7_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(trans_7_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(trans_7_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(trans_7_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(trans_7_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(trans_7_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(trans_7_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(trans_7_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(trans_7_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(trans_7_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(trans_7_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(trans_7_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(trans_7_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(trans_7_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(trans_7_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(trans_7_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(trans_7_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(trans_7_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(trans_7_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(trans_7_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(trans_7_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(trans_7_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(trans_7_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(trans_7_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(trans_7_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(trans_7_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(trans_7_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(trans_7_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(trans_7_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(trans_7_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(trans_7_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(trans_7_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(trans_7_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(trans_7_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(trans_7_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(trans_7_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(trans_7_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(trans_7_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(trans_7_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(trans_7_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(trans_7_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(trans_7_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(trans_7_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(trans_7_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(trans_7_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(trans_7_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(trans_7_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(trans_7_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(trans_7_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(trans_7_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(trans_7_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(trans_7_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(trans_7_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(trans_7_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(trans_7_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(trans_7_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(trans_7_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(trans_7_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(trans_7_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(trans_7_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(trans_7_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(trans_7_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(trans_7_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(trans_7_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(trans_7_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(trans_7_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(trans_7_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(trans_7_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(trans_7_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(trans_7_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(trans_7_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(trans_7_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(trans_7_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(trans_7_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(trans_7_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(trans_7_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(trans_7_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(trans_7_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(trans_7_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(trans_7_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(trans_7_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(trans_7_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(trans_7_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(trans_7_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(trans_7_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(trans_7_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(trans_7_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(trans_7_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(trans_7_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(trans_7_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(trans_7_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(trans_7_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(trans_7_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(trans_7_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(trans_7_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(trans_7_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(trans_7_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(trans_7_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(trans_7_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(trans_7_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(trans_7_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(trans_7_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(trans_7_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(trans_7_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(trans_7_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(trans_7_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(trans_7_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(trans_7_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(trans_7_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(trans_7_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(trans_7_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(trans_7_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(trans_7_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(trans_7_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(trans_7_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(trans_7_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(trans_7_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(trans_7_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(trans_7_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(trans_7_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(trans_7_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(trans_7_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(trans_7_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_header_0(trans_7_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(trans_7_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(trans_7_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(trans_7_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(trans_7_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(trans_7_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(trans_7_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(trans_7_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(trans_7_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(trans_7_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(trans_7_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(trans_7_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(trans_7_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(trans_7_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(trans_7_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(trans_7_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(trans_7_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(trans_7_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(trans_7_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(trans_7_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(trans_7_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(trans_7_io_pipe_phv_out_is_valid_processor),
    .io_pipe_phv_out_valid(trans_7_io_pipe_phv_out_valid),
    .io_pipe_phv_out_last(trans_7_io_pipe_phv_out_last),
    .io_next_proc_exist(trans_7_io_next_proc_exist)
  );
  InterProcessorTransfer trans_8 ( // @[ipsa.scala 79:25]
    .clock(trans_8_clock),
    .io_pipe_phv_in_data_0(trans_8_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(trans_8_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(trans_8_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(trans_8_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(trans_8_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(trans_8_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(trans_8_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(trans_8_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(trans_8_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(trans_8_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(trans_8_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(trans_8_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(trans_8_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(trans_8_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(trans_8_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(trans_8_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(trans_8_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(trans_8_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(trans_8_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(trans_8_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(trans_8_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(trans_8_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(trans_8_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(trans_8_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(trans_8_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(trans_8_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(trans_8_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(trans_8_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(trans_8_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(trans_8_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(trans_8_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(trans_8_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(trans_8_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(trans_8_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(trans_8_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(trans_8_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(trans_8_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(trans_8_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(trans_8_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(trans_8_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(trans_8_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(trans_8_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(trans_8_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(trans_8_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(trans_8_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(trans_8_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(trans_8_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(trans_8_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(trans_8_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(trans_8_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(trans_8_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(trans_8_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(trans_8_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(trans_8_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(trans_8_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(trans_8_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(trans_8_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(trans_8_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(trans_8_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(trans_8_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(trans_8_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(trans_8_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(trans_8_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(trans_8_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(trans_8_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(trans_8_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(trans_8_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(trans_8_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(trans_8_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(trans_8_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(trans_8_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(trans_8_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(trans_8_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(trans_8_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(trans_8_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(trans_8_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(trans_8_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(trans_8_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(trans_8_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(trans_8_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(trans_8_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(trans_8_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(trans_8_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(trans_8_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(trans_8_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(trans_8_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(trans_8_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(trans_8_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(trans_8_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(trans_8_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(trans_8_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(trans_8_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(trans_8_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(trans_8_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(trans_8_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(trans_8_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(trans_8_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(trans_8_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(trans_8_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(trans_8_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(trans_8_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(trans_8_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(trans_8_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(trans_8_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(trans_8_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(trans_8_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(trans_8_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(trans_8_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(trans_8_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(trans_8_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(trans_8_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(trans_8_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(trans_8_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(trans_8_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(trans_8_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(trans_8_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(trans_8_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(trans_8_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(trans_8_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(trans_8_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(trans_8_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(trans_8_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(trans_8_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(trans_8_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(trans_8_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(trans_8_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(trans_8_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(trans_8_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(trans_8_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(trans_8_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(trans_8_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(trans_8_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(trans_8_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(trans_8_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(trans_8_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(trans_8_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(trans_8_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(trans_8_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(trans_8_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(trans_8_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(trans_8_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(trans_8_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(trans_8_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(trans_8_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(trans_8_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(trans_8_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(trans_8_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(trans_8_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(trans_8_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(trans_8_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(trans_8_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(trans_8_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(trans_8_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(trans_8_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(trans_8_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(trans_8_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(trans_8_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(trans_8_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(trans_8_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(trans_8_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_header_0(trans_8_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(trans_8_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(trans_8_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(trans_8_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(trans_8_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(trans_8_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(trans_8_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(trans_8_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(trans_8_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(trans_8_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(trans_8_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(trans_8_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(trans_8_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(trans_8_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(trans_8_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(trans_8_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(trans_8_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(trans_8_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(trans_8_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(trans_8_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(trans_8_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_valid(trans_8_io_pipe_phv_in_valid),
    .io_pipe_phv_in_last(trans_8_io_pipe_phv_in_last),
    .io_pipe_phv_out_data_0(trans_8_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(trans_8_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(trans_8_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(trans_8_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(trans_8_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(trans_8_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(trans_8_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(trans_8_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(trans_8_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(trans_8_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(trans_8_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(trans_8_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(trans_8_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(trans_8_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(trans_8_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(trans_8_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(trans_8_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(trans_8_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(trans_8_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(trans_8_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(trans_8_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(trans_8_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(trans_8_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(trans_8_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(trans_8_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(trans_8_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(trans_8_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(trans_8_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(trans_8_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(trans_8_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(trans_8_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(trans_8_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(trans_8_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(trans_8_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(trans_8_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(trans_8_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(trans_8_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(trans_8_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(trans_8_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(trans_8_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(trans_8_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(trans_8_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(trans_8_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(trans_8_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(trans_8_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(trans_8_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(trans_8_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(trans_8_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(trans_8_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(trans_8_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(trans_8_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(trans_8_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(trans_8_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(trans_8_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(trans_8_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(trans_8_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(trans_8_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(trans_8_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(trans_8_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(trans_8_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(trans_8_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(trans_8_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(trans_8_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(trans_8_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(trans_8_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(trans_8_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(trans_8_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(trans_8_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(trans_8_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(trans_8_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(trans_8_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(trans_8_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(trans_8_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(trans_8_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(trans_8_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(trans_8_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(trans_8_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(trans_8_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(trans_8_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(trans_8_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(trans_8_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(trans_8_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(trans_8_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(trans_8_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(trans_8_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(trans_8_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(trans_8_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(trans_8_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(trans_8_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(trans_8_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(trans_8_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(trans_8_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(trans_8_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(trans_8_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(trans_8_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(trans_8_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(trans_8_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(trans_8_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(trans_8_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(trans_8_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(trans_8_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(trans_8_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(trans_8_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(trans_8_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(trans_8_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(trans_8_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(trans_8_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(trans_8_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(trans_8_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(trans_8_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(trans_8_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(trans_8_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(trans_8_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(trans_8_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(trans_8_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(trans_8_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(trans_8_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(trans_8_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(trans_8_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(trans_8_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(trans_8_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(trans_8_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(trans_8_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(trans_8_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(trans_8_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(trans_8_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(trans_8_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(trans_8_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(trans_8_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(trans_8_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(trans_8_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(trans_8_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(trans_8_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(trans_8_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(trans_8_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(trans_8_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(trans_8_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(trans_8_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(trans_8_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(trans_8_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(trans_8_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(trans_8_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(trans_8_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(trans_8_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(trans_8_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(trans_8_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(trans_8_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(trans_8_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(trans_8_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(trans_8_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(trans_8_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(trans_8_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(trans_8_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(trans_8_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(trans_8_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(trans_8_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(trans_8_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(trans_8_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(trans_8_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(trans_8_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_header_0(trans_8_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(trans_8_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(trans_8_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(trans_8_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(trans_8_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(trans_8_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(trans_8_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(trans_8_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(trans_8_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(trans_8_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(trans_8_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(trans_8_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(trans_8_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(trans_8_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(trans_8_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(trans_8_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(trans_8_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(trans_8_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(trans_8_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(trans_8_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(trans_8_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(trans_8_io_pipe_phv_out_is_valid_processor),
    .io_pipe_phv_out_valid(trans_8_io_pipe_phv_out_valid),
    .io_pipe_phv_out_last(trans_8_io_pipe_phv_out_last),
    .io_next_proc_exist(trans_8_io_next_proc_exist)
  );
  InterProcessorTransfer trans_9 ( // @[ipsa.scala 79:25]
    .clock(trans_9_clock),
    .io_pipe_phv_in_data_0(trans_9_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(trans_9_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(trans_9_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(trans_9_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(trans_9_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(trans_9_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(trans_9_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(trans_9_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(trans_9_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(trans_9_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(trans_9_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(trans_9_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(trans_9_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(trans_9_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(trans_9_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(trans_9_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(trans_9_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(trans_9_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(trans_9_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(trans_9_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(trans_9_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(trans_9_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(trans_9_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(trans_9_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(trans_9_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(trans_9_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(trans_9_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(trans_9_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(trans_9_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(trans_9_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(trans_9_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(trans_9_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(trans_9_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(trans_9_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(trans_9_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(trans_9_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(trans_9_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(trans_9_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(trans_9_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(trans_9_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(trans_9_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(trans_9_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(trans_9_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(trans_9_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(trans_9_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(trans_9_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(trans_9_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(trans_9_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(trans_9_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(trans_9_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(trans_9_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(trans_9_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(trans_9_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(trans_9_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(trans_9_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(trans_9_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(trans_9_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(trans_9_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(trans_9_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(trans_9_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(trans_9_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(trans_9_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(trans_9_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(trans_9_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(trans_9_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(trans_9_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(trans_9_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(trans_9_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(trans_9_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(trans_9_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(trans_9_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(trans_9_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(trans_9_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(trans_9_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(trans_9_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(trans_9_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(trans_9_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(trans_9_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(trans_9_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(trans_9_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(trans_9_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(trans_9_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(trans_9_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(trans_9_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(trans_9_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(trans_9_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(trans_9_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(trans_9_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(trans_9_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(trans_9_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(trans_9_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(trans_9_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(trans_9_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(trans_9_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(trans_9_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(trans_9_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(trans_9_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(trans_9_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(trans_9_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(trans_9_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(trans_9_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(trans_9_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(trans_9_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(trans_9_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(trans_9_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(trans_9_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(trans_9_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(trans_9_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(trans_9_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(trans_9_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(trans_9_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(trans_9_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(trans_9_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(trans_9_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(trans_9_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(trans_9_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(trans_9_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(trans_9_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(trans_9_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(trans_9_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(trans_9_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(trans_9_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(trans_9_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(trans_9_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(trans_9_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(trans_9_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(trans_9_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(trans_9_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(trans_9_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(trans_9_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(trans_9_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(trans_9_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(trans_9_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(trans_9_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(trans_9_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(trans_9_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(trans_9_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(trans_9_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(trans_9_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(trans_9_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(trans_9_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(trans_9_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(trans_9_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(trans_9_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(trans_9_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(trans_9_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(trans_9_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(trans_9_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(trans_9_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(trans_9_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(trans_9_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(trans_9_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(trans_9_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(trans_9_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(trans_9_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(trans_9_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(trans_9_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(trans_9_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(trans_9_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(trans_9_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_header_0(trans_9_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(trans_9_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(trans_9_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(trans_9_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(trans_9_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(trans_9_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(trans_9_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(trans_9_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(trans_9_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(trans_9_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(trans_9_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(trans_9_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(trans_9_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(trans_9_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(trans_9_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(trans_9_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(trans_9_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(trans_9_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(trans_9_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(trans_9_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(trans_9_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_valid(trans_9_io_pipe_phv_in_valid),
    .io_pipe_phv_in_last(trans_9_io_pipe_phv_in_last),
    .io_pipe_phv_out_data_0(trans_9_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(trans_9_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(trans_9_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(trans_9_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(trans_9_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(trans_9_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(trans_9_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(trans_9_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(trans_9_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(trans_9_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(trans_9_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(trans_9_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(trans_9_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(trans_9_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(trans_9_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(trans_9_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(trans_9_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(trans_9_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(trans_9_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(trans_9_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(trans_9_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(trans_9_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(trans_9_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(trans_9_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(trans_9_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(trans_9_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(trans_9_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(trans_9_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(trans_9_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(trans_9_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(trans_9_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(trans_9_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(trans_9_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(trans_9_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(trans_9_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(trans_9_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(trans_9_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(trans_9_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(trans_9_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(trans_9_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(trans_9_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(trans_9_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(trans_9_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(trans_9_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(trans_9_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(trans_9_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(trans_9_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(trans_9_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(trans_9_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(trans_9_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(trans_9_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(trans_9_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(trans_9_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(trans_9_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(trans_9_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(trans_9_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(trans_9_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(trans_9_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(trans_9_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(trans_9_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(trans_9_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(trans_9_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(trans_9_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(trans_9_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(trans_9_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(trans_9_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(trans_9_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(trans_9_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(trans_9_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(trans_9_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(trans_9_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(trans_9_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(trans_9_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(trans_9_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(trans_9_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(trans_9_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(trans_9_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(trans_9_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(trans_9_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(trans_9_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(trans_9_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(trans_9_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(trans_9_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(trans_9_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(trans_9_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(trans_9_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(trans_9_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(trans_9_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(trans_9_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(trans_9_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(trans_9_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(trans_9_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(trans_9_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(trans_9_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(trans_9_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(trans_9_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(trans_9_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(trans_9_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(trans_9_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(trans_9_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(trans_9_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(trans_9_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(trans_9_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(trans_9_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(trans_9_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(trans_9_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(trans_9_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(trans_9_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(trans_9_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(trans_9_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(trans_9_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(trans_9_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(trans_9_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(trans_9_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(trans_9_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(trans_9_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(trans_9_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(trans_9_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(trans_9_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(trans_9_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(trans_9_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(trans_9_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(trans_9_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(trans_9_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(trans_9_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(trans_9_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(trans_9_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(trans_9_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(trans_9_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(trans_9_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(trans_9_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(trans_9_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(trans_9_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(trans_9_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(trans_9_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(trans_9_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(trans_9_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(trans_9_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(trans_9_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(trans_9_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(trans_9_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(trans_9_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(trans_9_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(trans_9_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(trans_9_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(trans_9_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(trans_9_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(trans_9_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(trans_9_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(trans_9_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(trans_9_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(trans_9_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(trans_9_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(trans_9_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(trans_9_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(trans_9_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(trans_9_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(trans_9_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(trans_9_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(trans_9_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_header_0(trans_9_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(trans_9_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(trans_9_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(trans_9_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(trans_9_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(trans_9_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(trans_9_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(trans_9_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(trans_9_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(trans_9_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(trans_9_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(trans_9_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(trans_9_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(trans_9_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(trans_9_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(trans_9_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(trans_9_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(trans_9_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(trans_9_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(trans_9_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(trans_9_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(trans_9_io_pipe_phv_out_is_valid_processor),
    .io_pipe_phv_out_valid(trans_9_io_pipe_phv_out_valid),
    .io_pipe_phv_out_last(trans_9_io_pipe_phv_out_last),
    .io_next_proc_exist(trans_9_io_next_proc_exist)
  );
  InterProcessorTransfer trans_10 ( // @[ipsa.scala 79:25]
    .clock(trans_10_clock),
    .io_pipe_phv_in_data_0(trans_10_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(trans_10_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(trans_10_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(trans_10_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(trans_10_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(trans_10_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(trans_10_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(trans_10_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(trans_10_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(trans_10_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(trans_10_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(trans_10_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(trans_10_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(trans_10_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(trans_10_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(trans_10_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(trans_10_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(trans_10_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(trans_10_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(trans_10_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(trans_10_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(trans_10_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(trans_10_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(trans_10_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(trans_10_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(trans_10_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(trans_10_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(trans_10_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(trans_10_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(trans_10_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(trans_10_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(trans_10_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(trans_10_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(trans_10_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(trans_10_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(trans_10_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(trans_10_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(trans_10_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(trans_10_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(trans_10_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(trans_10_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(trans_10_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(trans_10_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(trans_10_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(trans_10_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(trans_10_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(trans_10_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(trans_10_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(trans_10_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(trans_10_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(trans_10_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(trans_10_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(trans_10_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(trans_10_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(trans_10_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(trans_10_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(trans_10_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(trans_10_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(trans_10_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(trans_10_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(trans_10_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(trans_10_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(trans_10_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(trans_10_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(trans_10_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(trans_10_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(trans_10_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(trans_10_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(trans_10_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(trans_10_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(trans_10_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(trans_10_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(trans_10_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(trans_10_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(trans_10_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(trans_10_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(trans_10_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(trans_10_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(trans_10_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(trans_10_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(trans_10_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(trans_10_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(trans_10_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(trans_10_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(trans_10_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(trans_10_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(trans_10_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(trans_10_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(trans_10_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(trans_10_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(trans_10_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(trans_10_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(trans_10_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(trans_10_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(trans_10_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(trans_10_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(trans_10_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(trans_10_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(trans_10_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(trans_10_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(trans_10_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(trans_10_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(trans_10_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(trans_10_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(trans_10_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(trans_10_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(trans_10_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(trans_10_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(trans_10_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(trans_10_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(trans_10_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(trans_10_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(trans_10_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(trans_10_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(trans_10_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(trans_10_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(trans_10_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(trans_10_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(trans_10_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(trans_10_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(trans_10_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(trans_10_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(trans_10_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(trans_10_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(trans_10_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(trans_10_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(trans_10_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(trans_10_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(trans_10_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(trans_10_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(trans_10_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(trans_10_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(trans_10_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(trans_10_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(trans_10_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(trans_10_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(trans_10_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(trans_10_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(trans_10_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(trans_10_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(trans_10_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(trans_10_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(trans_10_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(trans_10_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(trans_10_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(trans_10_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(trans_10_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(trans_10_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(trans_10_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(trans_10_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(trans_10_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(trans_10_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(trans_10_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(trans_10_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(trans_10_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(trans_10_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(trans_10_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(trans_10_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(trans_10_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(trans_10_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_header_0(trans_10_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(trans_10_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(trans_10_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(trans_10_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(trans_10_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(trans_10_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(trans_10_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(trans_10_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(trans_10_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(trans_10_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(trans_10_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(trans_10_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(trans_10_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(trans_10_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(trans_10_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(trans_10_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(trans_10_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(trans_10_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(trans_10_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(trans_10_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(trans_10_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_valid(trans_10_io_pipe_phv_in_valid),
    .io_pipe_phv_in_last(trans_10_io_pipe_phv_in_last),
    .io_pipe_phv_out_data_0(trans_10_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(trans_10_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(trans_10_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(trans_10_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(trans_10_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(trans_10_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(trans_10_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(trans_10_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(trans_10_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(trans_10_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(trans_10_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(trans_10_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(trans_10_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(trans_10_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(trans_10_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(trans_10_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(trans_10_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(trans_10_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(trans_10_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(trans_10_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(trans_10_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(trans_10_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(trans_10_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(trans_10_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(trans_10_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(trans_10_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(trans_10_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(trans_10_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(trans_10_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(trans_10_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(trans_10_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(trans_10_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(trans_10_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(trans_10_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(trans_10_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(trans_10_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(trans_10_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(trans_10_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(trans_10_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(trans_10_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(trans_10_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(trans_10_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(trans_10_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(trans_10_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(trans_10_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(trans_10_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(trans_10_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(trans_10_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(trans_10_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(trans_10_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(trans_10_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(trans_10_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(trans_10_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(trans_10_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(trans_10_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(trans_10_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(trans_10_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(trans_10_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(trans_10_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(trans_10_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(trans_10_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(trans_10_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(trans_10_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(trans_10_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(trans_10_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(trans_10_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(trans_10_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(trans_10_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(trans_10_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(trans_10_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(trans_10_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(trans_10_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(trans_10_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(trans_10_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(trans_10_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(trans_10_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(trans_10_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(trans_10_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(trans_10_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(trans_10_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(trans_10_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(trans_10_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(trans_10_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(trans_10_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(trans_10_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(trans_10_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(trans_10_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(trans_10_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(trans_10_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(trans_10_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(trans_10_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(trans_10_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(trans_10_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(trans_10_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(trans_10_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(trans_10_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(trans_10_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(trans_10_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(trans_10_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(trans_10_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(trans_10_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(trans_10_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(trans_10_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(trans_10_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(trans_10_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(trans_10_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(trans_10_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(trans_10_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(trans_10_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(trans_10_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(trans_10_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(trans_10_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(trans_10_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(trans_10_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(trans_10_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(trans_10_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(trans_10_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(trans_10_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(trans_10_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(trans_10_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(trans_10_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(trans_10_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(trans_10_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(trans_10_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(trans_10_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(trans_10_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(trans_10_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(trans_10_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(trans_10_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(trans_10_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(trans_10_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(trans_10_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(trans_10_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(trans_10_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(trans_10_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(trans_10_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(trans_10_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(trans_10_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(trans_10_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(trans_10_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(trans_10_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(trans_10_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(trans_10_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(trans_10_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(trans_10_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(trans_10_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(trans_10_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(trans_10_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(trans_10_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(trans_10_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(trans_10_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(trans_10_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(trans_10_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(trans_10_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(trans_10_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(trans_10_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(trans_10_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(trans_10_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(trans_10_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(trans_10_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_header_0(trans_10_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(trans_10_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(trans_10_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(trans_10_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(trans_10_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(trans_10_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(trans_10_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(trans_10_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(trans_10_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(trans_10_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(trans_10_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(trans_10_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(trans_10_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(trans_10_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(trans_10_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(trans_10_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(trans_10_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(trans_10_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(trans_10_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(trans_10_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(trans_10_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(trans_10_io_pipe_phv_out_is_valid_processor),
    .io_pipe_phv_out_valid(trans_10_io_pipe_phv_out_valid),
    .io_pipe_phv_out_last(trans_10_io_pipe_phv_out_last),
    .io_next_proc_exist(trans_10_io_next_proc_exist)
  );
  InterProcessorTransfer trans_11 ( // @[ipsa.scala 79:25]
    .clock(trans_11_clock),
    .io_pipe_phv_in_data_0(trans_11_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(trans_11_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(trans_11_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(trans_11_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(trans_11_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(trans_11_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(trans_11_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(trans_11_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(trans_11_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(trans_11_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(trans_11_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(trans_11_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(trans_11_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(trans_11_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(trans_11_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(trans_11_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(trans_11_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(trans_11_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(trans_11_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(trans_11_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(trans_11_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(trans_11_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(trans_11_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(trans_11_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(trans_11_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(trans_11_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(trans_11_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(trans_11_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(trans_11_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(trans_11_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(trans_11_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(trans_11_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(trans_11_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(trans_11_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(trans_11_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(trans_11_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(trans_11_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(trans_11_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(trans_11_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(trans_11_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(trans_11_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(trans_11_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(trans_11_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(trans_11_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(trans_11_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(trans_11_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(trans_11_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(trans_11_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(trans_11_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(trans_11_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(trans_11_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(trans_11_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(trans_11_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(trans_11_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(trans_11_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(trans_11_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(trans_11_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(trans_11_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(trans_11_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(trans_11_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(trans_11_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(trans_11_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(trans_11_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(trans_11_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(trans_11_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(trans_11_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(trans_11_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(trans_11_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(trans_11_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(trans_11_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(trans_11_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(trans_11_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(trans_11_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(trans_11_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(trans_11_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(trans_11_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(trans_11_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(trans_11_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(trans_11_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(trans_11_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(trans_11_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(trans_11_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(trans_11_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(trans_11_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(trans_11_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(trans_11_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(trans_11_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(trans_11_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(trans_11_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(trans_11_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(trans_11_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(trans_11_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(trans_11_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(trans_11_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(trans_11_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(trans_11_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(trans_11_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(trans_11_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(trans_11_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(trans_11_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(trans_11_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(trans_11_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(trans_11_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(trans_11_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(trans_11_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(trans_11_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(trans_11_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(trans_11_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(trans_11_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(trans_11_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(trans_11_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(trans_11_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(trans_11_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(trans_11_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(trans_11_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(trans_11_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(trans_11_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(trans_11_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(trans_11_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(trans_11_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(trans_11_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(trans_11_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(trans_11_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(trans_11_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(trans_11_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(trans_11_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(trans_11_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(trans_11_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(trans_11_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(trans_11_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(trans_11_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(trans_11_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(trans_11_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(trans_11_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(trans_11_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(trans_11_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(trans_11_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(trans_11_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(trans_11_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(trans_11_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(trans_11_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(trans_11_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(trans_11_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(trans_11_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(trans_11_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(trans_11_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(trans_11_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(trans_11_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(trans_11_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(trans_11_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(trans_11_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(trans_11_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(trans_11_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(trans_11_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(trans_11_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(trans_11_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(trans_11_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(trans_11_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(trans_11_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(trans_11_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_header_0(trans_11_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(trans_11_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(trans_11_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(trans_11_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(trans_11_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(trans_11_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(trans_11_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(trans_11_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(trans_11_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(trans_11_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(trans_11_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(trans_11_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(trans_11_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(trans_11_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(trans_11_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(trans_11_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(trans_11_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(trans_11_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(trans_11_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(trans_11_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(trans_11_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_valid(trans_11_io_pipe_phv_in_valid),
    .io_pipe_phv_in_last(trans_11_io_pipe_phv_in_last),
    .io_pipe_phv_out_data_0(trans_11_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(trans_11_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(trans_11_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(trans_11_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(trans_11_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(trans_11_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(trans_11_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(trans_11_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(trans_11_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(trans_11_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(trans_11_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(trans_11_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(trans_11_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(trans_11_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(trans_11_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(trans_11_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(trans_11_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(trans_11_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(trans_11_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(trans_11_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(trans_11_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(trans_11_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(trans_11_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(trans_11_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(trans_11_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(trans_11_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(trans_11_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(trans_11_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(trans_11_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(trans_11_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(trans_11_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(trans_11_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(trans_11_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(trans_11_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(trans_11_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(trans_11_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(trans_11_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(trans_11_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(trans_11_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(trans_11_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(trans_11_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(trans_11_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(trans_11_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(trans_11_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(trans_11_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(trans_11_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(trans_11_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(trans_11_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(trans_11_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(trans_11_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(trans_11_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(trans_11_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(trans_11_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(trans_11_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(trans_11_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(trans_11_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(trans_11_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(trans_11_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(trans_11_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(trans_11_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(trans_11_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(trans_11_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(trans_11_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(trans_11_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(trans_11_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(trans_11_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(trans_11_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(trans_11_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(trans_11_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(trans_11_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(trans_11_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(trans_11_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(trans_11_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(trans_11_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(trans_11_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(trans_11_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(trans_11_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(trans_11_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(trans_11_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(trans_11_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(trans_11_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(trans_11_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(trans_11_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(trans_11_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(trans_11_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(trans_11_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(trans_11_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(trans_11_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(trans_11_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(trans_11_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(trans_11_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(trans_11_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(trans_11_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(trans_11_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(trans_11_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(trans_11_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(trans_11_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(trans_11_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(trans_11_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(trans_11_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(trans_11_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(trans_11_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(trans_11_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(trans_11_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(trans_11_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(trans_11_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(trans_11_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(trans_11_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(trans_11_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(trans_11_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(trans_11_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(trans_11_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(trans_11_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(trans_11_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(trans_11_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(trans_11_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(trans_11_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(trans_11_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(trans_11_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(trans_11_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(trans_11_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(trans_11_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(trans_11_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(trans_11_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(trans_11_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(trans_11_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(trans_11_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(trans_11_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(trans_11_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(trans_11_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(trans_11_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(trans_11_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(trans_11_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(trans_11_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(trans_11_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(trans_11_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(trans_11_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(trans_11_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(trans_11_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(trans_11_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(trans_11_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(trans_11_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(trans_11_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(trans_11_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(trans_11_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(trans_11_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(trans_11_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(trans_11_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(trans_11_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(trans_11_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(trans_11_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(trans_11_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(trans_11_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(trans_11_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(trans_11_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(trans_11_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(trans_11_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(trans_11_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(trans_11_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(trans_11_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_header_0(trans_11_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(trans_11_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(trans_11_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(trans_11_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(trans_11_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(trans_11_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(trans_11_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(trans_11_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(trans_11_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(trans_11_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(trans_11_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(trans_11_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(trans_11_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(trans_11_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(trans_11_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(trans_11_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(trans_11_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(trans_11_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(trans_11_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(trans_11_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(trans_11_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(trans_11_io_pipe_phv_out_is_valid_processor),
    .io_pipe_phv_out_valid(trans_11_io_pipe_phv_out_valid),
    .io_pipe_phv_out_last(trans_11_io_pipe_phv_out_last),
    .io_next_proc_exist(trans_11_io_next_proc_exist)
  );
  InterProcessorTransfer trans_12 ( // @[ipsa.scala 79:25]
    .clock(trans_12_clock),
    .io_pipe_phv_in_data_0(trans_12_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(trans_12_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(trans_12_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(trans_12_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(trans_12_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(trans_12_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(trans_12_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(trans_12_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(trans_12_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(trans_12_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(trans_12_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(trans_12_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(trans_12_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(trans_12_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(trans_12_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(trans_12_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(trans_12_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(trans_12_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(trans_12_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(trans_12_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(trans_12_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(trans_12_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(trans_12_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(trans_12_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(trans_12_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(trans_12_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(trans_12_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(trans_12_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(trans_12_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(trans_12_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(trans_12_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(trans_12_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(trans_12_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(trans_12_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(trans_12_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(trans_12_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(trans_12_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(trans_12_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(trans_12_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(trans_12_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(trans_12_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(trans_12_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(trans_12_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(trans_12_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(trans_12_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(trans_12_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(trans_12_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(trans_12_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(trans_12_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(trans_12_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(trans_12_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(trans_12_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(trans_12_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(trans_12_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(trans_12_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(trans_12_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(trans_12_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(trans_12_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(trans_12_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(trans_12_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(trans_12_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(trans_12_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(trans_12_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(trans_12_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(trans_12_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(trans_12_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(trans_12_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(trans_12_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(trans_12_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(trans_12_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(trans_12_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(trans_12_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(trans_12_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(trans_12_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(trans_12_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(trans_12_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(trans_12_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(trans_12_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(trans_12_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(trans_12_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(trans_12_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(trans_12_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(trans_12_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(trans_12_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(trans_12_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(trans_12_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(trans_12_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(trans_12_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(trans_12_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(trans_12_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(trans_12_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(trans_12_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(trans_12_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(trans_12_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(trans_12_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(trans_12_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(trans_12_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(trans_12_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(trans_12_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(trans_12_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(trans_12_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(trans_12_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(trans_12_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(trans_12_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(trans_12_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(trans_12_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(trans_12_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(trans_12_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(trans_12_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(trans_12_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(trans_12_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(trans_12_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(trans_12_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(trans_12_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(trans_12_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(trans_12_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(trans_12_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(trans_12_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(trans_12_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(trans_12_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(trans_12_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(trans_12_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(trans_12_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(trans_12_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(trans_12_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(trans_12_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(trans_12_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(trans_12_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(trans_12_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(trans_12_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(trans_12_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(trans_12_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(trans_12_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(trans_12_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(trans_12_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(trans_12_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(trans_12_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(trans_12_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(trans_12_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(trans_12_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(trans_12_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(trans_12_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(trans_12_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(trans_12_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(trans_12_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(trans_12_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(trans_12_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(trans_12_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(trans_12_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(trans_12_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(trans_12_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(trans_12_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(trans_12_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(trans_12_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(trans_12_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(trans_12_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(trans_12_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(trans_12_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(trans_12_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(trans_12_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_header_0(trans_12_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(trans_12_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(trans_12_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(trans_12_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(trans_12_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(trans_12_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(trans_12_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(trans_12_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(trans_12_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(trans_12_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(trans_12_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(trans_12_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(trans_12_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(trans_12_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(trans_12_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(trans_12_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(trans_12_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(trans_12_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(trans_12_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(trans_12_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(trans_12_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_valid(trans_12_io_pipe_phv_in_valid),
    .io_pipe_phv_in_last(trans_12_io_pipe_phv_in_last),
    .io_pipe_phv_out_data_0(trans_12_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(trans_12_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(trans_12_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(trans_12_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(trans_12_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(trans_12_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(trans_12_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(trans_12_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(trans_12_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(trans_12_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(trans_12_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(trans_12_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(trans_12_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(trans_12_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(trans_12_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(trans_12_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(trans_12_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(trans_12_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(trans_12_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(trans_12_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(trans_12_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(trans_12_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(trans_12_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(trans_12_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(trans_12_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(trans_12_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(trans_12_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(trans_12_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(trans_12_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(trans_12_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(trans_12_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(trans_12_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(trans_12_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(trans_12_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(trans_12_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(trans_12_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(trans_12_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(trans_12_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(trans_12_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(trans_12_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(trans_12_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(trans_12_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(trans_12_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(trans_12_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(trans_12_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(trans_12_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(trans_12_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(trans_12_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(trans_12_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(trans_12_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(trans_12_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(trans_12_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(trans_12_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(trans_12_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(trans_12_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(trans_12_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(trans_12_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(trans_12_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(trans_12_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(trans_12_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(trans_12_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(trans_12_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(trans_12_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(trans_12_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(trans_12_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(trans_12_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(trans_12_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(trans_12_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(trans_12_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(trans_12_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(trans_12_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(trans_12_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(trans_12_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(trans_12_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(trans_12_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(trans_12_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(trans_12_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(trans_12_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(trans_12_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(trans_12_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(trans_12_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(trans_12_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(trans_12_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(trans_12_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(trans_12_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(trans_12_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(trans_12_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(trans_12_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(trans_12_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(trans_12_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(trans_12_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(trans_12_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(trans_12_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(trans_12_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(trans_12_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(trans_12_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(trans_12_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(trans_12_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(trans_12_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(trans_12_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(trans_12_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(trans_12_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(trans_12_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(trans_12_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(trans_12_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(trans_12_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(trans_12_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(trans_12_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(trans_12_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(trans_12_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(trans_12_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(trans_12_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(trans_12_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(trans_12_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(trans_12_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(trans_12_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(trans_12_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(trans_12_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(trans_12_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(trans_12_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(trans_12_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(trans_12_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(trans_12_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(trans_12_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(trans_12_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(trans_12_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(trans_12_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(trans_12_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(trans_12_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(trans_12_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(trans_12_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(trans_12_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(trans_12_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(trans_12_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(trans_12_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(trans_12_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(trans_12_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(trans_12_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(trans_12_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(trans_12_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(trans_12_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(trans_12_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(trans_12_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(trans_12_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(trans_12_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(trans_12_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(trans_12_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(trans_12_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(trans_12_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(trans_12_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(trans_12_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(trans_12_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(trans_12_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(trans_12_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(trans_12_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(trans_12_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(trans_12_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(trans_12_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(trans_12_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(trans_12_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_header_0(trans_12_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(trans_12_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(trans_12_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(trans_12_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(trans_12_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(trans_12_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(trans_12_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(trans_12_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(trans_12_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(trans_12_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(trans_12_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(trans_12_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(trans_12_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(trans_12_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(trans_12_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(trans_12_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(trans_12_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(trans_12_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(trans_12_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(trans_12_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(trans_12_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(trans_12_io_pipe_phv_out_is_valid_processor),
    .io_pipe_phv_out_valid(trans_12_io_pipe_phv_out_valid),
    .io_pipe_phv_out_last(trans_12_io_pipe_phv_out_last),
    .io_next_proc_exist(trans_12_io_next_proc_exist)
  );
  InterProcessorTransfer trans_13 ( // @[ipsa.scala 79:25]
    .clock(trans_13_clock),
    .io_pipe_phv_in_data_0(trans_13_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(trans_13_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(trans_13_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(trans_13_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(trans_13_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(trans_13_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(trans_13_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(trans_13_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(trans_13_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(trans_13_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(trans_13_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(trans_13_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(trans_13_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(trans_13_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(trans_13_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(trans_13_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(trans_13_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(trans_13_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(trans_13_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(trans_13_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(trans_13_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(trans_13_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(trans_13_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(trans_13_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(trans_13_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(trans_13_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(trans_13_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(trans_13_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(trans_13_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(trans_13_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(trans_13_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(trans_13_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(trans_13_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(trans_13_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(trans_13_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(trans_13_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(trans_13_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(trans_13_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(trans_13_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(trans_13_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(trans_13_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(trans_13_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(trans_13_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(trans_13_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(trans_13_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(trans_13_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(trans_13_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(trans_13_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(trans_13_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(trans_13_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(trans_13_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(trans_13_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(trans_13_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(trans_13_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(trans_13_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(trans_13_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(trans_13_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(trans_13_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(trans_13_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(trans_13_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(trans_13_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(trans_13_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(trans_13_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(trans_13_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(trans_13_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(trans_13_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(trans_13_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(trans_13_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(trans_13_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(trans_13_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(trans_13_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(trans_13_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(trans_13_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(trans_13_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(trans_13_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(trans_13_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(trans_13_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(trans_13_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(trans_13_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(trans_13_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(trans_13_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(trans_13_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(trans_13_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(trans_13_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(trans_13_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(trans_13_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(trans_13_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(trans_13_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(trans_13_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(trans_13_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(trans_13_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(trans_13_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(trans_13_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(trans_13_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(trans_13_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(trans_13_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(trans_13_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(trans_13_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(trans_13_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(trans_13_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(trans_13_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(trans_13_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(trans_13_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(trans_13_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(trans_13_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(trans_13_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(trans_13_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(trans_13_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(trans_13_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(trans_13_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(trans_13_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(trans_13_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(trans_13_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(trans_13_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(trans_13_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(trans_13_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(trans_13_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(trans_13_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(trans_13_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(trans_13_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(trans_13_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(trans_13_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(trans_13_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(trans_13_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(trans_13_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(trans_13_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(trans_13_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(trans_13_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(trans_13_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(trans_13_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(trans_13_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(trans_13_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(trans_13_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(trans_13_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(trans_13_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(trans_13_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(trans_13_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(trans_13_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(trans_13_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(trans_13_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(trans_13_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(trans_13_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(trans_13_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(trans_13_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(trans_13_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(trans_13_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(trans_13_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(trans_13_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(trans_13_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(trans_13_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(trans_13_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(trans_13_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(trans_13_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(trans_13_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(trans_13_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(trans_13_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(trans_13_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(trans_13_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(trans_13_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(trans_13_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_header_0(trans_13_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(trans_13_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(trans_13_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(trans_13_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(trans_13_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(trans_13_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(trans_13_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(trans_13_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(trans_13_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(trans_13_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(trans_13_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(trans_13_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(trans_13_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(trans_13_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(trans_13_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(trans_13_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(trans_13_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(trans_13_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(trans_13_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(trans_13_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(trans_13_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_valid(trans_13_io_pipe_phv_in_valid),
    .io_pipe_phv_in_last(trans_13_io_pipe_phv_in_last),
    .io_pipe_phv_out_data_0(trans_13_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(trans_13_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(trans_13_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(trans_13_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(trans_13_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(trans_13_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(trans_13_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(trans_13_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(trans_13_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(trans_13_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(trans_13_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(trans_13_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(trans_13_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(trans_13_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(trans_13_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(trans_13_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(trans_13_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(trans_13_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(trans_13_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(trans_13_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(trans_13_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(trans_13_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(trans_13_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(trans_13_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(trans_13_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(trans_13_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(trans_13_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(trans_13_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(trans_13_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(trans_13_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(trans_13_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(trans_13_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(trans_13_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(trans_13_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(trans_13_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(trans_13_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(trans_13_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(trans_13_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(trans_13_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(trans_13_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(trans_13_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(trans_13_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(trans_13_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(trans_13_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(trans_13_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(trans_13_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(trans_13_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(trans_13_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(trans_13_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(trans_13_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(trans_13_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(trans_13_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(trans_13_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(trans_13_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(trans_13_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(trans_13_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(trans_13_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(trans_13_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(trans_13_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(trans_13_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(trans_13_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(trans_13_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(trans_13_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(trans_13_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(trans_13_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(trans_13_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(trans_13_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(trans_13_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(trans_13_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(trans_13_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(trans_13_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(trans_13_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(trans_13_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(trans_13_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(trans_13_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(trans_13_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(trans_13_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(trans_13_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(trans_13_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(trans_13_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(trans_13_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(trans_13_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(trans_13_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(trans_13_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(trans_13_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(trans_13_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(trans_13_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(trans_13_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(trans_13_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(trans_13_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(trans_13_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(trans_13_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(trans_13_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(trans_13_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(trans_13_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(trans_13_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(trans_13_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(trans_13_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(trans_13_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(trans_13_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(trans_13_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(trans_13_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(trans_13_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(trans_13_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(trans_13_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(trans_13_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(trans_13_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(trans_13_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(trans_13_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(trans_13_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(trans_13_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(trans_13_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(trans_13_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(trans_13_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(trans_13_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(trans_13_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(trans_13_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(trans_13_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(trans_13_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(trans_13_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(trans_13_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(trans_13_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(trans_13_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(trans_13_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(trans_13_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(trans_13_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(trans_13_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(trans_13_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(trans_13_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(trans_13_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(trans_13_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(trans_13_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(trans_13_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(trans_13_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(trans_13_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(trans_13_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(trans_13_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(trans_13_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(trans_13_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(trans_13_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(trans_13_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(trans_13_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(trans_13_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(trans_13_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(trans_13_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(trans_13_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(trans_13_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(trans_13_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(trans_13_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(trans_13_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(trans_13_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(trans_13_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(trans_13_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(trans_13_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(trans_13_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(trans_13_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(trans_13_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(trans_13_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(trans_13_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(trans_13_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_header_0(trans_13_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(trans_13_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(trans_13_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(trans_13_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(trans_13_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(trans_13_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(trans_13_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(trans_13_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(trans_13_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(trans_13_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(trans_13_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(trans_13_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(trans_13_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(trans_13_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(trans_13_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(trans_13_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(trans_13_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(trans_13_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(trans_13_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(trans_13_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(trans_13_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(trans_13_io_pipe_phv_out_is_valid_processor),
    .io_pipe_phv_out_valid(trans_13_io_pipe_phv_out_valid),
    .io_pipe_phv_out_last(trans_13_io_pipe_phv_out_last),
    .io_next_proc_exist(trans_13_io_next_proc_exist)
  );
  InterProcessorTransfer trans_14 ( // @[ipsa.scala 79:25]
    .clock(trans_14_clock),
    .io_pipe_phv_in_data_0(trans_14_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(trans_14_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(trans_14_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(trans_14_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(trans_14_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(trans_14_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(trans_14_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(trans_14_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(trans_14_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(trans_14_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(trans_14_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(trans_14_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(trans_14_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(trans_14_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(trans_14_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(trans_14_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(trans_14_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(trans_14_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(trans_14_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(trans_14_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(trans_14_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(trans_14_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(trans_14_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(trans_14_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(trans_14_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(trans_14_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(trans_14_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(trans_14_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(trans_14_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(trans_14_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(trans_14_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(trans_14_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(trans_14_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(trans_14_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(trans_14_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(trans_14_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(trans_14_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(trans_14_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(trans_14_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(trans_14_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(trans_14_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(trans_14_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(trans_14_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(trans_14_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(trans_14_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(trans_14_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(trans_14_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(trans_14_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(trans_14_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(trans_14_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(trans_14_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(trans_14_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(trans_14_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(trans_14_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(trans_14_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(trans_14_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(trans_14_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(trans_14_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(trans_14_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(trans_14_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(trans_14_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(trans_14_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(trans_14_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(trans_14_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(trans_14_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(trans_14_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(trans_14_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(trans_14_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(trans_14_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(trans_14_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(trans_14_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(trans_14_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(trans_14_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(trans_14_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(trans_14_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(trans_14_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(trans_14_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(trans_14_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(trans_14_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(trans_14_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(trans_14_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(trans_14_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(trans_14_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(trans_14_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(trans_14_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(trans_14_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(trans_14_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(trans_14_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(trans_14_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(trans_14_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(trans_14_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(trans_14_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(trans_14_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(trans_14_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(trans_14_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(trans_14_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(trans_14_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(trans_14_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(trans_14_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(trans_14_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(trans_14_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(trans_14_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(trans_14_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(trans_14_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(trans_14_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(trans_14_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(trans_14_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(trans_14_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(trans_14_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(trans_14_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(trans_14_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(trans_14_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(trans_14_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(trans_14_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(trans_14_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(trans_14_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(trans_14_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(trans_14_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(trans_14_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(trans_14_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(trans_14_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(trans_14_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(trans_14_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(trans_14_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(trans_14_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(trans_14_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(trans_14_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(trans_14_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(trans_14_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(trans_14_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(trans_14_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(trans_14_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(trans_14_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(trans_14_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(trans_14_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(trans_14_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(trans_14_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(trans_14_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(trans_14_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(trans_14_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(trans_14_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(trans_14_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(trans_14_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(trans_14_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(trans_14_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(trans_14_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(trans_14_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(trans_14_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(trans_14_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(trans_14_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(trans_14_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(trans_14_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(trans_14_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(trans_14_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(trans_14_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(trans_14_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(trans_14_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(trans_14_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(trans_14_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(trans_14_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_header_0(trans_14_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(trans_14_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(trans_14_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(trans_14_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(trans_14_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(trans_14_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(trans_14_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(trans_14_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(trans_14_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(trans_14_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(trans_14_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(trans_14_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(trans_14_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(trans_14_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(trans_14_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(trans_14_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(trans_14_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(trans_14_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(trans_14_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(trans_14_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(trans_14_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_valid(trans_14_io_pipe_phv_in_valid),
    .io_pipe_phv_in_last(trans_14_io_pipe_phv_in_last),
    .io_pipe_phv_out_data_0(trans_14_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(trans_14_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(trans_14_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(trans_14_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(trans_14_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(trans_14_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(trans_14_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(trans_14_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(trans_14_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(trans_14_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(trans_14_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(trans_14_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(trans_14_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(trans_14_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(trans_14_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(trans_14_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(trans_14_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(trans_14_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(trans_14_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(trans_14_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(trans_14_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(trans_14_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(trans_14_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(trans_14_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(trans_14_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(trans_14_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(trans_14_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(trans_14_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(trans_14_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(trans_14_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(trans_14_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(trans_14_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(trans_14_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(trans_14_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(trans_14_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(trans_14_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(trans_14_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(trans_14_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(trans_14_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(trans_14_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(trans_14_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(trans_14_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(trans_14_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(trans_14_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(trans_14_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(trans_14_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(trans_14_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(trans_14_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(trans_14_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(trans_14_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(trans_14_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(trans_14_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(trans_14_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(trans_14_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(trans_14_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(trans_14_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(trans_14_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(trans_14_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(trans_14_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(trans_14_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(trans_14_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(trans_14_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(trans_14_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(trans_14_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(trans_14_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(trans_14_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(trans_14_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(trans_14_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(trans_14_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(trans_14_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(trans_14_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(trans_14_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(trans_14_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(trans_14_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(trans_14_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(trans_14_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(trans_14_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(trans_14_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(trans_14_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(trans_14_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(trans_14_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(trans_14_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(trans_14_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(trans_14_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(trans_14_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(trans_14_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(trans_14_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(trans_14_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(trans_14_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(trans_14_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(trans_14_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(trans_14_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(trans_14_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(trans_14_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(trans_14_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(trans_14_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(trans_14_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(trans_14_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(trans_14_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(trans_14_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(trans_14_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(trans_14_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(trans_14_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(trans_14_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(trans_14_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(trans_14_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(trans_14_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(trans_14_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(trans_14_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(trans_14_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(trans_14_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(trans_14_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(trans_14_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(trans_14_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(trans_14_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(trans_14_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(trans_14_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(trans_14_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(trans_14_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(trans_14_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(trans_14_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(trans_14_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(trans_14_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(trans_14_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(trans_14_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(trans_14_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(trans_14_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(trans_14_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(trans_14_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(trans_14_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(trans_14_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(trans_14_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(trans_14_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(trans_14_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(trans_14_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(trans_14_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(trans_14_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(trans_14_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(trans_14_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(trans_14_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(trans_14_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(trans_14_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(trans_14_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(trans_14_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(trans_14_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(trans_14_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(trans_14_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(trans_14_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(trans_14_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(trans_14_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(trans_14_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(trans_14_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(trans_14_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(trans_14_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(trans_14_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(trans_14_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(trans_14_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(trans_14_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(trans_14_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(trans_14_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_header_0(trans_14_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(trans_14_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(trans_14_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(trans_14_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(trans_14_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(trans_14_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(trans_14_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(trans_14_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(trans_14_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(trans_14_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(trans_14_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(trans_14_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(trans_14_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(trans_14_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(trans_14_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(trans_14_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(trans_14_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(trans_14_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(trans_14_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(trans_14_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(trans_14_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(trans_14_io_pipe_phv_out_is_valid_processor),
    .io_pipe_phv_out_valid(trans_14_io_pipe_phv_out_valid),
    .io_pipe_phv_out_last(trans_14_io_pipe_phv_out_last),
    .io_next_proc_exist(trans_14_io_next_proc_exist)
  );
  InterProcessorTransfer trans_15 ( // @[ipsa.scala 79:25]
    .clock(trans_15_clock),
    .io_pipe_phv_in_data_0(trans_15_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(trans_15_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(trans_15_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(trans_15_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(trans_15_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(trans_15_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(trans_15_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(trans_15_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(trans_15_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(trans_15_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(trans_15_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(trans_15_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(trans_15_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(trans_15_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(trans_15_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(trans_15_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(trans_15_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(trans_15_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(trans_15_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(trans_15_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(trans_15_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(trans_15_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(trans_15_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(trans_15_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(trans_15_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(trans_15_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(trans_15_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(trans_15_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(trans_15_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(trans_15_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(trans_15_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(trans_15_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(trans_15_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(trans_15_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(trans_15_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(trans_15_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(trans_15_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(trans_15_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(trans_15_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(trans_15_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(trans_15_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(trans_15_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(trans_15_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(trans_15_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(trans_15_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(trans_15_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(trans_15_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(trans_15_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(trans_15_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(trans_15_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(trans_15_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(trans_15_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(trans_15_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(trans_15_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(trans_15_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(trans_15_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(trans_15_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(trans_15_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(trans_15_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(trans_15_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(trans_15_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(trans_15_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(trans_15_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(trans_15_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(trans_15_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(trans_15_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(trans_15_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(trans_15_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(trans_15_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(trans_15_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(trans_15_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(trans_15_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(trans_15_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(trans_15_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(trans_15_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(trans_15_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(trans_15_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(trans_15_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(trans_15_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(trans_15_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(trans_15_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(trans_15_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(trans_15_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(trans_15_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(trans_15_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(trans_15_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(trans_15_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(trans_15_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(trans_15_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(trans_15_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(trans_15_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(trans_15_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(trans_15_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(trans_15_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(trans_15_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(trans_15_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(trans_15_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(trans_15_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(trans_15_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(trans_15_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(trans_15_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(trans_15_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(trans_15_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(trans_15_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(trans_15_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(trans_15_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(trans_15_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(trans_15_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(trans_15_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(trans_15_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(trans_15_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(trans_15_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(trans_15_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(trans_15_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(trans_15_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(trans_15_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(trans_15_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(trans_15_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(trans_15_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(trans_15_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(trans_15_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(trans_15_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(trans_15_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(trans_15_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(trans_15_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(trans_15_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(trans_15_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(trans_15_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(trans_15_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(trans_15_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(trans_15_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(trans_15_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(trans_15_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(trans_15_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(trans_15_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(trans_15_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(trans_15_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(trans_15_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(trans_15_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(trans_15_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(trans_15_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(trans_15_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(trans_15_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(trans_15_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(trans_15_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(trans_15_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(trans_15_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(trans_15_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(trans_15_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(trans_15_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(trans_15_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(trans_15_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(trans_15_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(trans_15_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(trans_15_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(trans_15_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(trans_15_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(trans_15_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(trans_15_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(trans_15_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_header_0(trans_15_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(trans_15_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(trans_15_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(trans_15_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(trans_15_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(trans_15_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(trans_15_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(trans_15_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(trans_15_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(trans_15_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(trans_15_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(trans_15_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(trans_15_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(trans_15_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(trans_15_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(trans_15_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(trans_15_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(trans_15_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(trans_15_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(trans_15_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(trans_15_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_valid(trans_15_io_pipe_phv_in_valid),
    .io_pipe_phv_in_last(trans_15_io_pipe_phv_in_last),
    .io_pipe_phv_out_data_0(trans_15_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(trans_15_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(trans_15_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(trans_15_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(trans_15_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(trans_15_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(trans_15_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(trans_15_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(trans_15_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(trans_15_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(trans_15_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(trans_15_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(trans_15_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(trans_15_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(trans_15_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(trans_15_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(trans_15_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(trans_15_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(trans_15_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(trans_15_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(trans_15_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(trans_15_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(trans_15_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(trans_15_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(trans_15_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(trans_15_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(trans_15_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(trans_15_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(trans_15_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(trans_15_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(trans_15_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(trans_15_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(trans_15_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(trans_15_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(trans_15_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(trans_15_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(trans_15_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(trans_15_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(trans_15_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(trans_15_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(trans_15_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(trans_15_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(trans_15_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(trans_15_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(trans_15_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(trans_15_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(trans_15_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(trans_15_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(trans_15_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(trans_15_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(trans_15_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(trans_15_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(trans_15_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(trans_15_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(trans_15_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(trans_15_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(trans_15_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(trans_15_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(trans_15_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(trans_15_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(trans_15_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(trans_15_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(trans_15_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(trans_15_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(trans_15_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(trans_15_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(trans_15_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(trans_15_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(trans_15_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(trans_15_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(trans_15_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(trans_15_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(trans_15_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(trans_15_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(trans_15_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(trans_15_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(trans_15_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(trans_15_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(trans_15_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(trans_15_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(trans_15_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(trans_15_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(trans_15_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(trans_15_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(trans_15_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(trans_15_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(trans_15_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(trans_15_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(trans_15_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(trans_15_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(trans_15_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(trans_15_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(trans_15_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(trans_15_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(trans_15_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(trans_15_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(trans_15_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(trans_15_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(trans_15_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(trans_15_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(trans_15_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(trans_15_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(trans_15_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(trans_15_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(trans_15_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(trans_15_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(trans_15_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(trans_15_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(trans_15_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(trans_15_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(trans_15_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(trans_15_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(trans_15_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(trans_15_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(trans_15_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(trans_15_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(trans_15_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(trans_15_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(trans_15_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(trans_15_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(trans_15_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(trans_15_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(trans_15_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(trans_15_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(trans_15_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(trans_15_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(trans_15_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(trans_15_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(trans_15_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(trans_15_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(trans_15_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(trans_15_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(trans_15_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(trans_15_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(trans_15_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(trans_15_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(trans_15_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(trans_15_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(trans_15_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(trans_15_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(trans_15_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(trans_15_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(trans_15_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(trans_15_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(trans_15_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(trans_15_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(trans_15_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(trans_15_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(trans_15_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(trans_15_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(trans_15_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(trans_15_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(trans_15_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(trans_15_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(trans_15_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(trans_15_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(trans_15_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(trans_15_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(trans_15_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(trans_15_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_header_0(trans_15_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(trans_15_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(trans_15_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(trans_15_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(trans_15_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(trans_15_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(trans_15_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(trans_15_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(trans_15_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(trans_15_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(trans_15_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(trans_15_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(trans_15_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(trans_15_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(trans_15_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(trans_15_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(trans_15_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(trans_15_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(trans_15_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(trans_15_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(trans_15_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(trans_15_io_pipe_phv_out_is_valid_processor),
    .io_pipe_phv_out_valid(trans_15_io_pipe_phv_out_valid),
    .io_pipe_phv_out_last(trans_15_io_pipe_phv_out_last),
    .io_next_proc_exist(trans_15_io_next_proc_exist)
  );
  assign io_pipe_phv_out_data_0 = trans_0_io_pipe_phv_out_data_0; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_1 = trans_0_io_pipe_phv_out_data_1; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_2 = trans_0_io_pipe_phv_out_data_2; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_3 = trans_0_io_pipe_phv_out_data_3; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_4 = trans_0_io_pipe_phv_out_data_4; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_5 = trans_0_io_pipe_phv_out_data_5; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_6 = trans_0_io_pipe_phv_out_data_6; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_7 = trans_0_io_pipe_phv_out_data_7; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_8 = trans_0_io_pipe_phv_out_data_8; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_9 = trans_0_io_pipe_phv_out_data_9; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_10 = trans_0_io_pipe_phv_out_data_10; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_11 = trans_0_io_pipe_phv_out_data_11; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_12 = trans_0_io_pipe_phv_out_data_12; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_13 = trans_0_io_pipe_phv_out_data_13; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_14 = trans_0_io_pipe_phv_out_data_14; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_15 = trans_0_io_pipe_phv_out_data_15; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_16 = trans_0_io_pipe_phv_out_data_16; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_17 = trans_0_io_pipe_phv_out_data_17; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_18 = trans_0_io_pipe_phv_out_data_18; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_19 = trans_0_io_pipe_phv_out_data_19; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_20 = trans_0_io_pipe_phv_out_data_20; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_21 = trans_0_io_pipe_phv_out_data_21; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_22 = trans_0_io_pipe_phv_out_data_22; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_23 = trans_0_io_pipe_phv_out_data_23; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_24 = trans_0_io_pipe_phv_out_data_24; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_25 = trans_0_io_pipe_phv_out_data_25; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_26 = trans_0_io_pipe_phv_out_data_26; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_27 = trans_0_io_pipe_phv_out_data_27; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_28 = trans_0_io_pipe_phv_out_data_28; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_29 = trans_0_io_pipe_phv_out_data_29; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_30 = trans_0_io_pipe_phv_out_data_30; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_31 = trans_0_io_pipe_phv_out_data_31; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_32 = trans_0_io_pipe_phv_out_data_32; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_33 = trans_0_io_pipe_phv_out_data_33; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_34 = trans_0_io_pipe_phv_out_data_34; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_35 = trans_0_io_pipe_phv_out_data_35; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_36 = trans_0_io_pipe_phv_out_data_36; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_37 = trans_0_io_pipe_phv_out_data_37; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_38 = trans_0_io_pipe_phv_out_data_38; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_39 = trans_0_io_pipe_phv_out_data_39; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_40 = trans_0_io_pipe_phv_out_data_40; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_41 = trans_0_io_pipe_phv_out_data_41; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_42 = trans_0_io_pipe_phv_out_data_42; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_43 = trans_0_io_pipe_phv_out_data_43; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_44 = trans_0_io_pipe_phv_out_data_44; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_45 = trans_0_io_pipe_phv_out_data_45; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_46 = trans_0_io_pipe_phv_out_data_46; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_47 = trans_0_io_pipe_phv_out_data_47; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_48 = trans_0_io_pipe_phv_out_data_48; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_49 = trans_0_io_pipe_phv_out_data_49; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_50 = trans_0_io_pipe_phv_out_data_50; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_51 = trans_0_io_pipe_phv_out_data_51; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_52 = trans_0_io_pipe_phv_out_data_52; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_53 = trans_0_io_pipe_phv_out_data_53; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_54 = trans_0_io_pipe_phv_out_data_54; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_55 = trans_0_io_pipe_phv_out_data_55; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_56 = trans_0_io_pipe_phv_out_data_56; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_57 = trans_0_io_pipe_phv_out_data_57; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_58 = trans_0_io_pipe_phv_out_data_58; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_59 = trans_0_io_pipe_phv_out_data_59; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_60 = trans_0_io_pipe_phv_out_data_60; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_61 = trans_0_io_pipe_phv_out_data_61; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_62 = trans_0_io_pipe_phv_out_data_62; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_63 = trans_0_io_pipe_phv_out_data_63; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_64 = trans_0_io_pipe_phv_out_data_64; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_65 = trans_0_io_pipe_phv_out_data_65; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_66 = trans_0_io_pipe_phv_out_data_66; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_67 = trans_0_io_pipe_phv_out_data_67; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_68 = trans_0_io_pipe_phv_out_data_68; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_69 = trans_0_io_pipe_phv_out_data_69; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_70 = trans_0_io_pipe_phv_out_data_70; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_71 = trans_0_io_pipe_phv_out_data_71; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_72 = trans_0_io_pipe_phv_out_data_72; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_73 = trans_0_io_pipe_phv_out_data_73; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_74 = trans_0_io_pipe_phv_out_data_74; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_75 = trans_0_io_pipe_phv_out_data_75; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_76 = trans_0_io_pipe_phv_out_data_76; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_77 = trans_0_io_pipe_phv_out_data_77; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_78 = trans_0_io_pipe_phv_out_data_78; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_79 = trans_0_io_pipe_phv_out_data_79; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_80 = trans_0_io_pipe_phv_out_data_80; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_81 = trans_0_io_pipe_phv_out_data_81; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_82 = trans_0_io_pipe_phv_out_data_82; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_83 = trans_0_io_pipe_phv_out_data_83; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_84 = trans_0_io_pipe_phv_out_data_84; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_85 = trans_0_io_pipe_phv_out_data_85; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_86 = trans_0_io_pipe_phv_out_data_86; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_87 = trans_0_io_pipe_phv_out_data_87; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_88 = trans_0_io_pipe_phv_out_data_88; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_89 = trans_0_io_pipe_phv_out_data_89; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_90 = trans_0_io_pipe_phv_out_data_90; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_91 = trans_0_io_pipe_phv_out_data_91; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_92 = trans_0_io_pipe_phv_out_data_92; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_93 = trans_0_io_pipe_phv_out_data_93; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_94 = trans_0_io_pipe_phv_out_data_94; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_95 = trans_0_io_pipe_phv_out_data_95; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_96 = trans_0_io_pipe_phv_out_data_96; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_97 = trans_0_io_pipe_phv_out_data_97; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_98 = trans_0_io_pipe_phv_out_data_98; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_99 = trans_0_io_pipe_phv_out_data_99; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_100 = trans_0_io_pipe_phv_out_data_100; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_101 = trans_0_io_pipe_phv_out_data_101; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_102 = trans_0_io_pipe_phv_out_data_102; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_103 = trans_0_io_pipe_phv_out_data_103; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_104 = trans_0_io_pipe_phv_out_data_104; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_105 = trans_0_io_pipe_phv_out_data_105; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_106 = trans_0_io_pipe_phv_out_data_106; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_107 = trans_0_io_pipe_phv_out_data_107; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_108 = trans_0_io_pipe_phv_out_data_108; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_109 = trans_0_io_pipe_phv_out_data_109; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_110 = trans_0_io_pipe_phv_out_data_110; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_111 = trans_0_io_pipe_phv_out_data_111; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_112 = trans_0_io_pipe_phv_out_data_112; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_113 = trans_0_io_pipe_phv_out_data_113; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_114 = trans_0_io_pipe_phv_out_data_114; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_115 = trans_0_io_pipe_phv_out_data_115; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_116 = trans_0_io_pipe_phv_out_data_116; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_117 = trans_0_io_pipe_phv_out_data_117; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_118 = trans_0_io_pipe_phv_out_data_118; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_119 = trans_0_io_pipe_phv_out_data_119; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_120 = trans_0_io_pipe_phv_out_data_120; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_121 = trans_0_io_pipe_phv_out_data_121; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_122 = trans_0_io_pipe_phv_out_data_122; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_123 = trans_0_io_pipe_phv_out_data_123; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_124 = trans_0_io_pipe_phv_out_data_124; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_125 = trans_0_io_pipe_phv_out_data_125; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_126 = trans_0_io_pipe_phv_out_data_126; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_127 = trans_0_io_pipe_phv_out_data_127; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_valid = trans_0_io_pipe_phv_out_valid; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign io_pipe_phv_out_last = trans_0_io_pipe_phv_out_last; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  assign proc_0_clock = clock;
  assign proc_0_io_pipe_phv_in_data_0 = trans_15_io_pipe_phv_out_data_0; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_1 = trans_15_io_pipe_phv_out_data_1; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_2 = trans_15_io_pipe_phv_out_data_2; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_3 = trans_15_io_pipe_phv_out_data_3; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_4 = trans_15_io_pipe_phv_out_data_4; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_5 = trans_15_io_pipe_phv_out_data_5; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_6 = trans_15_io_pipe_phv_out_data_6; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_7 = trans_15_io_pipe_phv_out_data_7; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_8 = trans_15_io_pipe_phv_out_data_8; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_9 = trans_15_io_pipe_phv_out_data_9; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_10 = trans_15_io_pipe_phv_out_data_10; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_11 = trans_15_io_pipe_phv_out_data_11; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_12 = trans_15_io_pipe_phv_out_data_12; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_13 = trans_15_io_pipe_phv_out_data_13; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_14 = trans_15_io_pipe_phv_out_data_14; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_15 = trans_15_io_pipe_phv_out_data_15; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_16 = trans_15_io_pipe_phv_out_data_16; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_17 = trans_15_io_pipe_phv_out_data_17; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_18 = trans_15_io_pipe_phv_out_data_18; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_19 = trans_15_io_pipe_phv_out_data_19; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_20 = trans_15_io_pipe_phv_out_data_20; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_21 = trans_15_io_pipe_phv_out_data_21; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_22 = trans_15_io_pipe_phv_out_data_22; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_23 = trans_15_io_pipe_phv_out_data_23; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_24 = trans_15_io_pipe_phv_out_data_24; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_25 = trans_15_io_pipe_phv_out_data_25; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_26 = trans_15_io_pipe_phv_out_data_26; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_27 = trans_15_io_pipe_phv_out_data_27; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_28 = trans_15_io_pipe_phv_out_data_28; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_29 = trans_15_io_pipe_phv_out_data_29; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_30 = trans_15_io_pipe_phv_out_data_30; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_31 = trans_15_io_pipe_phv_out_data_31; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_32 = trans_15_io_pipe_phv_out_data_32; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_33 = trans_15_io_pipe_phv_out_data_33; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_34 = trans_15_io_pipe_phv_out_data_34; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_35 = trans_15_io_pipe_phv_out_data_35; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_36 = trans_15_io_pipe_phv_out_data_36; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_37 = trans_15_io_pipe_phv_out_data_37; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_38 = trans_15_io_pipe_phv_out_data_38; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_39 = trans_15_io_pipe_phv_out_data_39; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_40 = trans_15_io_pipe_phv_out_data_40; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_41 = trans_15_io_pipe_phv_out_data_41; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_42 = trans_15_io_pipe_phv_out_data_42; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_43 = trans_15_io_pipe_phv_out_data_43; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_44 = trans_15_io_pipe_phv_out_data_44; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_45 = trans_15_io_pipe_phv_out_data_45; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_46 = trans_15_io_pipe_phv_out_data_46; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_47 = trans_15_io_pipe_phv_out_data_47; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_48 = trans_15_io_pipe_phv_out_data_48; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_49 = trans_15_io_pipe_phv_out_data_49; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_50 = trans_15_io_pipe_phv_out_data_50; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_51 = trans_15_io_pipe_phv_out_data_51; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_52 = trans_15_io_pipe_phv_out_data_52; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_53 = trans_15_io_pipe_phv_out_data_53; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_54 = trans_15_io_pipe_phv_out_data_54; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_55 = trans_15_io_pipe_phv_out_data_55; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_56 = trans_15_io_pipe_phv_out_data_56; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_57 = trans_15_io_pipe_phv_out_data_57; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_58 = trans_15_io_pipe_phv_out_data_58; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_59 = trans_15_io_pipe_phv_out_data_59; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_60 = trans_15_io_pipe_phv_out_data_60; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_61 = trans_15_io_pipe_phv_out_data_61; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_62 = trans_15_io_pipe_phv_out_data_62; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_63 = trans_15_io_pipe_phv_out_data_63; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_64 = trans_15_io_pipe_phv_out_data_64; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_65 = trans_15_io_pipe_phv_out_data_65; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_66 = trans_15_io_pipe_phv_out_data_66; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_67 = trans_15_io_pipe_phv_out_data_67; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_68 = trans_15_io_pipe_phv_out_data_68; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_69 = trans_15_io_pipe_phv_out_data_69; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_70 = trans_15_io_pipe_phv_out_data_70; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_71 = trans_15_io_pipe_phv_out_data_71; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_72 = trans_15_io_pipe_phv_out_data_72; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_73 = trans_15_io_pipe_phv_out_data_73; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_74 = trans_15_io_pipe_phv_out_data_74; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_75 = trans_15_io_pipe_phv_out_data_75; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_76 = trans_15_io_pipe_phv_out_data_76; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_77 = trans_15_io_pipe_phv_out_data_77; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_78 = trans_15_io_pipe_phv_out_data_78; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_79 = trans_15_io_pipe_phv_out_data_79; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_80 = trans_15_io_pipe_phv_out_data_80; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_81 = trans_15_io_pipe_phv_out_data_81; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_82 = trans_15_io_pipe_phv_out_data_82; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_83 = trans_15_io_pipe_phv_out_data_83; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_84 = trans_15_io_pipe_phv_out_data_84; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_85 = trans_15_io_pipe_phv_out_data_85; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_86 = trans_15_io_pipe_phv_out_data_86; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_87 = trans_15_io_pipe_phv_out_data_87; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_88 = trans_15_io_pipe_phv_out_data_88; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_89 = trans_15_io_pipe_phv_out_data_89; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_90 = trans_15_io_pipe_phv_out_data_90; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_91 = trans_15_io_pipe_phv_out_data_91; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_92 = trans_15_io_pipe_phv_out_data_92; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_93 = trans_15_io_pipe_phv_out_data_93; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_94 = trans_15_io_pipe_phv_out_data_94; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_95 = trans_15_io_pipe_phv_out_data_95; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_96 = trans_15_io_pipe_phv_out_data_96; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_97 = trans_15_io_pipe_phv_out_data_97; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_98 = trans_15_io_pipe_phv_out_data_98; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_99 = trans_15_io_pipe_phv_out_data_99; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_100 = trans_15_io_pipe_phv_out_data_100; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_101 = trans_15_io_pipe_phv_out_data_101; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_102 = trans_15_io_pipe_phv_out_data_102; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_103 = trans_15_io_pipe_phv_out_data_103; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_104 = trans_15_io_pipe_phv_out_data_104; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_105 = trans_15_io_pipe_phv_out_data_105; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_106 = trans_15_io_pipe_phv_out_data_106; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_107 = trans_15_io_pipe_phv_out_data_107; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_108 = trans_15_io_pipe_phv_out_data_108; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_109 = trans_15_io_pipe_phv_out_data_109; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_110 = trans_15_io_pipe_phv_out_data_110; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_111 = trans_15_io_pipe_phv_out_data_111; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_112 = trans_15_io_pipe_phv_out_data_112; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_113 = trans_15_io_pipe_phv_out_data_113; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_114 = trans_15_io_pipe_phv_out_data_114; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_115 = trans_15_io_pipe_phv_out_data_115; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_116 = trans_15_io_pipe_phv_out_data_116; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_117 = trans_15_io_pipe_phv_out_data_117; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_118 = trans_15_io_pipe_phv_out_data_118; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_119 = trans_15_io_pipe_phv_out_data_119; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_120 = trans_15_io_pipe_phv_out_data_120; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_121 = trans_15_io_pipe_phv_out_data_121; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_122 = trans_15_io_pipe_phv_out_data_122; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_123 = trans_15_io_pipe_phv_out_data_123; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_124 = trans_15_io_pipe_phv_out_data_124; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_125 = trans_15_io_pipe_phv_out_data_125; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_126 = trans_15_io_pipe_phv_out_data_126; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_127 = trans_15_io_pipe_phv_out_data_127; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_128 = trans_15_io_pipe_phv_out_data_128; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_129 = trans_15_io_pipe_phv_out_data_129; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_130 = trans_15_io_pipe_phv_out_data_130; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_131 = trans_15_io_pipe_phv_out_data_131; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_132 = trans_15_io_pipe_phv_out_data_132; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_133 = trans_15_io_pipe_phv_out_data_133; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_134 = trans_15_io_pipe_phv_out_data_134; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_135 = trans_15_io_pipe_phv_out_data_135; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_136 = trans_15_io_pipe_phv_out_data_136; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_137 = trans_15_io_pipe_phv_out_data_137; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_138 = trans_15_io_pipe_phv_out_data_138; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_139 = trans_15_io_pipe_phv_out_data_139; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_140 = trans_15_io_pipe_phv_out_data_140; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_141 = trans_15_io_pipe_phv_out_data_141; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_142 = trans_15_io_pipe_phv_out_data_142; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_143 = trans_15_io_pipe_phv_out_data_143; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_144 = trans_15_io_pipe_phv_out_data_144; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_145 = trans_15_io_pipe_phv_out_data_145; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_146 = trans_15_io_pipe_phv_out_data_146; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_147 = trans_15_io_pipe_phv_out_data_147; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_148 = trans_15_io_pipe_phv_out_data_148; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_149 = trans_15_io_pipe_phv_out_data_149; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_150 = trans_15_io_pipe_phv_out_data_150; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_151 = trans_15_io_pipe_phv_out_data_151; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_152 = trans_15_io_pipe_phv_out_data_152; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_153 = trans_15_io_pipe_phv_out_data_153; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_154 = trans_15_io_pipe_phv_out_data_154; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_155 = trans_15_io_pipe_phv_out_data_155; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_156 = trans_15_io_pipe_phv_out_data_156; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_157 = trans_15_io_pipe_phv_out_data_157; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_158 = trans_15_io_pipe_phv_out_data_158; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_data_159 = trans_15_io_pipe_phv_out_data_159; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_header_0 = trans_15_io_pipe_phv_out_header_0; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_header_1 = trans_15_io_pipe_phv_out_header_1; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_header_2 = trans_15_io_pipe_phv_out_header_2; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_header_3 = trans_15_io_pipe_phv_out_header_3; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_header_4 = trans_15_io_pipe_phv_out_header_4; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_header_5 = trans_15_io_pipe_phv_out_header_5; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_header_6 = trans_15_io_pipe_phv_out_header_6; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_header_7 = trans_15_io_pipe_phv_out_header_7; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_header_8 = trans_15_io_pipe_phv_out_header_8; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_header_9 = trans_15_io_pipe_phv_out_header_9; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_header_10 = trans_15_io_pipe_phv_out_header_10; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_header_11 = trans_15_io_pipe_phv_out_header_11; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_header_12 = trans_15_io_pipe_phv_out_header_12; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_header_13 = trans_15_io_pipe_phv_out_header_13; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_header_14 = trans_15_io_pipe_phv_out_header_14; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_header_15 = trans_15_io_pipe_phv_out_header_15; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_parse_current_state = trans_15_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_parse_current_offset = trans_15_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_parse_transition_field = trans_15_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_next_processor_id = trans_15_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_next_config_id = trans_15_io_pipe_phv_out_next_config_id; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_is_valid_processor = trans_15_io_pipe_phv_out_is_valid_processor; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_valid = trans_15_io_pipe_phv_out_valid; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_0_io_pipe_phv_in_last = trans_15_io_pipe_phv_out_last; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  assign proc_1_clock = clock;
  assign proc_1_io_pipe_phv_in_data_0 = init_io_pipe_phv_out_data_0; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_1 = init_io_pipe_phv_out_data_1; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_2 = init_io_pipe_phv_out_data_2; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_3 = init_io_pipe_phv_out_data_3; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_4 = init_io_pipe_phv_out_data_4; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_5 = init_io_pipe_phv_out_data_5; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_6 = init_io_pipe_phv_out_data_6; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_7 = init_io_pipe_phv_out_data_7; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_8 = init_io_pipe_phv_out_data_8; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_9 = init_io_pipe_phv_out_data_9; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_10 = init_io_pipe_phv_out_data_10; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_11 = init_io_pipe_phv_out_data_11; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_12 = init_io_pipe_phv_out_data_12; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_13 = init_io_pipe_phv_out_data_13; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_14 = init_io_pipe_phv_out_data_14; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_15 = init_io_pipe_phv_out_data_15; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_16 = init_io_pipe_phv_out_data_16; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_17 = init_io_pipe_phv_out_data_17; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_18 = init_io_pipe_phv_out_data_18; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_19 = init_io_pipe_phv_out_data_19; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_20 = init_io_pipe_phv_out_data_20; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_21 = init_io_pipe_phv_out_data_21; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_22 = init_io_pipe_phv_out_data_22; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_23 = init_io_pipe_phv_out_data_23; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_24 = init_io_pipe_phv_out_data_24; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_25 = init_io_pipe_phv_out_data_25; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_26 = init_io_pipe_phv_out_data_26; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_27 = init_io_pipe_phv_out_data_27; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_28 = init_io_pipe_phv_out_data_28; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_29 = init_io_pipe_phv_out_data_29; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_30 = init_io_pipe_phv_out_data_30; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_31 = init_io_pipe_phv_out_data_31; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_32 = init_io_pipe_phv_out_data_32; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_33 = init_io_pipe_phv_out_data_33; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_34 = init_io_pipe_phv_out_data_34; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_35 = init_io_pipe_phv_out_data_35; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_36 = init_io_pipe_phv_out_data_36; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_37 = init_io_pipe_phv_out_data_37; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_38 = init_io_pipe_phv_out_data_38; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_39 = init_io_pipe_phv_out_data_39; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_40 = init_io_pipe_phv_out_data_40; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_41 = init_io_pipe_phv_out_data_41; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_42 = init_io_pipe_phv_out_data_42; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_43 = init_io_pipe_phv_out_data_43; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_44 = init_io_pipe_phv_out_data_44; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_45 = init_io_pipe_phv_out_data_45; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_46 = init_io_pipe_phv_out_data_46; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_47 = init_io_pipe_phv_out_data_47; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_48 = init_io_pipe_phv_out_data_48; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_49 = init_io_pipe_phv_out_data_49; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_50 = init_io_pipe_phv_out_data_50; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_51 = init_io_pipe_phv_out_data_51; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_52 = init_io_pipe_phv_out_data_52; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_53 = init_io_pipe_phv_out_data_53; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_54 = init_io_pipe_phv_out_data_54; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_55 = init_io_pipe_phv_out_data_55; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_56 = init_io_pipe_phv_out_data_56; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_57 = init_io_pipe_phv_out_data_57; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_58 = init_io_pipe_phv_out_data_58; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_59 = init_io_pipe_phv_out_data_59; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_60 = init_io_pipe_phv_out_data_60; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_61 = init_io_pipe_phv_out_data_61; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_62 = init_io_pipe_phv_out_data_62; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_63 = init_io_pipe_phv_out_data_63; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_64 = init_io_pipe_phv_out_data_64; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_65 = init_io_pipe_phv_out_data_65; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_66 = init_io_pipe_phv_out_data_66; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_67 = init_io_pipe_phv_out_data_67; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_68 = init_io_pipe_phv_out_data_68; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_69 = init_io_pipe_phv_out_data_69; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_70 = init_io_pipe_phv_out_data_70; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_71 = init_io_pipe_phv_out_data_71; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_72 = init_io_pipe_phv_out_data_72; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_73 = init_io_pipe_phv_out_data_73; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_74 = init_io_pipe_phv_out_data_74; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_75 = init_io_pipe_phv_out_data_75; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_76 = init_io_pipe_phv_out_data_76; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_77 = init_io_pipe_phv_out_data_77; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_78 = init_io_pipe_phv_out_data_78; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_79 = init_io_pipe_phv_out_data_79; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_80 = init_io_pipe_phv_out_data_80; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_81 = init_io_pipe_phv_out_data_81; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_82 = init_io_pipe_phv_out_data_82; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_83 = init_io_pipe_phv_out_data_83; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_84 = init_io_pipe_phv_out_data_84; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_85 = init_io_pipe_phv_out_data_85; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_86 = init_io_pipe_phv_out_data_86; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_87 = init_io_pipe_phv_out_data_87; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_88 = init_io_pipe_phv_out_data_88; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_89 = init_io_pipe_phv_out_data_89; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_90 = init_io_pipe_phv_out_data_90; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_91 = init_io_pipe_phv_out_data_91; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_92 = init_io_pipe_phv_out_data_92; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_93 = init_io_pipe_phv_out_data_93; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_94 = init_io_pipe_phv_out_data_94; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_95 = init_io_pipe_phv_out_data_95; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_96 = init_io_pipe_phv_out_data_96; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_97 = init_io_pipe_phv_out_data_97; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_98 = init_io_pipe_phv_out_data_98; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_99 = init_io_pipe_phv_out_data_99; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_100 = init_io_pipe_phv_out_data_100; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_101 = init_io_pipe_phv_out_data_101; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_102 = init_io_pipe_phv_out_data_102; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_103 = init_io_pipe_phv_out_data_103; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_104 = init_io_pipe_phv_out_data_104; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_105 = init_io_pipe_phv_out_data_105; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_106 = init_io_pipe_phv_out_data_106; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_107 = init_io_pipe_phv_out_data_107; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_108 = init_io_pipe_phv_out_data_108; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_109 = init_io_pipe_phv_out_data_109; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_110 = init_io_pipe_phv_out_data_110; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_111 = init_io_pipe_phv_out_data_111; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_112 = init_io_pipe_phv_out_data_112; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_113 = init_io_pipe_phv_out_data_113; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_114 = init_io_pipe_phv_out_data_114; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_115 = init_io_pipe_phv_out_data_115; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_116 = init_io_pipe_phv_out_data_116; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_117 = init_io_pipe_phv_out_data_117; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_118 = init_io_pipe_phv_out_data_118; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_119 = init_io_pipe_phv_out_data_119; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_120 = init_io_pipe_phv_out_data_120; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_121 = init_io_pipe_phv_out_data_121; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_122 = init_io_pipe_phv_out_data_122; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_123 = init_io_pipe_phv_out_data_123; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_124 = init_io_pipe_phv_out_data_124; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_125 = init_io_pipe_phv_out_data_125; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_126 = init_io_pipe_phv_out_data_126; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_127 = init_io_pipe_phv_out_data_127; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_data_128 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_129 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_130 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_131 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_132 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_133 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_134 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_135 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_136 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_137 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_138 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_139 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_140 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_141 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_142 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_143 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_144 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_145 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_146 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_147 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_148 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_149 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_150 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_151 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_152 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_153 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_154 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_155 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_156 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_157 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_158 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_159 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_header_0 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_header_1 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_header_2 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_header_3 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_header_4 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_header_5 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_header_6 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_header_7 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_header_8 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_header_9 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_header_10 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_header_11 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_header_12 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_header_13 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_header_14 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_header_15 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_parse_current_state = 8'h0; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_parse_current_offset = 8'h0; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_parse_transition_field = 16'h0; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_next_processor_id = 4'h0; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_next_config_id = 1'h0; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_is_valid_processor = 1'h0; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_valid = init_io_pipe_phv_out_valid; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_1_io_pipe_phv_in_last = init_io_pipe_phv_out_last; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_clock = clock;
  assign proc_2_io_pipe_phv_in_data_0 = init_io_pipe_phv_out_data_0; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_1 = init_io_pipe_phv_out_data_1; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_2 = init_io_pipe_phv_out_data_2; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_3 = init_io_pipe_phv_out_data_3; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_4 = init_io_pipe_phv_out_data_4; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_5 = init_io_pipe_phv_out_data_5; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_6 = init_io_pipe_phv_out_data_6; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_7 = init_io_pipe_phv_out_data_7; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_8 = init_io_pipe_phv_out_data_8; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_9 = init_io_pipe_phv_out_data_9; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_10 = init_io_pipe_phv_out_data_10; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_11 = init_io_pipe_phv_out_data_11; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_12 = init_io_pipe_phv_out_data_12; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_13 = init_io_pipe_phv_out_data_13; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_14 = init_io_pipe_phv_out_data_14; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_15 = init_io_pipe_phv_out_data_15; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_16 = init_io_pipe_phv_out_data_16; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_17 = init_io_pipe_phv_out_data_17; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_18 = init_io_pipe_phv_out_data_18; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_19 = init_io_pipe_phv_out_data_19; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_20 = init_io_pipe_phv_out_data_20; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_21 = init_io_pipe_phv_out_data_21; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_22 = init_io_pipe_phv_out_data_22; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_23 = init_io_pipe_phv_out_data_23; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_24 = init_io_pipe_phv_out_data_24; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_25 = init_io_pipe_phv_out_data_25; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_26 = init_io_pipe_phv_out_data_26; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_27 = init_io_pipe_phv_out_data_27; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_28 = init_io_pipe_phv_out_data_28; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_29 = init_io_pipe_phv_out_data_29; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_30 = init_io_pipe_phv_out_data_30; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_31 = init_io_pipe_phv_out_data_31; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_32 = init_io_pipe_phv_out_data_32; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_33 = init_io_pipe_phv_out_data_33; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_34 = init_io_pipe_phv_out_data_34; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_35 = init_io_pipe_phv_out_data_35; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_36 = init_io_pipe_phv_out_data_36; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_37 = init_io_pipe_phv_out_data_37; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_38 = init_io_pipe_phv_out_data_38; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_39 = init_io_pipe_phv_out_data_39; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_40 = init_io_pipe_phv_out_data_40; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_41 = init_io_pipe_phv_out_data_41; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_42 = init_io_pipe_phv_out_data_42; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_43 = init_io_pipe_phv_out_data_43; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_44 = init_io_pipe_phv_out_data_44; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_45 = init_io_pipe_phv_out_data_45; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_46 = init_io_pipe_phv_out_data_46; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_47 = init_io_pipe_phv_out_data_47; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_48 = init_io_pipe_phv_out_data_48; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_49 = init_io_pipe_phv_out_data_49; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_50 = init_io_pipe_phv_out_data_50; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_51 = init_io_pipe_phv_out_data_51; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_52 = init_io_pipe_phv_out_data_52; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_53 = init_io_pipe_phv_out_data_53; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_54 = init_io_pipe_phv_out_data_54; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_55 = init_io_pipe_phv_out_data_55; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_56 = init_io_pipe_phv_out_data_56; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_57 = init_io_pipe_phv_out_data_57; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_58 = init_io_pipe_phv_out_data_58; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_59 = init_io_pipe_phv_out_data_59; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_60 = init_io_pipe_phv_out_data_60; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_61 = init_io_pipe_phv_out_data_61; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_62 = init_io_pipe_phv_out_data_62; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_63 = init_io_pipe_phv_out_data_63; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_64 = init_io_pipe_phv_out_data_64; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_65 = init_io_pipe_phv_out_data_65; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_66 = init_io_pipe_phv_out_data_66; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_67 = init_io_pipe_phv_out_data_67; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_68 = init_io_pipe_phv_out_data_68; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_69 = init_io_pipe_phv_out_data_69; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_70 = init_io_pipe_phv_out_data_70; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_71 = init_io_pipe_phv_out_data_71; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_72 = init_io_pipe_phv_out_data_72; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_73 = init_io_pipe_phv_out_data_73; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_74 = init_io_pipe_phv_out_data_74; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_75 = init_io_pipe_phv_out_data_75; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_76 = init_io_pipe_phv_out_data_76; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_77 = init_io_pipe_phv_out_data_77; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_78 = init_io_pipe_phv_out_data_78; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_79 = init_io_pipe_phv_out_data_79; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_80 = init_io_pipe_phv_out_data_80; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_81 = init_io_pipe_phv_out_data_81; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_82 = init_io_pipe_phv_out_data_82; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_83 = init_io_pipe_phv_out_data_83; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_84 = init_io_pipe_phv_out_data_84; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_85 = init_io_pipe_phv_out_data_85; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_86 = init_io_pipe_phv_out_data_86; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_87 = init_io_pipe_phv_out_data_87; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_88 = init_io_pipe_phv_out_data_88; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_89 = init_io_pipe_phv_out_data_89; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_90 = init_io_pipe_phv_out_data_90; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_91 = init_io_pipe_phv_out_data_91; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_92 = init_io_pipe_phv_out_data_92; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_93 = init_io_pipe_phv_out_data_93; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_94 = init_io_pipe_phv_out_data_94; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_95 = init_io_pipe_phv_out_data_95; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_96 = init_io_pipe_phv_out_data_96; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_97 = init_io_pipe_phv_out_data_97; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_98 = init_io_pipe_phv_out_data_98; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_99 = init_io_pipe_phv_out_data_99; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_100 = init_io_pipe_phv_out_data_100; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_101 = init_io_pipe_phv_out_data_101; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_102 = init_io_pipe_phv_out_data_102; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_103 = init_io_pipe_phv_out_data_103; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_104 = init_io_pipe_phv_out_data_104; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_105 = init_io_pipe_phv_out_data_105; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_106 = init_io_pipe_phv_out_data_106; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_107 = init_io_pipe_phv_out_data_107; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_108 = init_io_pipe_phv_out_data_108; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_109 = init_io_pipe_phv_out_data_109; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_110 = init_io_pipe_phv_out_data_110; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_111 = init_io_pipe_phv_out_data_111; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_112 = init_io_pipe_phv_out_data_112; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_113 = init_io_pipe_phv_out_data_113; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_114 = init_io_pipe_phv_out_data_114; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_115 = init_io_pipe_phv_out_data_115; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_116 = init_io_pipe_phv_out_data_116; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_117 = init_io_pipe_phv_out_data_117; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_118 = init_io_pipe_phv_out_data_118; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_119 = init_io_pipe_phv_out_data_119; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_120 = init_io_pipe_phv_out_data_120; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_121 = init_io_pipe_phv_out_data_121; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_122 = init_io_pipe_phv_out_data_122; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_123 = init_io_pipe_phv_out_data_123; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_124 = init_io_pipe_phv_out_data_124; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_125 = init_io_pipe_phv_out_data_125; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_126 = init_io_pipe_phv_out_data_126; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_127 = init_io_pipe_phv_out_data_127; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_data_128 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_129 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_130 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_131 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_132 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_133 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_134 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_135 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_136 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_137 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_138 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_139 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_140 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_141 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_142 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_143 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_144 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_145 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_146 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_147 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_148 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_149 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_150 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_151 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_152 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_153 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_154 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_155 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_156 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_157 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_158 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_159 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_header_0 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_header_1 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_header_2 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_header_3 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_header_4 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_header_5 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_header_6 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_header_7 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_header_8 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_header_9 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_header_10 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_header_11 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_header_12 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_header_13 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_header_14 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_header_15 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_parse_current_state = 8'h0; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_parse_current_offset = 8'h0; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_parse_transition_field = 16'h0; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_next_processor_id = 4'h0; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_next_config_id = 1'h0; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_is_valid_processor = 1'h0; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_valid = init_io_pipe_phv_out_valid; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_2_io_pipe_phv_in_last = init_io_pipe_phv_out_last; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_clock = clock;
  assign proc_3_io_pipe_phv_in_data_0 = init_io_pipe_phv_out_data_0; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_1 = init_io_pipe_phv_out_data_1; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_2 = init_io_pipe_phv_out_data_2; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_3 = init_io_pipe_phv_out_data_3; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_4 = init_io_pipe_phv_out_data_4; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_5 = init_io_pipe_phv_out_data_5; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_6 = init_io_pipe_phv_out_data_6; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_7 = init_io_pipe_phv_out_data_7; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_8 = init_io_pipe_phv_out_data_8; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_9 = init_io_pipe_phv_out_data_9; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_10 = init_io_pipe_phv_out_data_10; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_11 = init_io_pipe_phv_out_data_11; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_12 = init_io_pipe_phv_out_data_12; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_13 = init_io_pipe_phv_out_data_13; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_14 = init_io_pipe_phv_out_data_14; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_15 = init_io_pipe_phv_out_data_15; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_16 = init_io_pipe_phv_out_data_16; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_17 = init_io_pipe_phv_out_data_17; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_18 = init_io_pipe_phv_out_data_18; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_19 = init_io_pipe_phv_out_data_19; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_20 = init_io_pipe_phv_out_data_20; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_21 = init_io_pipe_phv_out_data_21; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_22 = init_io_pipe_phv_out_data_22; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_23 = init_io_pipe_phv_out_data_23; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_24 = init_io_pipe_phv_out_data_24; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_25 = init_io_pipe_phv_out_data_25; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_26 = init_io_pipe_phv_out_data_26; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_27 = init_io_pipe_phv_out_data_27; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_28 = init_io_pipe_phv_out_data_28; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_29 = init_io_pipe_phv_out_data_29; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_30 = init_io_pipe_phv_out_data_30; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_31 = init_io_pipe_phv_out_data_31; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_32 = init_io_pipe_phv_out_data_32; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_33 = init_io_pipe_phv_out_data_33; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_34 = init_io_pipe_phv_out_data_34; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_35 = init_io_pipe_phv_out_data_35; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_36 = init_io_pipe_phv_out_data_36; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_37 = init_io_pipe_phv_out_data_37; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_38 = init_io_pipe_phv_out_data_38; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_39 = init_io_pipe_phv_out_data_39; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_40 = init_io_pipe_phv_out_data_40; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_41 = init_io_pipe_phv_out_data_41; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_42 = init_io_pipe_phv_out_data_42; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_43 = init_io_pipe_phv_out_data_43; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_44 = init_io_pipe_phv_out_data_44; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_45 = init_io_pipe_phv_out_data_45; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_46 = init_io_pipe_phv_out_data_46; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_47 = init_io_pipe_phv_out_data_47; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_48 = init_io_pipe_phv_out_data_48; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_49 = init_io_pipe_phv_out_data_49; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_50 = init_io_pipe_phv_out_data_50; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_51 = init_io_pipe_phv_out_data_51; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_52 = init_io_pipe_phv_out_data_52; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_53 = init_io_pipe_phv_out_data_53; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_54 = init_io_pipe_phv_out_data_54; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_55 = init_io_pipe_phv_out_data_55; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_56 = init_io_pipe_phv_out_data_56; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_57 = init_io_pipe_phv_out_data_57; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_58 = init_io_pipe_phv_out_data_58; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_59 = init_io_pipe_phv_out_data_59; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_60 = init_io_pipe_phv_out_data_60; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_61 = init_io_pipe_phv_out_data_61; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_62 = init_io_pipe_phv_out_data_62; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_63 = init_io_pipe_phv_out_data_63; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_64 = init_io_pipe_phv_out_data_64; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_65 = init_io_pipe_phv_out_data_65; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_66 = init_io_pipe_phv_out_data_66; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_67 = init_io_pipe_phv_out_data_67; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_68 = init_io_pipe_phv_out_data_68; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_69 = init_io_pipe_phv_out_data_69; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_70 = init_io_pipe_phv_out_data_70; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_71 = init_io_pipe_phv_out_data_71; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_72 = init_io_pipe_phv_out_data_72; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_73 = init_io_pipe_phv_out_data_73; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_74 = init_io_pipe_phv_out_data_74; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_75 = init_io_pipe_phv_out_data_75; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_76 = init_io_pipe_phv_out_data_76; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_77 = init_io_pipe_phv_out_data_77; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_78 = init_io_pipe_phv_out_data_78; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_79 = init_io_pipe_phv_out_data_79; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_80 = init_io_pipe_phv_out_data_80; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_81 = init_io_pipe_phv_out_data_81; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_82 = init_io_pipe_phv_out_data_82; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_83 = init_io_pipe_phv_out_data_83; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_84 = init_io_pipe_phv_out_data_84; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_85 = init_io_pipe_phv_out_data_85; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_86 = init_io_pipe_phv_out_data_86; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_87 = init_io_pipe_phv_out_data_87; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_88 = init_io_pipe_phv_out_data_88; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_89 = init_io_pipe_phv_out_data_89; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_90 = init_io_pipe_phv_out_data_90; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_91 = init_io_pipe_phv_out_data_91; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_92 = init_io_pipe_phv_out_data_92; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_93 = init_io_pipe_phv_out_data_93; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_94 = init_io_pipe_phv_out_data_94; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_95 = init_io_pipe_phv_out_data_95; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_96 = init_io_pipe_phv_out_data_96; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_97 = init_io_pipe_phv_out_data_97; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_98 = init_io_pipe_phv_out_data_98; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_99 = init_io_pipe_phv_out_data_99; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_100 = init_io_pipe_phv_out_data_100; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_101 = init_io_pipe_phv_out_data_101; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_102 = init_io_pipe_phv_out_data_102; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_103 = init_io_pipe_phv_out_data_103; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_104 = init_io_pipe_phv_out_data_104; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_105 = init_io_pipe_phv_out_data_105; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_106 = init_io_pipe_phv_out_data_106; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_107 = init_io_pipe_phv_out_data_107; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_108 = init_io_pipe_phv_out_data_108; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_109 = init_io_pipe_phv_out_data_109; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_110 = init_io_pipe_phv_out_data_110; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_111 = init_io_pipe_phv_out_data_111; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_112 = init_io_pipe_phv_out_data_112; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_113 = init_io_pipe_phv_out_data_113; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_114 = init_io_pipe_phv_out_data_114; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_115 = init_io_pipe_phv_out_data_115; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_116 = init_io_pipe_phv_out_data_116; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_117 = init_io_pipe_phv_out_data_117; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_118 = init_io_pipe_phv_out_data_118; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_119 = init_io_pipe_phv_out_data_119; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_120 = init_io_pipe_phv_out_data_120; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_121 = init_io_pipe_phv_out_data_121; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_122 = init_io_pipe_phv_out_data_122; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_123 = init_io_pipe_phv_out_data_123; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_124 = init_io_pipe_phv_out_data_124; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_125 = init_io_pipe_phv_out_data_125; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_126 = init_io_pipe_phv_out_data_126; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_127 = init_io_pipe_phv_out_data_127; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_data_128 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_129 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_130 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_131 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_132 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_133 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_134 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_135 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_136 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_137 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_138 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_139 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_140 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_141 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_142 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_143 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_144 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_145 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_146 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_147 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_148 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_149 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_150 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_151 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_152 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_153 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_154 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_155 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_156 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_157 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_158 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_159 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_header_0 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_header_1 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_header_2 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_header_3 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_header_4 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_header_5 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_header_6 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_header_7 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_header_8 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_header_9 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_header_10 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_header_11 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_header_12 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_header_13 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_header_14 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_header_15 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_parse_current_state = 8'h0; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_parse_current_offset = 8'h0; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_parse_transition_field = 16'h0; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_next_processor_id = 4'h0; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_next_config_id = 1'h0; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_is_valid_processor = 1'h0; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_valid = init_io_pipe_phv_out_valid; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_3_io_pipe_phv_in_last = init_io_pipe_phv_out_last; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_clock = clock;
  assign proc_4_io_pipe_phv_in_data_0 = init_io_pipe_phv_out_data_0; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_1 = init_io_pipe_phv_out_data_1; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_2 = init_io_pipe_phv_out_data_2; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_3 = init_io_pipe_phv_out_data_3; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_4 = init_io_pipe_phv_out_data_4; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_5 = init_io_pipe_phv_out_data_5; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_6 = init_io_pipe_phv_out_data_6; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_7 = init_io_pipe_phv_out_data_7; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_8 = init_io_pipe_phv_out_data_8; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_9 = init_io_pipe_phv_out_data_9; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_10 = init_io_pipe_phv_out_data_10; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_11 = init_io_pipe_phv_out_data_11; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_12 = init_io_pipe_phv_out_data_12; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_13 = init_io_pipe_phv_out_data_13; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_14 = init_io_pipe_phv_out_data_14; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_15 = init_io_pipe_phv_out_data_15; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_16 = init_io_pipe_phv_out_data_16; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_17 = init_io_pipe_phv_out_data_17; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_18 = init_io_pipe_phv_out_data_18; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_19 = init_io_pipe_phv_out_data_19; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_20 = init_io_pipe_phv_out_data_20; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_21 = init_io_pipe_phv_out_data_21; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_22 = init_io_pipe_phv_out_data_22; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_23 = init_io_pipe_phv_out_data_23; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_24 = init_io_pipe_phv_out_data_24; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_25 = init_io_pipe_phv_out_data_25; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_26 = init_io_pipe_phv_out_data_26; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_27 = init_io_pipe_phv_out_data_27; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_28 = init_io_pipe_phv_out_data_28; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_29 = init_io_pipe_phv_out_data_29; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_30 = init_io_pipe_phv_out_data_30; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_31 = init_io_pipe_phv_out_data_31; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_32 = init_io_pipe_phv_out_data_32; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_33 = init_io_pipe_phv_out_data_33; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_34 = init_io_pipe_phv_out_data_34; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_35 = init_io_pipe_phv_out_data_35; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_36 = init_io_pipe_phv_out_data_36; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_37 = init_io_pipe_phv_out_data_37; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_38 = init_io_pipe_phv_out_data_38; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_39 = init_io_pipe_phv_out_data_39; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_40 = init_io_pipe_phv_out_data_40; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_41 = init_io_pipe_phv_out_data_41; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_42 = init_io_pipe_phv_out_data_42; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_43 = init_io_pipe_phv_out_data_43; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_44 = init_io_pipe_phv_out_data_44; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_45 = init_io_pipe_phv_out_data_45; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_46 = init_io_pipe_phv_out_data_46; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_47 = init_io_pipe_phv_out_data_47; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_48 = init_io_pipe_phv_out_data_48; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_49 = init_io_pipe_phv_out_data_49; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_50 = init_io_pipe_phv_out_data_50; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_51 = init_io_pipe_phv_out_data_51; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_52 = init_io_pipe_phv_out_data_52; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_53 = init_io_pipe_phv_out_data_53; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_54 = init_io_pipe_phv_out_data_54; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_55 = init_io_pipe_phv_out_data_55; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_56 = init_io_pipe_phv_out_data_56; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_57 = init_io_pipe_phv_out_data_57; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_58 = init_io_pipe_phv_out_data_58; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_59 = init_io_pipe_phv_out_data_59; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_60 = init_io_pipe_phv_out_data_60; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_61 = init_io_pipe_phv_out_data_61; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_62 = init_io_pipe_phv_out_data_62; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_63 = init_io_pipe_phv_out_data_63; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_64 = init_io_pipe_phv_out_data_64; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_65 = init_io_pipe_phv_out_data_65; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_66 = init_io_pipe_phv_out_data_66; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_67 = init_io_pipe_phv_out_data_67; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_68 = init_io_pipe_phv_out_data_68; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_69 = init_io_pipe_phv_out_data_69; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_70 = init_io_pipe_phv_out_data_70; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_71 = init_io_pipe_phv_out_data_71; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_72 = init_io_pipe_phv_out_data_72; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_73 = init_io_pipe_phv_out_data_73; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_74 = init_io_pipe_phv_out_data_74; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_75 = init_io_pipe_phv_out_data_75; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_76 = init_io_pipe_phv_out_data_76; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_77 = init_io_pipe_phv_out_data_77; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_78 = init_io_pipe_phv_out_data_78; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_79 = init_io_pipe_phv_out_data_79; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_80 = init_io_pipe_phv_out_data_80; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_81 = init_io_pipe_phv_out_data_81; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_82 = init_io_pipe_phv_out_data_82; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_83 = init_io_pipe_phv_out_data_83; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_84 = init_io_pipe_phv_out_data_84; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_85 = init_io_pipe_phv_out_data_85; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_86 = init_io_pipe_phv_out_data_86; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_87 = init_io_pipe_phv_out_data_87; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_88 = init_io_pipe_phv_out_data_88; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_89 = init_io_pipe_phv_out_data_89; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_90 = init_io_pipe_phv_out_data_90; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_91 = init_io_pipe_phv_out_data_91; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_92 = init_io_pipe_phv_out_data_92; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_93 = init_io_pipe_phv_out_data_93; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_94 = init_io_pipe_phv_out_data_94; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_95 = init_io_pipe_phv_out_data_95; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_96 = init_io_pipe_phv_out_data_96; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_97 = init_io_pipe_phv_out_data_97; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_98 = init_io_pipe_phv_out_data_98; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_99 = init_io_pipe_phv_out_data_99; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_100 = init_io_pipe_phv_out_data_100; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_101 = init_io_pipe_phv_out_data_101; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_102 = init_io_pipe_phv_out_data_102; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_103 = init_io_pipe_phv_out_data_103; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_104 = init_io_pipe_phv_out_data_104; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_105 = init_io_pipe_phv_out_data_105; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_106 = init_io_pipe_phv_out_data_106; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_107 = init_io_pipe_phv_out_data_107; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_108 = init_io_pipe_phv_out_data_108; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_109 = init_io_pipe_phv_out_data_109; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_110 = init_io_pipe_phv_out_data_110; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_111 = init_io_pipe_phv_out_data_111; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_112 = init_io_pipe_phv_out_data_112; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_113 = init_io_pipe_phv_out_data_113; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_114 = init_io_pipe_phv_out_data_114; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_115 = init_io_pipe_phv_out_data_115; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_116 = init_io_pipe_phv_out_data_116; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_117 = init_io_pipe_phv_out_data_117; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_118 = init_io_pipe_phv_out_data_118; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_119 = init_io_pipe_phv_out_data_119; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_120 = init_io_pipe_phv_out_data_120; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_121 = init_io_pipe_phv_out_data_121; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_122 = init_io_pipe_phv_out_data_122; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_123 = init_io_pipe_phv_out_data_123; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_124 = init_io_pipe_phv_out_data_124; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_125 = init_io_pipe_phv_out_data_125; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_126 = init_io_pipe_phv_out_data_126; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_127 = init_io_pipe_phv_out_data_127; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_data_128 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_4_io_pipe_phv_in_data_129 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_4_io_pipe_phv_in_data_130 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_4_io_pipe_phv_in_data_131 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_4_io_pipe_phv_in_data_132 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_4_io_pipe_phv_in_data_133 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_4_io_pipe_phv_in_data_134 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_4_io_pipe_phv_in_data_135 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_4_io_pipe_phv_in_data_136 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_4_io_pipe_phv_in_data_137 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_4_io_pipe_phv_in_data_138 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_4_io_pipe_phv_in_data_139 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_4_io_pipe_phv_in_data_140 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_4_io_pipe_phv_in_data_141 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_4_io_pipe_phv_in_data_142 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_4_io_pipe_phv_in_data_143 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_4_io_pipe_phv_in_data_144 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_4_io_pipe_phv_in_data_145 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_4_io_pipe_phv_in_data_146 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_4_io_pipe_phv_in_data_147 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_4_io_pipe_phv_in_data_148 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_4_io_pipe_phv_in_data_149 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_4_io_pipe_phv_in_data_150 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_4_io_pipe_phv_in_data_151 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_4_io_pipe_phv_in_data_152 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_4_io_pipe_phv_in_data_153 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_4_io_pipe_phv_in_data_154 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_4_io_pipe_phv_in_data_155 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_4_io_pipe_phv_in_data_156 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_4_io_pipe_phv_in_data_157 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_4_io_pipe_phv_in_data_158 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_4_io_pipe_phv_in_data_159 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_4_io_pipe_phv_in_header_0 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_4_io_pipe_phv_in_header_1 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_4_io_pipe_phv_in_header_2 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_4_io_pipe_phv_in_header_3 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_4_io_pipe_phv_in_header_4 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_4_io_pipe_phv_in_header_5 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_4_io_pipe_phv_in_header_6 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_4_io_pipe_phv_in_header_7 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_4_io_pipe_phv_in_header_8 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_4_io_pipe_phv_in_header_9 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_4_io_pipe_phv_in_header_10 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_4_io_pipe_phv_in_header_11 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_4_io_pipe_phv_in_header_12 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_4_io_pipe_phv_in_header_13 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_4_io_pipe_phv_in_header_14 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_4_io_pipe_phv_in_header_15 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_4_io_pipe_phv_in_parse_current_state = 8'h0; // @[ipsa.scala 94:65]
  assign proc_4_io_pipe_phv_in_parse_current_offset = 8'h0; // @[ipsa.scala 94:65]
  assign proc_4_io_pipe_phv_in_parse_transition_field = 16'h0; // @[ipsa.scala 94:65]
  assign proc_4_io_pipe_phv_in_next_processor_id = 4'h0; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_next_config_id = 1'h0; // @[ipsa.scala 94:65]
  assign proc_4_io_pipe_phv_in_is_valid_processor = 1'h0; // @[ipsa.scala 94:65]
  assign proc_4_io_pipe_phv_in_valid = init_io_pipe_phv_out_valid; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_4_io_pipe_phv_in_last = init_io_pipe_phv_out_last; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_clock = clock;
  assign proc_5_io_pipe_phv_in_data_0 = init_io_pipe_phv_out_data_0; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_1 = init_io_pipe_phv_out_data_1; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_2 = init_io_pipe_phv_out_data_2; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_3 = init_io_pipe_phv_out_data_3; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_4 = init_io_pipe_phv_out_data_4; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_5 = init_io_pipe_phv_out_data_5; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_6 = init_io_pipe_phv_out_data_6; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_7 = init_io_pipe_phv_out_data_7; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_8 = init_io_pipe_phv_out_data_8; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_9 = init_io_pipe_phv_out_data_9; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_10 = init_io_pipe_phv_out_data_10; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_11 = init_io_pipe_phv_out_data_11; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_12 = init_io_pipe_phv_out_data_12; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_13 = init_io_pipe_phv_out_data_13; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_14 = init_io_pipe_phv_out_data_14; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_15 = init_io_pipe_phv_out_data_15; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_16 = init_io_pipe_phv_out_data_16; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_17 = init_io_pipe_phv_out_data_17; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_18 = init_io_pipe_phv_out_data_18; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_19 = init_io_pipe_phv_out_data_19; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_20 = init_io_pipe_phv_out_data_20; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_21 = init_io_pipe_phv_out_data_21; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_22 = init_io_pipe_phv_out_data_22; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_23 = init_io_pipe_phv_out_data_23; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_24 = init_io_pipe_phv_out_data_24; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_25 = init_io_pipe_phv_out_data_25; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_26 = init_io_pipe_phv_out_data_26; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_27 = init_io_pipe_phv_out_data_27; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_28 = init_io_pipe_phv_out_data_28; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_29 = init_io_pipe_phv_out_data_29; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_30 = init_io_pipe_phv_out_data_30; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_31 = init_io_pipe_phv_out_data_31; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_32 = init_io_pipe_phv_out_data_32; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_33 = init_io_pipe_phv_out_data_33; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_34 = init_io_pipe_phv_out_data_34; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_35 = init_io_pipe_phv_out_data_35; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_36 = init_io_pipe_phv_out_data_36; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_37 = init_io_pipe_phv_out_data_37; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_38 = init_io_pipe_phv_out_data_38; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_39 = init_io_pipe_phv_out_data_39; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_40 = init_io_pipe_phv_out_data_40; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_41 = init_io_pipe_phv_out_data_41; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_42 = init_io_pipe_phv_out_data_42; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_43 = init_io_pipe_phv_out_data_43; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_44 = init_io_pipe_phv_out_data_44; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_45 = init_io_pipe_phv_out_data_45; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_46 = init_io_pipe_phv_out_data_46; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_47 = init_io_pipe_phv_out_data_47; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_48 = init_io_pipe_phv_out_data_48; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_49 = init_io_pipe_phv_out_data_49; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_50 = init_io_pipe_phv_out_data_50; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_51 = init_io_pipe_phv_out_data_51; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_52 = init_io_pipe_phv_out_data_52; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_53 = init_io_pipe_phv_out_data_53; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_54 = init_io_pipe_phv_out_data_54; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_55 = init_io_pipe_phv_out_data_55; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_56 = init_io_pipe_phv_out_data_56; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_57 = init_io_pipe_phv_out_data_57; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_58 = init_io_pipe_phv_out_data_58; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_59 = init_io_pipe_phv_out_data_59; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_60 = init_io_pipe_phv_out_data_60; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_61 = init_io_pipe_phv_out_data_61; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_62 = init_io_pipe_phv_out_data_62; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_63 = init_io_pipe_phv_out_data_63; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_64 = init_io_pipe_phv_out_data_64; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_65 = init_io_pipe_phv_out_data_65; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_66 = init_io_pipe_phv_out_data_66; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_67 = init_io_pipe_phv_out_data_67; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_68 = init_io_pipe_phv_out_data_68; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_69 = init_io_pipe_phv_out_data_69; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_70 = init_io_pipe_phv_out_data_70; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_71 = init_io_pipe_phv_out_data_71; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_72 = init_io_pipe_phv_out_data_72; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_73 = init_io_pipe_phv_out_data_73; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_74 = init_io_pipe_phv_out_data_74; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_75 = init_io_pipe_phv_out_data_75; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_76 = init_io_pipe_phv_out_data_76; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_77 = init_io_pipe_phv_out_data_77; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_78 = init_io_pipe_phv_out_data_78; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_79 = init_io_pipe_phv_out_data_79; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_80 = init_io_pipe_phv_out_data_80; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_81 = init_io_pipe_phv_out_data_81; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_82 = init_io_pipe_phv_out_data_82; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_83 = init_io_pipe_phv_out_data_83; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_84 = init_io_pipe_phv_out_data_84; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_85 = init_io_pipe_phv_out_data_85; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_86 = init_io_pipe_phv_out_data_86; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_87 = init_io_pipe_phv_out_data_87; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_88 = init_io_pipe_phv_out_data_88; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_89 = init_io_pipe_phv_out_data_89; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_90 = init_io_pipe_phv_out_data_90; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_91 = init_io_pipe_phv_out_data_91; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_92 = init_io_pipe_phv_out_data_92; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_93 = init_io_pipe_phv_out_data_93; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_94 = init_io_pipe_phv_out_data_94; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_95 = init_io_pipe_phv_out_data_95; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_96 = init_io_pipe_phv_out_data_96; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_97 = init_io_pipe_phv_out_data_97; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_98 = init_io_pipe_phv_out_data_98; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_99 = init_io_pipe_phv_out_data_99; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_100 = init_io_pipe_phv_out_data_100; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_101 = init_io_pipe_phv_out_data_101; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_102 = init_io_pipe_phv_out_data_102; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_103 = init_io_pipe_phv_out_data_103; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_104 = init_io_pipe_phv_out_data_104; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_105 = init_io_pipe_phv_out_data_105; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_106 = init_io_pipe_phv_out_data_106; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_107 = init_io_pipe_phv_out_data_107; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_108 = init_io_pipe_phv_out_data_108; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_109 = init_io_pipe_phv_out_data_109; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_110 = init_io_pipe_phv_out_data_110; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_111 = init_io_pipe_phv_out_data_111; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_112 = init_io_pipe_phv_out_data_112; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_113 = init_io_pipe_phv_out_data_113; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_114 = init_io_pipe_phv_out_data_114; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_115 = init_io_pipe_phv_out_data_115; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_116 = init_io_pipe_phv_out_data_116; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_117 = init_io_pipe_phv_out_data_117; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_118 = init_io_pipe_phv_out_data_118; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_119 = init_io_pipe_phv_out_data_119; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_120 = init_io_pipe_phv_out_data_120; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_121 = init_io_pipe_phv_out_data_121; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_122 = init_io_pipe_phv_out_data_122; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_123 = init_io_pipe_phv_out_data_123; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_124 = init_io_pipe_phv_out_data_124; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_125 = init_io_pipe_phv_out_data_125; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_126 = init_io_pipe_phv_out_data_126; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_127 = init_io_pipe_phv_out_data_127; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_data_128 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_5_io_pipe_phv_in_data_129 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_5_io_pipe_phv_in_data_130 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_5_io_pipe_phv_in_data_131 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_5_io_pipe_phv_in_data_132 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_5_io_pipe_phv_in_data_133 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_5_io_pipe_phv_in_data_134 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_5_io_pipe_phv_in_data_135 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_5_io_pipe_phv_in_data_136 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_5_io_pipe_phv_in_data_137 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_5_io_pipe_phv_in_data_138 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_5_io_pipe_phv_in_data_139 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_5_io_pipe_phv_in_data_140 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_5_io_pipe_phv_in_data_141 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_5_io_pipe_phv_in_data_142 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_5_io_pipe_phv_in_data_143 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_5_io_pipe_phv_in_data_144 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_5_io_pipe_phv_in_data_145 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_5_io_pipe_phv_in_data_146 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_5_io_pipe_phv_in_data_147 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_5_io_pipe_phv_in_data_148 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_5_io_pipe_phv_in_data_149 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_5_io_pipe_phv_in_data_150 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_5_io_pipe_phv_in_data_151 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_5_io_pipe_phv_in_data_152 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_5_io_pipe_phv_in_data_153 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_5_io_pipe_phv_in_data_154 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_5_io_pipe_phv_in_data_155 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_5_io_pipe_phv_in_data_156 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_5_io_pipe_phv_in_data_157 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_5_io_pipe_phv_in_data_158 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_5_io_pipe_phv_in_data_159 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_5_io_pipe_phv_in_header_0 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_5_io_pipe_phv_in_header_1 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_5_io_pipe_phv_in_header_2 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_5_io_pipe_phv_in_header_3 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_5_io_pipe_phv_in_header_4 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_5_io_pipe_phv_in_header_5 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_5_io_pipe_phv_in_header_6 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_5_io_pipe_phv_in_header_7 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_5_io_pipe_phv_in_header_8 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_5_io_pipe_phv_in_header_9 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_5_io_pipe_phv_in_header_10 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_5_io_pipe_phv_in_header_11 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_5_io_pipe_phv_in_header_12 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_5_io_pipe_phv_in_header_13 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_5_io_pipe_phv_in_header_14 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_5_io_pipe_phv_in_header_15 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_5_io_pipe_phv_in_parse_current_state = 8'h0; // @[ipsa.scala 94:65]
  assign proc_5_io_pipe_phv_in_parse_current_offset = 8'h0; // @[ipsa.scala 94:65]
  assign proc_5_io_pipe_phv_in_parse_transition_field = 16'h0; // @[ipsa.scala 94:65]
  assign proc_5_io_pipe_phv_in_next_processor_id = 4'h0; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_next_config_id = 1'h0; // @[ipsa.scala 94:65]
  assign proc_5_io_pipe_phv_in_is_valid_processor = 1'h0; // @[ipsa.scala 94:65]
  assign proc_5_io_pipe_phv_in_valid = init_io_pipe_phv_out_valid; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_5_io_pipe_phv_in_last = init_io_pipe_phv_out_last; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_clock = clock;
  assign proc_6_io_pipe_phv_in_data_0 = init_io_pipe_phv_out_data_0; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_1 = init_io_pipe_phv_out_data_1; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_2 = init_io_pipe_phv_out_data_2; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_3 = init_io_pipe_phv_out_data_3; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_4 = init_io_pipe_phv_out_data_4; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_5 = init_io_pipe_phv_out_data_5; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_6 = init_io_pipe_phv_out_data_6; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_7 = init_io_pipe_phv_out_data_7; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_8 = init_io_pipe_phv_out_data_8; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_9 = init_io_pipe_phv_out_data_9; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_10 = init_io_pipe_phv_out_data_10; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_11 = init_io_pipe_phv_out_data_11; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_12 = init_io_pipe_phv_out_data_12; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_13 = init_io_pipe_phv_out_data_13; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_14 = init_io_pipe_phv_out_data_14; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_15 = init_io_pipe_phv_out_data_15; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_16 = init_io_pipe_phv_out_data_16; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_17 = init_io_pipe_phv_out_data_17; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_18 = init_io_pipe_phv_out_data_18; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_19 = init_io_pipe_phv_out_data_19; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_20 = init_io_pipe_phv_out_data_20; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_21 = init_io_pipe_phv_out_data_21; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_22 = init_io_pipe_phv_out_data_22; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_23 = init_io_pipe_phv_out_data_23; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_24 = init_io_pipe_phv_out_data_24; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_25 = init_io_pipe_phv_out_data_25; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_26 = init_io_pipe_phv_out_data_26; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_27 = init_io_pipe_phv_out_data_27; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_28 = init_io_pipe_phv_out_data_28; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_29 = init_io_pipe_phv_out_data_29; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_30 = init_io_pipe_phv_out_data_30; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_31 = init_io_pipe_phv_out_data_31; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_32 = init_io_pipe_phv_out_data_32; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_33 = init_io_pipe_phv_out_data_33; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_34 = init_io_pipe_phv_out_data_34; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_35 = init_io_pipe_phv_out_data_35; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_36 = init_io_pipe_phv_out_data_36; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_37 = init_io_pipe_phv_out_data_37; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_38 = init_io_pipe_phv_out_data_38; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_39 = init_io_pipe_phv_out_data_39; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_40 = init_io_pipe_phv_out_data_40; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_41 = init_io_pipe_phv_out_data_41; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_42 = init_io_pipe_phv_out_data_42; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_43 = init_io_pipe_phv_out_data_43; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_44 = init_io_pipe_phv_out_data_44; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_45 = init_io_pipe_phv_out_data_45; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_46 = init_io_pipe_phv_out_data_46; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_47 = init_io_pipe_phv_out_data_47; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_48 = init_io_pipe_phv_out_data_48; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_49 = init_io_pipe_phv_out_data_49; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_50 = init_io_pipe_phv_out_data_50; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_51 = init_io_pipe_phv_out_data_51; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_52 = init_io_pipe_phv_out_data_52; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_53 = init_io_pipe_phv_out_data_53; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_54 = init_io_pipe_phv_out_data_54; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_55 = init_io_pipe_phv_out_data_55; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_56 = init_io_pipe_phv_out_data_56; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_57 = init_io_pipe_phv_out_data_57; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_58 = init_io_pipe_phv_out_data_58; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_59 = init_io_pipe_phv_out_data_59; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_60 = init_io_pipe_phv_out_data_60; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_61 = init_io_pipe_phv_out_data_61; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_62 = init_io_pipe_phv_out_data_62; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_63 = init_io_pipe_phv_out_data_63; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_64 = init_io_pipe_phv_out_data_64; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_65 = init_io_pipe_phv_out_data_65; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_66 = init_io_pipe_phv_out_data_66; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_67 = init_io_pipe_phv_out_data_67; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_68 = init_io_pipe_phv_out_data_68; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_69 = init_io_pipe_phv_out_data_69; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_70 = init_io_pipe_phv_out_data_70; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_71 = init_io_pipe_phv_out_data_71; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_72 = init_io_pipe_phv_out_data_72; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_73 = init_io_pipe_phv_out_data_73; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_74 = init_io_pipe_phv_out_data_74; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_75 = init_io_pipe_phv_out_data_75; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_76 = init_io_pipe_phv_out_data_76; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_77 = init_io_pipe_phv_out_data_77; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_78 = init_io_pipe_phv_out_data_78; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_79 = init_io_pipe_phv_out_data_79; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_80 = init_io_pipe_phv_out_data_80; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_81 = init_io_pipe_phv_out_data_81; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_82 = init_io_pipe_phv_out_data_82; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_83 = init_io_pipe_phv_out_data_83; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_84 = init_io_pipe_phv_out_data_84; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_85 = init_io_pipe_phv_out_data_85; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_86 = init_io_pipe_phv_out_data_86; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_87 = init_io_pipe_phv_out_data_87; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_88 = init_io_pipe_phv_out_data_88; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_89 = init_io_pipe_phv_out_data_89; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_90 = init_io_pipe_phv_out_data_90; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_91 = init_io_pipe_phv_out_data_91; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_92 = init_io_pipe_phv_out_data_92; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_93 = init_io_pipe_phv_out_data_93; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_94 = init_io_pipe_phv_out_data_94; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_95 = init_io_pipe_phv_out_data_95; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_96 = init_io_pipe_phv_out_data_96; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_97 = init_io_pipe_phv_out_data_97; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_98 = init_io_pipe_phv_out_data_98; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_99 = init_io_pipe_phv_out_data_99; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_100 = init_io_pipe_phv_out_data_100; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_101 = init_io_pipe_phv_out_data_101; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_102 = init_io_pipe_phv_out_data_102; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_103 = init_io_pipe_phv_out_data_103; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_104 = init_io_pipe_phv_out_data_104; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_105 = init_io_pipe_phv_out_data_105; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_106 = init_io_pipe_phv_out_data_106; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_107 = init_io_pipe_phv_out_data_107; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_108 = init_io_pipe_phv_out_data_108; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_109 = init_io_pipe_phv_out_data_109; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_110 = init_io_pipe_phv_out_data_110; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_111 = init_io_pipe_phv_out_data_111; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_112 = init_io_pipe_phv_out_data_112; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_113 = init_io_pipe_phv_out_data_113; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_114 = init_io_pipe_phv_out_data_114; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_115 = init_io_pipe_phv_out_data_115; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_116 = init_io_pipe_phv_out_data_116; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_117 = init_io_pipe_phv_out_data_117; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_118 = init_io_pipe_phv_out_data_118; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_119 = init_io_pipe_phv_out_data_119; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_120 = init_io_pipe_phv_out_data_120; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_121 = init_io_pipe_phv_out_data_121; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_122 = init_io_pipe_phv_out_data_122; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_123 = init_io_pipe_phv_out_data_123; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_124 = init_io_pipe_phv_out_data_124; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_125 = init_io_pipe_phv_out_data_125; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_126 = init_io_pipe_phv_out_data_126; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_127 = init_io_pipe_phv_out_data_127; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_data_128 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_6_io_pipe_phv_in_data_129 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_6_io_pipe_phv_in_data_130 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_6_io_pipe_phv_in_data_131 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_6_io_pipe_phv_in_data_132 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_6_io_pipe_phv_in_data_133 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_6_io_pipe_phv_in_data_134 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_6_io_pipe_phv_in_data_135 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_6_io_pipe_phv_in_data_136 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_6_io_pipe_phv_in_data_137 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_6_io_pipe_phv_in_data_138 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_6_io_pipe_phv_in_data_139 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_6_io_pipe_phv_in_data_140 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_6_io_pipe_phv_in_data_141 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_6_io_pipe_phv_in_data_142 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_6_io_pipe_phv_in_data_143 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_6_io_pipe_phv_in_data_144 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_6_io_pipe_phv_in_data_145 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_6_io_pipe_phv_in_data_146 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_6_io_pipe_phv_in_data_147 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_6_io_pipe_phv_in_data_148 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_6_io_pipe_phv_in_data_149 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_6_io_pipe_phv_in_data_150 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_6_io_pipe_phv_in_data_151 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_6_io_pipe_phv_in_data_152 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_6_io_pipe_phv_in_data_153 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_6_io_pipe_phv_in_data_154 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_6_io_pipe_phv_in_data_155 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_6_io_pipe_phv_in_data_156 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_6_io_pipe_phv_in_data_157 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_6_io_pipe_phv_in_data_158 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_6_io_pipe_phv_in_data_159 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_6_io_pipe_phv_in_header_0 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_6_io_pipe_phv_in_header_1 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_6_io_pipe_phv_in_header_2 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_6_io_pipe_phv_in_header_3 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_6_io_pipe_phv_in_header_4 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_6_io_pipe_phv_in_header_5 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_6_io_pipe_phv_in_header_6 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_6_io_pipe_phv_in_header_7 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_6_io_pipe_phv_in_header_8 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_6_io_pipe_phv_in_header_9 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_6_io_pipe_phv_in_header_10 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_6_io_pipe_phv_in_header_11 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_6_io_pipe_phv_in_header_12 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_6_io_pipe_phv_in_header_13 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_6_io_pipe_phv_in_header_14 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_6_io_pipe_phv_in_header_15 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_6_io_pipe_phv_in_parse_current_state = 8'h0; // @[ipsa.scala 94:65]
  assign proc_6_io_pipe_phv_in_parse_current_offset = 8'h0; // @[ipsa.scala 94:65]
  assign proc_6_io_pipe_phv_in_parse_transition_field = 16'h0; // @[ipsa.scala 94:65]
  assign proc_6_io_pipe_phv_in_next_processor_id = 4'h0; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_next_config_id = 1'h0; // @[ipsa.scala 94:65]
  assign proc_6_io_pipe_phv_in_is_valid_processor = 1'h0; // @[ipsa.scala 94:65]
  assign proc_6_io_pipe_phv_in_valid = init_io_pipe_phv_out_valid; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_6_io_pipe_phv_in_last = init_io_pipe_phv_out_last; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_clock = clock;
  assign proc_7_io_pipe_phv_in_data_0 = init_io_pipe_phv_out_data_0; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_1 = init_io_pipe_phv_out_data_1; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_2 = init_io_pipe_phv_out_data_2; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_3 = init_io_pipe_phv_out_data_3; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_4 = init_io_pipe_phv_out_data_4; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_5 = init_io_pipe_phv_out_data_5; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_6 = init_io_pipe_phv_out_data_6; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_7 = init_io_pipe_phv_out_data_7; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_8 = init_io_pipe_phv_out_data_8; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_9 = init_io_pipe_phv_out_data_9; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_10 = init_io_pipe_phv_out_data_10; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_11 = init_io_pipe_phv_out_data_11; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_12 = init_io_pipe_phv_out_data_12; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_13 = init_io_pipe_phv_out_data_13; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_14 = init_io_pipe_phv_out_data_14; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_15 = init_io_pipe_phv_out_data_15; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_16 = init_io_pipe_phv_out_data_16; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_17 = init_io_pipe_phv_out_data_17; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_18 = init_io_pipe_phv_out_data_18; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_19 = init_io_pipe_phv_out_data_19; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_20 = init_io_pipe_phv_out_data_20; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_21 = init_io_pipe_phv_out_data_21; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_22 = init_io_pipe_phv_out_data_22; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_23 = init_io_pipe_phv_out_data_23; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_24 = init_io_pipe_phv_out_data_24; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_25 = init_io_pipe_phv_out_data_25; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_26 = init_io_pipe_phv_out_data_26; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_27 = init_io_pipe_phv_out_data_27; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_28 = init_io_pipe_phv_out_data_28; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_29 = init_io_pipe_phv_out_data_29; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_30 = init_io_pipe_phv_out_data_30; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_31 = init_io_pipe_phv_out_data_31; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_32 = init_io_pipe_phv_out_data_32; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_33 = init_io_pipe_phv_out_data_33; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_34 = init_io_pipe_phv_out_data_34; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_35 = init_io_pipe_phv_out_data_35; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_36 = init_io_pipe_phv_out_data_36; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_37 = init_io_pipe_phv_out_data_37; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_38 = init_io_pipe_phv_out_data_38; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_39 = init_io_pipe_phv_out_data_39; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_40 = init_io_pipe_phv_out_data_40; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_41 = init_io_pipe_phv_out_data_41; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_42 = init_io_pipe_phv_out_data_42; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_43 = init_io_pipe_phv_out_data_43; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_44 = init_io_pipe_phv_out_data_44; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_45 = init_io_pipe_phv_out_data_45; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_46 = init_io_pipe_phv_out_data_46; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_47 = init_io_pipe_phv_out_data_47; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_48 = init_io_pipe_phv_out_data_48; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_49 = init_io_pipe_phv_out_data_49; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_50 = init_io_pipe_phv_out_data_50; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_51 = init_io_pipe_phv_out_data_51; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_52 = init_io_pipe_phv_out_data_52; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_53 = init_io_pipe_phv_out_data_53; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_54 = init_io_pipe_phv_out_data_54; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_55 = init_io_pipe_phv_out_data_55; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_56 = init_io_pipe_phv_out_data_56; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_57 = init_io_pipe_phv_out_data_57; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_58 = init_io_pipe_phv_out_data_58; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_59 = init_io_pipe_phv_out_data_59; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_60 = init_io_pipe_phv_out_data_60; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_61 = init_io_pipe_phv_out_data_61; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_62 = init_io_pipe_phv_out_data_62; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_63 = init_io_pipe_phv_out_data_63; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_64 = init_io_pipe_phv_out_data_64; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_65 = init_io_pipe_phv_out_data_65; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_66 = init_io_pipe_phv_out_data_66; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_67 = init_io_pipe_phv_out_data_67; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_68 = init_io_pipe_phv_out_data_68; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_69 = init_io_pipe_phv_out_data_69; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_70 = init_io_pipe_phv_out_data_70; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_71 = init_io_pipe_phv_out_data_71; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_72 = init_io_pipe_phv_out_data_72; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_73 = init_io_pipe_phv_out_data_73; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_74 = init_io_pipe_phv_out_data_74; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_75 = init_io_pipe_phv_out_data_75; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_76 = init_io_pipe_phv_out_data_76; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_77 = init_io_pipe_phv_out_data_77; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_78 = init_io_pipe_phv_out_data_78; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_79 = init_io_pipe_phv_out_data_79; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_80 = init_io_pipe_phv_out_data_80; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_81 = init_io_pipe_phv_out_data_81; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_82 = init_io_pipe_phv_out_data_82; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_83 = init_io_pipe_phv_out_data_83; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_84 = init_io_pipe_phv_out_data_84; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_85 = init_io_pipe_phv_out_data_85; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_86 = init_io_pipe_phv_out_data_86; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_87 = init_io_pipe_phv_out_data_87; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_88 = init_io_pipe_phv_out_data_88; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_89 = init_io_pipe_phv_out_data_89; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_90 = init_io_pipe_phv_out_data_90; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_91 = init_io_pipe_phv_out_data_91; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_92 = init_io_pipe_phv_out_data_92; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_93 = init_io_pipe_phv_out_data_93; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_94 = init_io_pipe_phv_out_data_94; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_95 = init_io_pipe_phv_out_data_95; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_96 = init_io_pipe_phv_out_data_96; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_97 = init_io_pipe_phv_out_data_97; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_98 = init_io_pipe_phv_out_data_98; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_99 = init_io_pipe_phv_out_data_99; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_100 = init_io_pipe_phv_out_data_100; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_101 = init_io_pipe_phv_out_data_101; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_102 = init_io_pipe_phv_out_data_102; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_103 = init_io_pipe_phv_out_data_103; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_104 = init_io_pipe_phv_out_data_104; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_105 = init_io_pipe_phv_out_data_105; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_106 = init_io_pipe_phv_out_data_106; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_107 = init_io_pipe_phv_out_data_107; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_108 = init_io_pipe_phv_out_data_108; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_109 = init_io_pipe_phv_out_data_109; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_110 = init_io_pipe_phv_out_data_110; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_111 = init_io_pipe_phv_out_data_111; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_112 = init_io_pipe_phv_out_data_112; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_113 = init_io_pipe_phv_out_data_113; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_114 = init_io_pipe_phv_out_data_114; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_115 = init_io_pipe_phv_out_data_115; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_116 = init_io_pipe_phv_out_data_116; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_117 = init_io_pipe_phv_out_data_117; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_118 = init_io_pipe_phv_out_data_118; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_119 = init_io_pipe_phv_out_data_119; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_120 = init_io_pipe_phv_out_data_120; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_121 = init_io_pipe_phv_out_data_121; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_122 = init_io_pipe_phv_out_data_122; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_123 = init_io_pipe_phv_out_data_123; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_124 = init_io_pipe_phv_out_data_124; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_125 = init_io_pipe_phv_out_data_125; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_126 = init_io_pipe_phv_out_data_126; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_127 = init_io_pipe_phv_out_data_127; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_data_128 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_7_io_pipe_phv_in_data_129 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_7_io_pipe_phv_in_data_130 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_7_io_pipe_phv_in_data_131 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_7_io_pipe_phv_in_data_132 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_7_io_pipe_phv_in_data_133 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_7_io_pipe_phv_in_data_134 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_7_io_pipe_phv_in_data_135 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_7_io_pipe_phv_in_data_136 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_7_io_pipe_phv_in_data_137 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_7_io_pipe_phv_in_data_138 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_7_io_pipe_phv_in_data_139 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_7_io_pipe_phv_in_data_140 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_7_io_pipe_phv_in_data_141 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_7_io_pipe_phv_in_data_142 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_7_io_pipe_phv_in_data_143 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_7_io_pipe_phv_in_data_144 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_7_io_pipe_phv_in_data_145 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_7_io_pipe_phv_in_data_146 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_7_io_pipe_phv_in_data_147 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_7_io_pipe_phv_in_data_148 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_7_io_pipe_phv_in_data_149 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_7_io_pipe_phv_in_data_150 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_7_io_pipe_phv_in_data_151 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_7_io_pipe_phv_in_data_152 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_7_io_pipe_phv_in_data_153 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_7_io_pipe_phv_in_data_154 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_7_io_pipe_phv_in_data_155 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_7_io_pipe_phv_in_data_156 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_7_io_pipe_phv_in_data_157 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_7_io_pipe_phv_in_data_158 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_7_io_pipe_phv_in_data_159 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_7_io_pipe_phv_in_header_0 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_7_io_pipe_phv_in_header_1 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_7_io_pipe_phv_in_header_2 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_7_io_pipe_phv_in_header_3 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_7_io_pipe_phv_in_header_4 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_7_io_pipe_phv_in_header_5 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_7_io_pipe_phv_in_header_6 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_7_io_pipe_phv_in_header_7 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_7_io_pipe_phv_in_header_8 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_7_io_pipe_phv_in_header_9 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_7_io_pipe_phv_in_header_10 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_7_io_pipe_phv_in_header_11 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_7_io_pipe_phv_in_header_12 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_7_io_pipe_phv_in_header_13 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_7_io_pipe_phv_in_header_14 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_7_io_pipe_phv_in_header_15 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_7_io_pipe_phv_in_parse_current_state = 8'h0; // @[ipsa.scala 94:65]
  assign proc_7_io_pipe_phv_in_parse_current_offset = 8'h0; // @[ipsa.scala 94:65]
  assign proc_7_io_pipe_phv_in_parse_transition_field = 16'h0; // @[ipsa.scala 94:65]
  assign proc_7_io_pipe_phv_in_next_processor_id = 4'h0; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_next_config_id = 1'h0; // @[ipsa.scala 94:65]
  assign proc_7_io_pipe_phv_in_is_valid_processor = 1'h0; // @[ipsa.scala 94:65]
  assign proc_7_io_pipe_phv_in_valid = init_io_pipe_phv_out_valid; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_7_io_pipe_phv_in_last = init_io_pipe_phv_out_last; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_clock = clock;
  assign proc_8_io_pipe_phv_in_data_0 = init_io_pipe_phv_out_data_0; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_1 = init_io_pipe_phv_out_data_1; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_2 = init_io_pipe_phv_out_data_2; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_3 = init_io_pipe_phv_out_data_3; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_4 = init_io_pipe_phv_out_data_4; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_5 = init_io_pipe_phv_out_data_5; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_6 = init_io_pipe_phv_out_data_6; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_7 = init_io_pipe_phv_out_data_7; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_8 = init_io_pipe_phv_out_data_8; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_9 = init_io_pipe_phv_out_data_9; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_10 = init_io_pipe_phv_out_data_10; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_11 = init_io_pipe_phv_out_data_11; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_12 = init_io_pipe_phv_out_data_12; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_13 = init_io_pipe_phv_out_data_13; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_14 = init_io_pipe_phv_out_data_14; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_15 = init_io_pipe_phv_out_data_15; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_16 = init_io_pipe_phv_out_data_16; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_17 = init_io_pipe_phv_out_data_17; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_18 = init_io_pipe_phv_out_data_18; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_19 = init_io_pipe_phv_out_data_19; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_20 = init_io_pipe_phv_out_data_20; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_21 = init_io_pipe_phv_out_data_21; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_22 = init_io_pipe_phv_out_data_22; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_23 = init_io_pipe_phv_out_data_23; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_24 = init_io_pipe_phv_out_data_24; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_25 = init_io_pipe_phv_out_data_25; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_26 = init_io_pipe_phv_out_data_26; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_27 = init_io_pipe_phv_out_data_27; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_28 = init_io_pipe_phv_out_data_28; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_29 = init_io_pipe_phv_out_data_29; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_30 = init_io_pipe_phv_out_data_30; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_31 = init_io_pipe_phv_out_data_31; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_32 = init_io_pipe_phv_out_data_32; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_33 = init_io_pipe_phv_out_data_33; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_34 = init_io_pipe_phv_out_data_34; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_35 = init_io_pipe_phv_out_data_35; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_36 = init_io_pipe_phv_out_data_36; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_37 = init_io_pipe_phv_out_data_37; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_38 = init_io_pipe_phv_out_data_38; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_39 = init_io_pipe_phv_out_data_39; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_40 = init_io_pipe_phv_out_data_40; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_41 = init_io_pipe_phv_out_data_41; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_42 = init_io_pipe_phv_out_data_42; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_43 = init_io_pipe_phv_out_data_43; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_44 = init_io_pipe_phv_out_data_44; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_45 = init_io_pipe_phv_out_data_45; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_46 = init_io_pipe_phv_out_data_46; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_47 = init_io_pipe_phv_out_data_47; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_48 = init_io_pipe_phv_out_data_48; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_49 = init_io_pipe_phv_out_data_49; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_50 = init_io_pipe_phv_out_data_50; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_51 = init_io_pipe_phv_out_data_51; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_52 = init_io_pipe_phv_out_data_52; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_53 = init_io_pipe_phv_out_data_53; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_54 = init_io_pipe_phv_out_data_54; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_55 = init_io_pipe_phv_out_data_55; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_56 = init_io_pipe_phv_out_data_56; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_57 = init_io_pipe_phv_out_data_57; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_58 = init_io_pipe_phv_out_data_58; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_59 = init_io_pipe_phv_out_data_59; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_60 = init_io_pipe_phv_out_data_60; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_61 = init_io_pipe_phv_out_data_61; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_62 = init_io_pipe_phv_out_data_62; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_63 = init_io_pipe_phv_out_data_63; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_64 = init_io_pipe_phv_out_data_64; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_65 = init_io_pipe_phv_out_data_65; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_66 = init_io_pipe_phv_out_data_66; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_67 = init_io_pipe_phv_out_data_67; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_68 = init_io_pipe_phv_out_data_68; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_69 = init_io_pipe_phv_out_data_69; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_70 = init_io_pipe_phv_out_data_70; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_71 = init_io_pipe_phv_out_data_71; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_72 = init_io_pipe_phv_out_data_72; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_73 = init_io_pipe_phv_out_data_73; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_74 = init_io_pipe_phv_out_data_74; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_75 = init_io_pipe_phv_out_data_75; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_76 = init_io_pipe_phv_out_data_76; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_77 = init_io_pipe_phv_out_data_77; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_78 = init_io_pipe_phv_out_data_78; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_79 = init_io_pipe_phv_out_data_79; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_80 = init_io_pipe_phv_out_data_80; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_81 = init_io_pipe_phv_out_data_81; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_82 = init_io_pipe_phv_out_data_82; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_83 = init_io_pipe_phv_out_data_83; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_84 = init_io_pipe_phv_out_data_84; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_85 = init_io_pipe_phv_out_data_85; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_86 = init_io_pipe_phv_out_data_86; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_87 = init_io_pipe_phv_out_data_87; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_88 = init_io_pipe_phv_out_data_88; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_89 = init_io_pipe_phv_out_data_89; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_90 = init_io_pipe_phv_out_data_90; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_91 = init_io_pipe_phv_out_data_91; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_92 = init_io_pipe_phv_out_data_92; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_93 = init_io_pipe_phv_out_data_93; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_94 = init_io_pipe_phv_out_data_94; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_95 = init_io_pipe_phv_out_data_95; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_96 = init_io_pipe_phv_out_data_96; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_97 = init_io_pipe_phv_out_data_97; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_98 = init_io_pipe_phv_out_data_98; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_99 = init_io_pipe_phv_out_data_99; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_100 = init_io_pipe_phv_out_data_100; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_101 = init_io_pipe_phv_out_data_101; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_102 = init_io_pipe_phv_out_data_102; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_103 = init_io_pipe_phv_out_data_103; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_104 = init_io_pipe_phv_out_data_104; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_105 = init_io_pipe_phv_out_data_105; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_106 = init_io_pipe_phv_out_data_106; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_107 = init_io_pipe_phv_out_data_107; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_108 = init_io_pipe_phv_out_data_108; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_109 = init_io_pipe_phv_out_data_109; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_110 = init_io_pipe_phv_out_data_110; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_111 = init_io_pipe_phv_out_data_111; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_112 = init_io_pipe_phv_out_data_112; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_113 = init_io_pipe_phv_out_data_113; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_114 = init_io_pipe_phv_out_data_114; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_115 = init_io_pipe_phv_out_data_115; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_116 = init_io_pipe_phv_out_data_116; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_117 = init_io_pipe_phv_out_data_117; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_118 = init_io_pipe_phv_out_data_118; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_119 = init_io_pipe_phv_out_data_119; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_120 = init_io_pipe_phv_out_data_120; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_121 = init_io_pipe_phv_out_data_121; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_122 = init_io_pipe_phv_out_data_122; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_123 = init_io_pipe_phv_out_data_123; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_124 = init_io_pipe_phv_out_data_124; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_125 = init_io_pipe_phv_out_data_125; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_126 = init_io_pipe_phv_out_data_126; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_127 = init_io_pipe_phv_out_data_127; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_data_128 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_8_io_pipe_phv_in_data_129 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_8_io_pipe_phv_in_data_130 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_8_io_pipe_phv_in_data_131 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_8_io_pipe_phv_in_data_132 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_8_io_pipe_phv_in_data_133 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_8_io_pipe_phv_in_data_134 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_8_io_pipe_phv_in_data_135 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_8_io_pipe_phv_in_data_136 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_8_io_pipe_phv_in_data_137 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_8_io_pipe_phv_in_data_138 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_8_io_pipe_phv_in_data_139 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_8_io_pipe_phv_in_data_140 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_8_io_pipe_phv_in_data_141 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_8_io_pipe_phv_in_data_142 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_8_io_pipe_phv_in_data_143 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_8_io_pipe_phv_in_data_144 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_8_io_pipe_phv_in_data_145 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_8_io_pipe_phv_in_data_146 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_8_io_pipe_phv_in_data_147 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_8_io_pipe_phv_in_data_148 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_8_io_pipe_phv_in_data_149 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_8_io_pipe_phv_in_data_150 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_8_io_pipe_phv_in_data_151 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_8_io_pipe_phv_in_data_152 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_8_io_pipe_phv_in_data_153 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_8_io_pipe_phv_in_data_154 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_8_io_pipe_phv_in_data_155 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_8_io_pipe_phv_in_data_156 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_8_io_pipe_phv_in_data_157 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_8_io_pipe_phv_in_data_158 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_8_io_pipe_phv_in_data_159 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_8_io_pipe_phv_in_header_0 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_8_io_pipe_phv_in_header_1 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_8_io_pipe_phv_in_header_2 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_8_io_pipe_phv_in_header_3 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_8_io_pipe_phv_in_header_4 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_8_io_pipe_phv_in_header_5 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_8_io_pipe_phv_in_header_6 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_8_io_pipe_phv_in_header_7 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_8_io_pipe_phv_in_header_8 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_8_io_pipe_phv_in_header_9 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_8_io_pipe_phv_in_header_10 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_8_io_pipe_phv_in_header_11 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_8_io_pipe_phv_in_header_12 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_8_io_pipe_phv_in_header_13 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_8_io_pipe_phv_in_header_14 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_8_io_pipe_phv_in_header_15 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_8_io_pipe_phv_in_parse_current_state = 8'h0; // @[ipsa.scala 94:65]
  assign proc_8_io_pipe_phv_in_parse_current_offset = 8'h0; // @[ipsa.scala 94:65]
  assign proc_8_io_pipe_phv_in_parse_transition_field = 16'h0; // @[ipsa.scala 94:65]
  assign proc_8_io_pipe_phv_in_next_processor_id = 4'h0; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_next_config_id = 1'h0; // @[ipsa.scala 94:65]
  assign proc_8_io_pipe_phv_in_is_valid_processor = 1'h0; // @[ipsa.scala 94:65]
  assign proc_8_io_pipe_phv_in_valid = init_io_pipe_phv_out_valid; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_8_io_pipe_phv_in_last = init_io_pipe_phv_out_last; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_clock = clock;
  assign proc_9_io_pipe_phv_in_data_0 = init_io_pipe_phv_out_data_0; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_1 = init_io_pipe_phv_out_data_1; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_2 = init_io_pipe_phv_out_data_2; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_3 = init_io_pipe_phv_out_data_3; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_4 = init_io_pipe_phv_out_data_4; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_5 = init_io_pipe_phv_out_data_5; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_6 = init_io_pipe_phv_out_data_6; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_7 = init_io_pipe_phv_out_data_7; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_8 = init_io_pipe_phv_out_data_8; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_9 = init_io_pipe_phv_out_data_9; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_10 = init_io_pipe_phv_out_data_10; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_11 = init_io_pipe_phv_out_data_11; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_12 = init_io_pipe_phv_out_data_12; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_13 = init_io_pipe_phv_out_data_13; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_14 = init_io_pipe_phv_out_data_14; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_15 = init_io_pipe_phv_out_data_15; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_16 = init_io_pipe_phv_out_data_16; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_17 = init_io_pipe_phv_out_data_17; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_18 = init_io_pipe_phv_out_data_18; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_19 = init_io_pipe_phv_out_data_19; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_20 = init_io_pipe_phv_out_data_20; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_21 = init_io_pipe_phv_out_data_21; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_22 = init_io_pipe_phv_out_data_22; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_23 = init_io_pipe_phv_out_data_23; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_24 = init_io_pipe_phv_out_data_24; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_25 = init_io_pipe_phv_out_data_25; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_26 = init_io_pipe_phv_out_data_26; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_27 = init_io_pipe_phv_out_data_27; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_28 = init_io_pipe_phv_out_data_28; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_29 = init_io_pipe_phv_out_data_29; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_30 = init_io_pipe_phv_out_data_30; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_31 = init_io_pipe_phv_out_data_31; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_32 = init_io_pipe_phv_out_data_32; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_33 = init_io_pipe_phv_out_data_33; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_34 = init_io_pipe_phv_out_data_34; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_35 = init_io_pipe_phv_out_data_35; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_36 = init_io_pipe_phv_out_data_36; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_37 = init_io_pipe_phv_out_data_37; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_38 = init_io_pipe_phv_out_data_38; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_39 = init_io_pipe_phv_out_data_39; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_40 = init_io_pipe_phv_out_data_40; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_41 = init_io_pipe_phv_out_data_41; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_42 = init_io_pipe_phv_out_data_42; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_43 = init_io_pipe_phv_out_data_43; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_44 = init_io_pipe_phv_out_data_44; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_45 = init_io_pipe_phv_out_data_45; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_46 = init_io_pipe_phv_out_data_46; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_47 = init_io_pipe_phv_out_data_47; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_48 = init_io_pipe_phv_out_data_48; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_49 = init_io_pipe_phv_out_data_49; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_50 = init_io_pipe_phv_out_data_50; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_51 = init_io_pipe_phv_out_data_51; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_52 = init_io_pipe_phv_out_data_52; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_53 = init_io_pipe_phv_out_data_53; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_54 = init_io_pipe_phv_out_data_54; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_55 = init_io_pipe_phv_out_data_55; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_56 = init_io_pipe_phv_out_data_56; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_57 = init_io_pipe_phv_out_data_57; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_58 = init_io_pipe_phv_out_data_58; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_59 = init_io_pipe_phv_out_data_59; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_60 = init_io_pipe_phv_out_data_60; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_61 = init_io_pipe_phv_out_data_61; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_62 = init_io_pipe_phv_out_data_62; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_63 = init_io_pipe_phv_out_data_63; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_64 = init_io_pipe_phv_out_data_64; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_65 = init_io_pipe_phv_out_data_65; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_66 = init_io_pipe_phv_out_data_66; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_67 = init_io_pipe_phv_out_data_67; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_68 = init_io_pipe_phv_out_data_68; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_69 = init_io_pipe_phv_out_data_69; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_70 = init_io_pipe_phv_out_data_70; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_71 = init_io_pipe_phv_out_data_71; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_72 = init_io_pipe_phv_out_data_72; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_73 = init_io_pipe_phv_out_data_73; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_74 = init_io_pipe_phv_out_data_74; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_75 = init_io_pipe_phv_out_data_75; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_76 = init_io_pipe_phv_out_data_76; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_77 = init_io_pipe_phv_out_data_77; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_78 = init_io_pipe_phv_out_data_78; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_79 = init_io_pipe_phv_out_data_79; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_80 = init_io_pipe_phv_out_data_80; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_81 = init_io_pipe_phv_out_data_81; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_82 = init_io_pipe_phv_out_data_82; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_83 = init_io_pipe_phv_out_data_83; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_84 = init_io_pipe_phv_out_data_84; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_85 = init_io_pipe_phv_out_data_85; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_86 = init_io_pipe_phv_out_data_86; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_87 = init_io_pipe_phv_out_data_87; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_88 = init_io_pipe_phv_out_data_88; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_89 = init_io_pipe_phv_out_data_89; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_90 = init_io_pipe_phv_out_data_90; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_91 = init_io_pipe_phv_out_data_91; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_92 = init_io_pipe_phv_out_data_92; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_93 = init_io_pipe_phv_out_data_93; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_94 = init_io_pipe_phv_out_data_94; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_95 = init_io_pipe_phv_out_data_95; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_96 = init_io_pipe_phv_out_data_96; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_97 = init_io_pipe_phv_out_data_97; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_98 = init_io_pipe_phv_out_data_98; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_99 = init_io_pipe_phv_out_data_99; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_100 = init_io_pipe_phv_out_data_100; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_101 = init_io_pipe_phv_out_data_101; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_102 = init_io_pipe_phv_out_data_102; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_103 = init_io_pipe_phv_out_data_103; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_104 = init_io_pipe_phv_out_data_104; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_105 = init_io_pipe_phv_out_data_105; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_106 = init_io_pipe_phv_out_data_106; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_107 = init_io_pipe_phv_out_data_107; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_108 = init_io_pipe_phv_out_data_108; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_109 = init_io_pipe_phv_out_data_109; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_110 = init_io_pipe_phv_out_data_110; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_111 = init_io_pipe_phv_out_data_111; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_112 = init_io_pipe_phv_out_data_112; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_113 = init_io_pipe_phv_out_data_113; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_114 = init_io_pipe_phv_out_data_114; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_115 = init_io_pipe_phv_out_data_115; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_116 = init_io_pipe_phv_out_data_116; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_117 = init_io_pipe_phv_out_data_117; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_118 = init_io_pipe_phv_out_data_118; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_119 = init_io_pipe_phv_out_data_119; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_120 = init_io_pipe_phv_out_data_120; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_121 = init_io_pipe_phv_out_data_121; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_122 = init_io_pipe_phv_out_data_122; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_123 = init_io_pipe_phv_out_data_123; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_124 = init_io_pipe_phv_out_data_124; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_125 = init_io_pipe_phv_out_data_125; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_126 = init_io_pipe_phv_out_data_126; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_127 = init_io_pipe_phv_out_data_127; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_data_128 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_9_io_pipe_phv_in_data_129 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_9_io_pipe_phv_in_data_130 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_9_io_pipe_phv_in_data_131 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_9_io_pipe_phv_in_data_132 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_9_io_pipe_phv_in_data_133 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_9_io_pipe_phv_in_data_134 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_9_io_pipe_phv_in_data_135 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_9_io_pipe_phv_in_data_136 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_9_io_pipe_phv_in_data_137 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_9_io_pipe_phv_in_data_138 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_9_io_pipe_phv_in_data_139 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_9_io_pipe_phv_in_data_140 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_9_io_pipe_phv_in_data_141 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_9_io_pipe_phv_in_data_142 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_9_io_pipe_phv_in_data_143 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_9_io_pipe_phv_in_data_144 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_9_io_pipe_phv_in_data_145 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_9_io_pipe_phv_in_data_146 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_9_io_pipe_phv_in_data_147 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_9_io_pipe_phv_in_data_148 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_9_io_pipe_phv_in_data_149 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_9_io_pipe_phv_in_data_150 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_9_io_pipe_phv_in_data_151 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_9_io_pipe_phv_in_data_152 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_9_io_pipe_phv_in_data_153 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_9_io_pipe_phv_in_data_154 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_9_io_pipe_phv_in_data_155 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_9_io_pipe_phv_in_data_156 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_9_io_pipe_phv_in_data_157 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_9_io_pipe_phv_in_data_158 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_9_io_pipe_phv_in_data_159 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_9_io_pipe_phv_in_header_0 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_9_io_pipe_phv_in_header_1 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_9_io_pipe_phv_in_header_2 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_9_io_pipe_phv_in_header_3 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_9_io_pipe_phv_in_header_4 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_9_io_pipe_phv_in_header_5 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_9_io_pipe_phv_in_header_6 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_9_io_pipe_phv_in_header_7 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_9_io_pipe_phv_in_header_8 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_9_io_pipe_phv_in_header_9 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_9_io_pipe_phv_in_header_10 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_9_io_pipe_phv_in_header_11 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_9_io_pipe_phv_in_header_12 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_9_io_pipe_phv_in_header_13 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_9_io_pipe_phv_in_header_14 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_9_io_pipe_phv_in_header_15 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_9_io_pipe_phv_in_parse_current_state = 8'h0; // @[ipsa.scala 94:65]
  assign proc_9_io_pipe_phv_in_parse_current_offset = 8'h0; // @[ipsa.scala 94:65]
  assign proc_9_io_pipe_phv_in_parse_transition_field = 16'h0; // @[ipsa.scala 94:65]
  assign proc_9_io_pipe_phv_in_next_processor_id = 4'h0; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_next_config_id = 1'h0; // @[ipsa.scala 94:65]
  assign proc_9_io_pipe_phv_in_is_valid_processor = 1'h0; // @[ipsa.scala 94:65]
  assign proc_9_io_pipe_phv_in_valid = init_io_pipe_phv_out_valid; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_9_io_pipe_phv_in_last = init_io_pipe_phv_out_last; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_clock = clock;
  assign proc_10_io_pipe_phv_in_data_0 = init_io_pipe_phv_out_data_0; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_1 = init_io_pipe_phv_out_data_1; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_2 = init_io_pipe_phv_out_data_2; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_3 = init_io_pipe_phv_out_data_3; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_4 = init_io_pipe_phv_out_data_4; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_5 = init_io_pipe_phv_out_data_5; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_6 = init_io_pipe_phv_out_data_6; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_7 = init_io_pipe_phv_out_data_7; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_8 = init_io_pipe_phv_out_data_8; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_9 = init_io_pipe_phv_out_data_9; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_10 = init_io_pipe_phv_out_data_10; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_11 = init_io_pipe_phv_out_data_11; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_12 = init_io_pipe_phv_out_data_12; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_13 = init_io_pipe_phv_out_data_13; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_14 = init_io_pipe_phv_out_data_14; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_15 = init_io_pipe_phv_out_data_15; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_16 = init_io_pipe_phv_out_data_16; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_17 = init_io_pipe_phv_out_data_17; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_18 = init_io_pipe_phv_out_data_18; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_19 = init_io_pipe_phv_out_data_19; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_20 = init_io_pipe_phv_out_data_20; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_21 = init_io_pipe_phv_out_data_21; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_22 = init_io_pipe_phv_out_data_22; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_23 = init_io_pipe_phv_out_data_23; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_24 = init_io_pipe_phv_out_data_24; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_25 = init_io_pipe_phv_out_data_25; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_26 = init_io_pipe_phv_out_data_26; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_27 = init_io_pipe_phv_out_data_27; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_28 = init_io_pipe_phv_out_data_28; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_29 = init_io_pipe_phv_out_data_29; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_30 = init_io_pipe_phv_out_data_30; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_31 = init_io_pipe_phv_out_data_31; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_32 = init_io_pipe_phv_out_data_32; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_33 = init_io_pipe_phv_out_data_33; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_34 = init_io_pipe_phv_out_data_34; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_35 = init_io_pipe_phv_out_data_35; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_36 = init_io_pipe_phv_out_data_36; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_37 = init_io_pipe_phv_out_data_37; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_38 = init_io_pipe_phv_out_data_38; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_39 = init_io_pipe_phv_out_data_39; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_40 = init_io_pipe_phv_out_data_40; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_41 = init_io_pipe_phv_out_data_41; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_42 = init_io_pipe_phv_out_data_42; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_43 = init_io_pipe_phv_out_data_43; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_44 = init_io_pipe_phv_out_data_44; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_45 = init_io_pipe_phv_out_data_45; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_46 = init_io_pipe_phv_out_data_46; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_47 = init_io_pipe_phv_out_data_47; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_48 = init_io_pipe_phv_out_data_48; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_49 = init_io_pipe_phv_out_data_49; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_50 = init_io_pipe_phv_out_data_50; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_51 = init_io_pipe_phv_out_data_51; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_52 = init_io_pipe_phv_out_data_52; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_53 = init_io_pipe_phv_out_data_53; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_54 = init_io_pipe_phv_out_data_54; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_55 = init_io_pipe_phv_out_data_55; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_56 = init_io_pipe_phv_out_data_56; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_57 = init_io_pipe_phv_out_data_57; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_58 = init_io_pipe_phv_out_data_58; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_59 = init_io_pipe_phv_out_data_59; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_60 = init_io_pipe_phv_out_data_60; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_61 = init_io_pipe_phv_out_data_61; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_62 = init_io_pipe_phv_out_data_62; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_63 = init_io_pipe_phv_out_data_63; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_64 = init_io_pipe_phv_out_data_64; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_65 = init_io_pipe_phv_out_data_65; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_66 = init_io_pipe_phv_out_data_66; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_67 = init_io_pipe_phv_out_data_67; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_68 = init_io_pipe_phv_out_data_68; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_69 = init_io_pipe_phv_out_data_69; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_70 = init_io_pipe_phv_out_data_70; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_71 = init_io_pipe_phv_out_data_71; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_72 = init_io_pipe_phv_out_data_72; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_73 = init_io_pipe_phv_out_data_73; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_74 = init_io_pipe_phv_out_data_74; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_75 = init_io_pipe_phv_out_data_75; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_76 = init_io_pipe_phv_out_data_76; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_77 = init_io_pipe_phv_out_data_77; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_78 = init_io_pipe_phv_out_data_78; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_79 = init_io_pipe_phv_out_data_79; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_80 = init_io_pipe_phv_out_data_80; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_81 = init_io_pipe_phv_out_data_81; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_82 = init_io_pipe_phv_out_data_82; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_83 = init_io_pipe_phv_out_data_83; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_84 = init_io_pipe_phv_out_data_84; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_85 = init_io_pipe_phv_out_data_85; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_86 = init_io_pipe_phv_out_data_86; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_87 = init_io_pipe_phv_out_data_87; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_88 = init_io_pipe_phv_out_data_88; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_89 = init_io_pipe_phv_out_data_89; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_90 = init_io_pipe_phv_out_data_90; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_91 = init_io_pipe_phv_out_data_91; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_92 = init_io_pipe_phv_out_data_92; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_93 = init_io_pipe_phv_out_data_93; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_94 = init_io_pipe_phv_out_data_94; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_95 = init_io_pipe_phv_out_data_95; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_96 = init_io_pipe_phv_out_data_96; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_97 = init_io_pipe_phv_out_data_97; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_98 = init_io_pipe_phv_out_data_98; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_99 = init_io_pipe_phv_out_data_99; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_100 = init_io_pipe_phv_out_data_100; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_101 = init_io_pipe_phv_out_data_101; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_102 = init_io_pipe_phv_out_data_102; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_103 = init_io_pipe_phv_out_data_103; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_104 = init_io_pipe_phv_out_data_104; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_105 = init_io_pipe_phv_out_data_105; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_106 = init_io_pipe_phv_out_data_106; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_107 = init_io_pipe_phv_out_data_107; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_108 = init_io_pipe_phv_out_data_108; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_109 = init_io_pipe_phv_out_data_109; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_110 = init_io_pipe_phv_out_data_110; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_111 = init_io_pipe_phv_out_data_111; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_112 = init_io_pipe_phv_out_data_112; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_113 = init_io_pipe_phv_out_data_113; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_114 = init_io_pipe_phv_out_data_114; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_115 = init_io_pipe_phv_out_data_115; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_116 = init_io_pipe_phv_out_data_116; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_117 = init_io_pipe_phv_out_data_117; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_118 = init_io_pipe_phv_out_data_118; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_119 = init_io_pipe_phv_out_data_119; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_120 = init_io_pipe_phv_out_data_120; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_121 = init_io_pipe_phv_out_data_121; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_122 = init_io_pipe_phv_out_data_122; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_123 = init_io_pipe_phv_out_data_123; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_124 = init_io_pipe_phv_out_data_124; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_125 = init_io_pipe_phv_out_data_125; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_126 = init_io_pipe_phv_out_data_126; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_127 = init_io_pipe_phv_out_data_127; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_data_128 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_10_io_pipe_phv_in_data_129 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_10_io_pipe_phv_in_data_130 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_10_io_pipe_phv_in_data_131 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_10_io_pipe_phv_in_data_132 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_10_io_pipe_phv_in_data_133 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_10_io_pipe_phv_in_data_134 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_10_io_pipe_phv_in_data_135 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_10_io_pipe_phv_in_data_136 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_10_io_pipe_phv_in_data_137 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_10_io_pipe_phv_in_data_138 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_10_io_pipe_phv_in_data_139 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_10_io_pipe_phv_in_data_140 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_10_io_pipe_phv_in_data_141 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_10_io_pipe_phv_in_data_142 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_10_io_pipe_phv_in_data_143 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_10_io_pipe_phv_in_data_144 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_10_io_pipe_phv_in_data_145 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_10_io_pipe_phv_in_data_146 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_10_io_pipe_phv_in_data_147 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_10_io_pipe_phv_in_data_148 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_10_io_pipe_phv_in_data_149 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_10_io_pipe_phv_in_data_150 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_10_io_pipe_phv_in_data_151 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_10_io_pipe_phv_in_data_152 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_10_io_pipe_phv_in_data_153 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_10_io_pipe_phv_in_data_154 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_10_io_pipe_phv_in_data_155 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_10_io_pipe_phv_in_data_156 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_10_io_pipe_phv_in_data_157 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_10_io_pipe_phv_in_data_158 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_10_io_pipe_phv_in_data_159 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_10_io_pipe_phv_in_header_0 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_10_io_pipe_phv_in_header_1 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_10_io_pipe_phv_in_header_2 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_10_io_pipe_phv_in_header_3 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_10_io_pipe_phv_in_header_4 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_10_io_pipe_phv_in_header_5 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_10_io_pipe_phv_in_header_6 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_10_io_pipe_phv_in_header_7 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_10_io_pipe_phv_in_header_8 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_10_io_pipe_phv_in_header_9 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_10_io_pipe_phv_in_header_10 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_10_io_pipe_phv_in_header_11 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_10_io_pipe_phv_in_header_12 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_10_io_pipe_phv_in_header_13 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_10_io_pipe_phv_in_header_14 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_10_io_pipe_phv_in_header_15 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_10_io_pipe_phv_in_parse_current_state = 8'h0; // @[ipsa.scala 94:65]
  assign proc_10_io_pipe_phv_in_parse_current_offset = 8'h0; // @[ipsa.scala 94:65]
  assign proc_10_io_pipe_phv_in_parse_transition_field = 16'h0; // @[ipsa.scala 94:65]
  assign proc_10_io_pipe_phv_in_next_processor_id = 4'h0; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_next_config_id = 1'h0; // @[ipsa.scala 94:65]
  assign proc_10_io_pipe_phv_in_is_valid_processor = 1'h0; // @[ipsa.scala 94:65]
  assign proc_10_io_pipe_phv_in_valid = init_io_pipe_phv_out_valid; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_10_io_pipe_phv_in_last = init_io_pipe_phv_out_last; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_clock = clock;
  assign proc_11_io_pipe_phv_in_data_0 = init_io_pipe_phv_out_data_0; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_1 = init_io_pipe_phv_out_data_1; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_2 = init_io_pipe_phv_out_data_2; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_3 = init_io_pipe_phv_out_data_3; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_4 = init_io_pipe_phv_out_data_4; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_5 = init_io_pipe_phv_out_data_5; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_6 = init_io_pipe_phv_out_data_6; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_7 = init_io_pipe_phv_out_data_7; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_8 = init_io_pipe_phv_out_data_8; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_9 = init_io_pipe_phv_out_data_9; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_10 = init_io_pipe_phv_out_data_10; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_11 = init_io_pipe_phv_out_data_11; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_12 = init_io_pipe_phv_out_data_12; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_13 = init_io_pipe_phv_out_data_13; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_14 = init_io_pipe_phv_out_data_14; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_15 = init_io_pipe_phv_out_data_15; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_16 = init_io_pipe_phv_out_data_16; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_17 = init_io_pipe_phv_out_data_17; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_18 = init_io_pipe_phv_out_data_18; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_19 = init_io_pipe_phv_out_data_19; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_20 = init_io_pipe_phv_out_data_20; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_21 = init_io_pipe_phv_out_data_21; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_22 = init_io_pipe_phv_out_data_22; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_23 = init_io_pipe_phv_out_data_23; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_24 = init_io_pipe_phv_out_data_24; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_25 = init_io_pipe_phv_out_data_25; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_26 = init_io_pipe_phv_out_data_26; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_27 = init_io_pipe_phv_out_data_27; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_28 = init_io_pipe_phv_out_data_28; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_29 = init_io_pipe_phv_out_data_29; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_30 = init_io_pipe_phv_out_data_30; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_31 = init_io_pipe_phv_out_data_31; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_32 = init_io_pipe_phv_out_data_32; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_33 = init_io_pipe_phv_out_data_33; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_34 = init_io_pipe_phv_out_data_34; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_35 = init_io_pipe_phv_out_data_35; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_36 = init_io_pipe_phv_out_data_36; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_37 = init_io_pipe_phv_out_data_37; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_38 = init_io_pipe_phv_out_data_38; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_39 = init_io_pipe_phv_out_data_39; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_40 = init_io_pipe_phv_out_data_40; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_41 = init_io_pipe_phv_out_data_41; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_42 = init_io_pipe_phv_out_data_42; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_43 = init_io_pipe_phv_out_data_43; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_44 = init_io_pipe_phv_out_data_44; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_45 = init_io_pipe_phv_out_data_45; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_46 = init_io_pipe_phv_out_data_46; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_47 = init_io_pipe_phv_out_data_47; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_48 = init_io_pipe_phv_out_data_48; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_49 = init_io_pipe_phv_out_data_49; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_50 = init_io_pipe_phv_out_data_50; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_51 = init_io_pipe_phv_out_data_51; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_52 = init_io_pipe_phv_out_data_52; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_53 = init_io_pipe_phv_out_data_53; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_54 = init_io_pipe_phv_out_data_54; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_55 = init_io_pipe_phv_out_data_55; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_56 = init_io_pipe_phv_out_data_56; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_57 = init_io_pipe_phv_out_data_57; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_58 = init_io_pipe_phv_out_data_58; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_59 = init_io_pipe_phv_out_data_59; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_60 = init_io_pipe_phv_out_data_60; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_61 = init_io_pipe_phv_out_data_61; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_62 = init_io_pipe_phv_out_data_62; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_63 = init_io_pipe_phv_out_data_63; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_64 = init_io_pipe_phv_out_data_64; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_65 = init_io_pipe_phv_out_data_65; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_66 = init_io_pipe_phv_out_data_66; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_67 = init_io_pipe_phv_out_data_67; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_68 = init_io_pipe_phv_out_data_68; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_69 = init_io_pipe_phv_out_data_69; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_70 = init_io_pipe_phv_out_data_70; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_71 = init_io_pipe_phv_out_data_71; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_72 = init_io_pipe_phv_out_data_72; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_73 = init_io_pipe_phv_out_data_73; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_74 = init_io_pipe_phv_out_data_74; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_75 = init_io_pipe_phv_out_data_75; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_76 = init_io_pipe_phv_out_data_76; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_77 = init_io_pipe_phv_out_data_77; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_78 = init_io_pipe_phv_out_data_78; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_79 = init_io_pipe_phv_out_data_79; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_80 = init_io_pipe_phv_out_data_80; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_81 = init_io_pipe_phv_out_data_81; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_82 = init_io_pipe_phv_out_data_82; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_83 = init_io_pipe_phv_out_data_83; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_84 = init_io_pipe_phv_out_data_84; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_85 = init_io_pipe_phv_out_data_85; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_86 = init_io_pipe_phv_out_data_86; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_87 = init_io_pipe_phv_out_data_87; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_88 = init_io_pipe_phv_out_data_88; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_89 = init_io_pipe_phv_out_data_89; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_90 = init_io_pipe_phv_out_data_90; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_91 = init_io_pipe_phv_out_data_91; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_92 = init_io_pipe_phv_out_data_92; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_93 = init_io_pipe_phv_out_data_93; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_94 = init_io_pipe_phv_out_data_94; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_95 = init_io_pipe_phv_out_data_95; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_96 = init_io_pipe_phv_out_data_96; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_97 = init_io_pipe_phv_out_data_97; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_98 = init_io_pipe_phv_out_data_98; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_99 = init_io_pipe_phv_out_data_99; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_100 = init_io_pipe_phv_out_data_100; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_101 = init_io_pipe_phv_out_data_101; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_102 = init_io_pipe_phv_out_data_102; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_103 = init_io_pipe_phv_out_data_103; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_104 = init_io_pipe_phv_out_data_104; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_105 = init_io_pipe_phv_out_data_105; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_106 = init_io_pipe_phv_out_data_106; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_107 = init_io_pipe_phv_out_data_107; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_108 = init_io_pipe_phv_out_data_108; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_109 = init_io_pipe_phv_out_data_109; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_110 = init_io_pipe_phv_out_data_110; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_111 = init_io_pipe_phv_out_data_111; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_112 = init_io_pipe_phv_out_data_112; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_113 = init_io_pipe_phv_out_data_113; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_114 = init_io_pipe_phv_out_data_114; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_115 = init_io_pipe_phv_out_data_115; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_116 = init_io_pipe_phv_out_data_116; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_117 = init_io_pipe_phv_out_data_117; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_118 = init_io_pipe_phv_out_data_118; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_119 = init_io_pipe_phv_out_data_119; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_120 = init_io_pipe_phv_out_data_120; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_121 = init_io_pipe_phv_out_data_121; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_122 = init_io_pipe_phv_out_data_122; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_123 = init_io_pipe_phv_out_data_123; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_124 = init_io_pipe_phv_out_data_124; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_125 = init_io_pipe_phv_out_data_125; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_126 = init_io_pipe_phv_out_data_126; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_127 = init_io_pipe_phv_out_data_127; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_data_128 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_11_io_pipe_phv_in_data_129 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_11_io_pipe_phv_in_data_130 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_11_io_pipe_phv_in_data_131 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_11_io_pipe_phv_in_data_132 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_11_io_pipe_phv_in_data_133 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_11_io_pipe_phv_in_data_134 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_11_io_pipe_phv_in_data_135 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_11_io_pipe_phv_in_data_136 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_11_io_pipe_phv_in_data_137 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_11_io_pipe_phv_in_data_138 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_11_io_pipe_phv_in_data_139 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_11_io_pipe_phv_in_data_140 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_11_io_pipe_phv_in_data_141 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_11_io_pipe_phv_in_data_142 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_11_io_pipe_phv_in_data_143 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_11_io_pipe_phv_in_data_144 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_11_io_pipe_phv_in_data_145 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_11_io_pipe_phv_in_data_146 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_11_io_pipe_phv_in_data_147 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_11_io_pipe_phv_in_data_148 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_11_io_pipe_phv_in_data_149 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_11_io_pipe_phv_in_data_150 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_11_io_pipe_phv_in_data_151 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_11_io_pipe_phv_in_data_152 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_11_io_pipe_phv_in_data_153 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_11_io_pipe_phv_in_data_154 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_11_io_pipe_phv_in_data_155 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_11_io_pipe_phv_in_data_156 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_11_io_pipe_phv_in_data_157 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_11_io_pipe_phv_in_data_158 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_11_io_pipe_phv_in_data_159 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_11_io_pipe_phv_in_header_0 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_11_io_pipe_phv_in_header_1 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_11_io_pipe_phv_in_header_2 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_11_io_pipe_phv_in_header_3 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_11_io_pipe_phv_in_header_4 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_11_io_pipe_phv_in_header_5 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_11_io_pipe_phv_in_header_6 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_11_io_pipe_phv_in_header_7 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_11_io_pipe_phv_in_header_8 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_11_io_pipe_phv_in_header_9 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_11_io_pipe_phv_in_header_10 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_11_io_pipe_phv_in_header_11 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_11_io_pipe_phv_in_header_12 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_11_io_pipe_phv_in_header_13 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_11_io_pipe_phv_in_header_14 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_11_io_pipe_phv_in_header_15 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_11_io_pipe_phv_in_parse_current_state = 8'h0; // @[ipsa.scala 94:65]
  assign proc_11_io_pipe_phv_in_parse_current_offset = 8'h0; // @[ipsa.scala 94:65]
  assign proc_11_io_pipe_phv_in_parse_transition_field = 16'h0; // @[ipsa.scala 94:65]
  assign proc_11_io_pipe_phv_in_next_processor_id = 4'h0; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_next_config_id = 1'h0; // @[ipsa.scala 94:65]
  assign proc_11_io_pipe_phv_in_is_valid_processor = 1'h0; // @[ipsa.scala 94:65]
  assign proc_11_io_pipe_phv_in_valid = init_io_pipe_phv_out_valid; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_11_io_pipe_phv_in_last = init_io_pipe_phv_out_last; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_clock = clock;
  assign proc_12_io_pipe_phv_in_data_0 = init_io_pipe_phv_out_data_0; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_1 = init_io_pipe_phv_out_data_1; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_2 = init_io_pipe_phv_out_data_2; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_3 = init_io_pipe_phv_out_data_3; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_4 = init_io_pipe_phv_out_data_4; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_5 = init_io_pipe_phv_out_data_5; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_6 = init_io_pipe_phv_out_data_6; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_7 = init_io_pipe_phv_out_data_7; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_8 = init_io_pipe_phv_out_data_8; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_9 = init_io_pipe_phv_out_data_9; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_10 = init_io_pipe_phv_out_data_10; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_11 = init_io_pipe_phv_out_data_11; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_12 = init_io_pipe_phv_out_data_12; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_13 = init_io_pipe_phv_out_data_13; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_14 = init_io_pipe_phv_out_data_14; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_15 = init_io_pipe_phv_out_data_15; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_16 = init_io_pipe_phv_out_data_16; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_17 = init_io_pipe_phv_out_data_17; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_18 = init_io_pipe_phv_out_data_18; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_19 = init_io_pipe_phv_out_data_19; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_20 = init_io_pipe_phv_out_data_20; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_21 = init_io_pipe_phv_out_data_21; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_22 = init_io_pipe_phv_out_data_22; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_23 = init_io_pipe_phv_out_data_23; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_24 = init_io_pipe_phv_out_data_24; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_25 = init_io_pipe_phv_out_data_25; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_26 = init_io_pipe_phv_out_data_26; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_27 = init_io_pipe_phv_out_data_27; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_28 = init_io_pipe_phv_out_data_28; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_29 = init_io_pipe_phv_out_data_29; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_30 = init_io_pipe_phv_out_data_30; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_31 = init_io_pipe_phv_out_data_31; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_32 = init_io_pipe_phv_out_data_32; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_33 = init_io_pipe_phv_out_data_33; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_34 = init_io_pipe_phv_out_data_34; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_35 = init_io_pipe_phv_out_data_35; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_36 = init_io_pipe_phv_out_data_36; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_37 = init_io_pipe_phv_out_data_37; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_38 = init_io_pipe_phv_out_data_38; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_39 = init_io_pipe_phv_out_data_39; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_40 = init_io_pipe_phv_out_data_40; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_41 = init_io_pipe_phv_out_data_41; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_42 = init_io_pipe_phv_out_data_42; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_43 = init_io_pipe_phv_out_data_43; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_44 = init_io_pipe_phv_out_data_44; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_45 = init_io_pipe_phv_out_data_45; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_46 = init_io_pipe_phv_out_data_46; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_47 = init_io_pipe_phv_out_data_47; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_48 = init_io_pipe_phv_out_data_48; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_49 = init_io_pipe_phv_out_data_49; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_50 = init_io_pipe_phv_out_data_50; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_51 = init_io_pipe_phv_out_data_51; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_52 = init_io_pipe_phv_out_data_52; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_53 = init_io_pipe_phv_out_data_53; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_54 = init_io_pipe_phv_out_data_54; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_55 = init_io_pipe_phv_out_data_55; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_56 = init_io_pipe_phv_out_data_56; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_57 = init_io_pipe_phv_out_data_57; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_58 = init_io_pipe_phv_out_data_58; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_59 = init_io_pipe_phv_out_data_59; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_60 = init_io_pipe_phv_out_data_60; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_61 = init_io_pipe_phv_out_data_61; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_62 = init_io_pipe_phv_out_data_62; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_63 = init_io_pipe_phv_out_data_63; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_64 = init_io_pipe_phv_out_data_64; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_65 = init_io_pipe_phv_out_data_65; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_66 = init_io_pipe_phv_out_data_66; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_67 = init_io_pipe_phv_out_data_67; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_68 = init_io_pipe_phv_out_data_68; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_69 = init_io_pipe_phv_out_data_69; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_70 = init_io_pipe_phv_out_data_70; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_71 = init_io_pipe_phv_out_data_71; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_72 = init_io_pipe_phv_out_data_72; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_73 = init_io_pipe_phv_out_data_73; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_74 = init_io_pipe_phv_out_data_74; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_75 = init_io_pipe_phv_out_data_75; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_76 = init_io_pipe_phv_out_data_76; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_77 = init_io_pipe_phv_out_data_77; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_78 = init_io_pipe_phv_out_data_78; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_79 = init_io_pipe_phv_out_data_79; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_80 = init_io_pipe_phv_out_data_80; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_81 = init_io_pipe_phv_out_data_81; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_82 = init_io_pipe_phv_out_data_82; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_83 = init_io_pipe_phv_out_data_83; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_84 = init_io_pipe_phv_out_data_84; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_85 = init_io_pipe_phv_out_data_85; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_86 = init_io_pipe_phv_out_data_86; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_87 = init_io_pipe_phv_out_data_87; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_88 = init_io_pipe_phv_out_data_88; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_89 = init_io_pipe_phv_out_data_89; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_90 = init_io_pipe_phv_out_data_90; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_91 = init_io_pipe_phv_out_data_91; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_92 = init_io_pipe_phv_out_data_92; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_93 = init_io_pipe_phv_out_data_93; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_94 = init_io_pipe_phv_out_data_94; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_95 = init_io_pipe_phv_out_data_95; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_96 = init_io_pipe_phv_out_data_96; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_97 = init_io_pipe_phv_out_data_97; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_98 = init_io_pipe_phv_out_data_98; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_99 = init_io_pipe_phv_out_data_99; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_100 = init_io_pipe_phv_out_data_100; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_101 = init_io_pipe_phv_out_data_101; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_102 = init_io_pipe_phv_out_data_102; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_103 = init_io_pipe_phv_out_data_103; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_104 = init_io_pipe_phv_out_data_104; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_105 = init_io_pipe_phv_out_data_105; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_106 = init_io_pipe_phv_out_data_106; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_107 = init_io_pipe_phv_out_data_107; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_108 = init_io_pipe_phv_out_data_108; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_109 = init_io_pipe_phv_out_data_109; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_110 = init_io_pipe_phv_out_data_110; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_111 = init_io_pipe_phv_out_data_111; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_112 = init_io_pipe_phv_out_data_112; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_113 = init_io_pipe_phv_out_data_113; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_114 = init_io_pipe_phv_out_data_114; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_115 = init_io_pipe_phv_out_data_115; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_116 = init_io_pipe_phv_out_data_116; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_117 = init_io_pipe_phv_out_data_117; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_118 = init_io_pipe_phv_out_data_118; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_119 = init_io_pipe_phv_out_data_119; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_120 = init_io_pipe_phv_out_data_120; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_121 = init_io_pipe_phv_out_data_121; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_122 = init_io_pipe_phv_out_data_122; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_123 = init_io_pipe_phv_out_data_123; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_124 = init_io_pipe_phv_out_data_124; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_125 = init_io_pipe_phv_out_data_125; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_126 = init_io_pipe_phv_out_data_126; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_127 = init_io_pipe_phv_out_data_127; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_data_128 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_12_io_pipe_phv_in_data_129 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_12_io_pipe_phv_in_data_130 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_12_io_pipe_phv_in_data_131 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_12_io_pipe_phv_in_data_132 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_12_io_pipe_phv_in_data_133 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_12_io_pipe_phv_in_data_134 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_12_io_pipe_phv_in_data_135 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_12_io_pipe_phv_in_data_136 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_12_io_pipe_phv_in_data_137 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_12_io_pipe_phv_in_data_138 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_12_io_pipe_phv_in_data_139 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_12_io_pipe_phv_in_data_140 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_12_io_pipe_phv_in_data_141 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_12_io_pipe_phv_in_data_142 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_12_io_pipe_phv_in_data_143 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_12_io_pipe_phv_in_data_144 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_12_io_pipe_phv_in_data_145 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_12_io_pipe_phv_in_data_146 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_12_io_pipe_phv_in_data_147 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_12_io_pipe_phv_in_data_148 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_12_io_pipe_phv_in_data_149 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_12_io_pipe_phv_in_data_150 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_12_io_pipe_phv_in_data_151 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_12_io_pipe_phv_in_data_152 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_12_io_pipe_phv_in_data_153 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_12_io_pipe_phv_in_data_154 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_12_io_pipe_phv_in_data_155 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_12_io_pipe_phv_in_data_156 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_12_io_pipe_phv_in_data_157 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_12_io_pipe_phv_in_data_158 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_12_io_pipe_phv_in_data_159 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_12_io_pipe_phv_in_header_0 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_12_io_pipe_phv_in_header_1 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_12_io_pipe_phv_in_header_2 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_12_io_pipe_phv_in_header_3 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_12_io_pipe_phv_in_header_4 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_12_io_pipe_phv_in_header_5 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_12_io_pipe_phv_in_header_6 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_12_io_pipe_phv_in_header_7 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_12_io_pipe_phv_in_header_8 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_12_io_pipe_phv_in_header_9 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_12_io_pipe_phv_in_header_10 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_12_io_pipe_phv_in_header_11 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_12_io_pipe_phv_in_header_12 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_12_io_pipe_phv_in_header_13 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_12_io_pipe_phv_in_header_14 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_12_io_pipe_phv_in_header_15 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_12_io_pipe_phv_in_parse_current_state = 8'h0; // @[ipsa.scala 94:65]
  assign proc_12_io_pipe_phv_in_parse_current_offset = 8'h0; // @[ipsa.scala 94:65]
  assign proc_12_io_pipe_phv_in_parse_transition_field = 16'h0; // @[ipsa.scala 94:65]
  assign proc_12_io_pipe_phv_in_next_processor_id = 4'h0; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_next_config_id = 1'h0; // @[ipsa.scala 94:65]
  assign proc_12_io_pipe_phv_in_is_valid_processor = 1'h0; // @[ipsa.scala 94:65]
  assign proc_12_io_pipe_phv_in_valid = init_io_pipe_phv_out_valid; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_12_io_pipe_phv_in_last = init_io_pipe_phv_out_last; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_clock = clock;
  assign proc_13_io_pipe_phv_in_data_0 = init_io_pipe_phv_out_data_0; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_1 = init_io_pipe_phv_out_data_1; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_2 = init_io_pipe_phv_out_data_2; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_3 = init_io_pipe_phv_out_data_3; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_4 = init_io_pipe_phv_out_data_4; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_5 = init_io_pipe_phv_out_data_5; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_6 = init_io_pipe_phv_out_data_6; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_7 = init_io_pipe_phv_out_data_7; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_8 = init_io_pipe_phv_out_data_8; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_9 = init_io_pipe_phv_out_data_9; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_10 = init_io_pipe_phv_out_data_10; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_11 = init_io_pipe_phv_out_data_11; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_12 = init_io_pipe_phv_out_data_12; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_13 = init_io_pipe_phv_out_data_13; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_14 = init_io_pipe_phv_out_data_14; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_15 = init_io_pipe_phv_out_data_15; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_16 = init_io_pipe_phv_out_data_16; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_17 = init_io_pipe_phv_out_data_17; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_18 = init_io_pipe_phv_out_data_18; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_19 = init_io_pipe_phv_out_data_19; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_20 = init_io_pipe_phv_out_data_20; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_21 = init_io_pipe_phv_out_data_21; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_22 = init_io_pipe_phv_out_data_22; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_23 = init_io_pipe_phv_out_data_23; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_24 = init_io_pipe_phv_out_data_24; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_25 = init_io_pipe_phv_out_data_25; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_26 = init_io_pipe_phv_out_data_26; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_27 = init_io_pipe_phv_out_data_27; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_28 = init_io_pipe_phv_out_data_28; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_29 = init_io_pipe_phv_out_data_29; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_30 = init_io_pipe_phv_out_data_30; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_31 = init_io_pipe_phv_out_data_31; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_32 = init_io_pipe_phv_out_data_32; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_33 = init_io_pipe_phv_out_data_33; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_34 = init_io_pipe_phv_out_data_34; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_35 = init_io_pipe_phv_out_data_35; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_36 = init_io_pipe_phv_out_data_36; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_37 = init_io_pipe_phv_out_data_37; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_38 = init_io_pipe_phv_out_data_38; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_39 = init_io_pipe_phv_out_data_39; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_40 = init_io_pipe_phv_out_data_40; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_41 = init_io_pipe_phv_out_data_41; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_42 = init_io_pipe_phv_out_data_42; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_43 = init_io_pipe_phv_out_data_43; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_44 = init_io_pipe_phv_out_data_44; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_45 = init_io_pipe_phv_out_data_45; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_46 = init_io_pipe_phv_out_data_46; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_47 = init_io_pipe_phv_out_data_47; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_48 = init_io_pipe_phv_out_data_48; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_49 = init_io_pipe_phv_out_data_49; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_50 = init_io_pipe_phv_out_data_50; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_51 = init_io_pipe_phv_out_data_51; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_52 = init_io_pipe_phv_out_data_52; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_53 = init_io_pipe_phv_out_data_53; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_54 = init_io_pipe_phv_out_data_54; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_55 = init_io_pipe_phv_out_data_55; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_56 = init_io_pipe_phv_out_data_56; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_57 = init_io_pipe_phv_out_data_57; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_58 = init_io_pipe_phv_out_data_58; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_59 = init_io_pipe_phv_out_data_59; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_60 = init_io_pipe_phv_out_data_60; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_61 = init_io_pipe_phv_out_data_61; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_62 = init_io_pipe_phv_out_data_62; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_63 = init_io_pipe_phv_out_data_63; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_64 = init_io_pipe_phv_out_data_64; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_65 = init_io_pipe_phv_out_data_65; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_66 = init_io_pipe_phv_out_data_66; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_67 = init_io_pipe_phv_out_data_67; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_68 = init_io_pipe_phv_out_data_68; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_69 = init_io_pipe_phv_out_data_69; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_70 = init_io_pipe_phv_out_data_70; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_71 = init_io_pipe_phv_out_data_71; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_72 = init_io_pipe_phv_out_data_72; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_73 = init_io_pipe_phv_out_data_73; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_74 = init_io_pipe_phv_out_data_74; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_75 = init_io_pipe_phv_out_data_75; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_76 = init_io_pipe_phv_out_data_76; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_77 = init_io_pipe_phv_out_data_77; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_78 = init_io_pipe_phv_out_data_78; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_79 = init_io_pipe_phv_out_data_79; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_80 = init_io_pipe_phv_out_data_80; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_81 = init_io_pipe_phv_out_data_81; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_82 = init_io_pipe_phv_out_data_82; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_83 = init_io_pipe_phv_out_data_83; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_84 = init_io_pipe_phv_out_data_84; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_85 = init_io_pipe_phv_out_data_85; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_86 = init_io_pipe_phv_out_data_86; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_87 = init_io_pipe_phv_out_data_87; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_88 = init_io_pipe_phv_out_data_88; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_89 = init_io_pipe_phv_out_data_89; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_90 = init_io_pipe_phv_out_data_90; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_91 = init_io_pipe_phv_out_data_91; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_92 = init_io_pipe_phv_out_data_92; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_93 = init_io_pipe_phv_out_data_93; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_94 = init_io_pipe_phv_out_data_94; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_95 = init_io_pipe_phv_out_data_95; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_96 = init_io_pipe_phv_out_data_96; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_97 = init_io_pipe_phv_out_data_97; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_98 = init_io_pipe_phv_out_data_98; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_99 = init_io_pipe_phv_out_data_99; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_100 = init_io_pipe_phv_out_data_100; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_101 = init_io_pipe_phv_out_data_101; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_102 = init_io_pipe_phv_out_data_102; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_103 = init_io_pipe_phv_out_data_103; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_104 = init_io_pipe_phv_out_data_104; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_105 = init_io_pipe_phv_out_data_105; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_106 = init_io_pipe_phv_out_data_106; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_107 = init_io_pipe_phv_out_data_107; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_108 = init_io_pipe_phv_out_data_108; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_109 = init_io_pipe_phv_out_data_109; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_110 = init_io_pipe_phv_out_data_110; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_111 = init_io_pipe_phv_out_data_111; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_112 = init_io_pipe_phv_out_data_112; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_113 = init_io_pipe_phv_out_data_113; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_114 = init_io_pipe_phv_out_data_114; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_115 = init_io_pipe_phv_out_data_115; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_116 = init_io_pipe_phv_out_data_116; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_117 = init_io_pipe_phv_out_data_117; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_118 = init_io_pipe_phv_out_data_118; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_119 = init_io_pipe_phv_out_data_119; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_120 = init_io_pipe_phv_out_data_120; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_121 = init_io_pipe_phv_out_data_121; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_122 = init_io_pipe_phv_out_data_122; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_123 = init_io_pipe_phv_out_data_123; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_124 = init_io_pipe_phv_out_data_124; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_125 = init_io_pipe_phv_out_data_125; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_126 = init_io_pipe_phv_out_data_126; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_127 = init_io_pipe_phv_out_data_127; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_data_128 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_13_io_pipe_phv_in_data_129 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_13_io_pipe_phv_in_data_130 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_13_io_pipe_phv_in_data_131 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_13_io_pipe_phv_in_data_132 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_13_io_pipe_phv_in_data_133 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_13_io_pipe_phv_in_data_134 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_13_io_pipe_phv_in_data_135 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_13_io_pipe_phv_in_data_136 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_13_io_pipe_phv_in_data_137 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_13_io_pipe_phv_in_data_138 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_13_io_pipe_phv_in_data_139 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_13_io_pipe_phv_in_data_140 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_13_io_pipe_phv_in_data_141 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_13_io_pipe_phv_in_data_142 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_13_io_pipe_phv_in_data_143 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_13_io_pipe_phv_in_data_144 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_13_io_pipe_phv_in_data_145 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_13_io_pipe_phv_in_data_146 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_13_io_pipe_phv_in_data_147 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_13_io_pipe_phv_in_data_148 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_13_io_pipe_phv_in_data_149 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_13_io_pipe_phv_in_data_150 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_13_io_pipe_phv_in_data_151 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_13_io_pipe_phv_in_data_152 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_13_io_pipe_phv_in_data_153 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_13_io_pipe_phv_in_data_154 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_13_io_pipe_phv_in_data_155 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_13_io_pipe_phv_in_data_156 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_13_io_pipe_phv_in_data_157 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_13_io_pipe_phv_in_data_158 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_13_io_pipe_phv_in_data_159 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_13_io_pipe_phv_in_header_0 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_13_io_pipe_phv_in_header_1 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_13_io_pipe_phv_in_header_2 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_13_io_pipe_phv_in_header_3 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_13_io_pipe_phv_in_header_4 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_13_io_pipe_phv_in_header_5 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_13_io_pipe_phv_in_header_6 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_13_io_pipe_phv_in_header_7 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_13_io_pipe_phv_in_header_8 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_13_io_pipe_phv_in_header_9 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_13_io_pipe_phv_in_header_10 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_13_io_pipe_phv_in_header_11 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_13_io_pipe_phv_in_header_12 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_13_io_pipe_phv_in_header_13 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_13_io_pipe_phv_in_header_14 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_13_io_pipe_phv_in_header_15 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_13_io_pipe_phv_in_parse_current_state = 8'h0; // @[ipsa.scala 94:65]
  assign proc_13_io_pipe_phv_in_parse_current_offset = 8'h0; // @[ipsa.scala 94:65]
  assign proc_13_io_pipe_phv_in_parse_transition_field = 16'h0; // @[ipsa.scala 94:65]
  assign proc_13_io_pipe_phv_in_next_processor_id = 4'h0; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_next_config_id = 1'h0; // @[ipsa.scala 94:65]
  assign proc_13_io_pipe_phv_in_is_valid_processor = 1'h0; // @[ipsa.scala 94:65]
  assign proc_13_io_pipe_phv_in_valid = init_io_pipe_phv_out_valid; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_13_io_pipe_phv_in_last = init_io_pipe_phv_out_last; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_clock = clock;
  assign proc_14_io_pipe_phv_in_data_0 = init_io_pipe_phv_out_data_0; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_1 = init_io_pipe_phv_out_data_1; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_2 = init_io_pipe_phv_out_data_2; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_3 = init_io_pipe_phv_out_data_3; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_4 = init_io_pipe_phv_out_data_4; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_5 = init_io_pipe_phv_out_data_5; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_6 = init_io_pipe_phv_out_data_6; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_7 = init_io_pipe_phv_out_data_7; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_8 = init_io_pipe_phv_out_data_8; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_9 = init_io_pipe_phv_out_data_9; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_10 = init_io_pipe_phv_out_data_10; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_11 = init_io_pipe_phv_out_data_11; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_12 = init_io_pipe_phv_out_data_12; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_13 = init_io_pipe_phv_out_data_13; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_14 = init_io_pipe_phv_out_data_14; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_15 = init_io_pipe_phv_out_data_15; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_16 = init_io_pipe_phv_out_data_16; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_17 = init_io_pipe_phv_out_data_17; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_18 = init_io_pipe_phv_out_data_18; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_19 = init_io_pipe_phv_out_data_19; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_20 = init_io_pipe_phv_out_data_20; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_21 = init_io_pipe_phv_out_data_21; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_22 = init_io_pipe_phv_out_data_22; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_23 = init_io_pipe_phv_out_data_23; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_24 = init_io_pipe_phv_out_data_24; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_25 = init_io_pipe_phv_out_data_25; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_26 = init_io_pipe_phv_out_data_26; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_27 = init_io_pipe_phv_out_data_27; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_28 = init_io_pipe_phv_out_data_28; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_29 = init_io_pipe_phv_out_data_29; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_30 = init_io_pipe_phv_out_data_30; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_31 = init_io_pipe_phv_out_data_31; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_32 = init_io_pipe_phv_out_data_32; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_33 = init_io_pipe_phv_out_data_33; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_34 = init_io_pipe_phv_out_data_34; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_35 = init_io_pipe_phv_out_data_35; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_36 = init_io_pipe_phv_out_data_36; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_37 = init_io_pipe_phv_out_data_37; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_38 = init_io_pipe_phv_out_data_38; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_39 = init_io_pipe_phv_out_data_39; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_40 = init_io_pipe_phv_out_data_40; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_41 = init_io_pipe_phv_out_data_41; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_42 = init_io_pipe_phv_out_data_42; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_43 = init_io_pipe_phv_out_data_43; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_44 = init_io_pipe_phv_out_data_44; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_45 = init_io_pipe_phv_out_data_45; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_46 = init_io_pipe_phv_out_data_46; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_47 = init_io_pipe_phv_out_data_47; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_48 = init_io_pipe_phv_out_data_48; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_49 = init_io_pipe_phv_out_data_49; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_50 = init_io_pipe_phv_out_data_50; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_51 = init_io_pipe_phv_out_data_51; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_52 = init_io_pipe_phv_out_data_52; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_53 = init_io_pipe_phv_out_data_53; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_54 = init_io_pipe_phv_out_data_54; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_55 = init_io_pipe_phv_out_data_55; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_56 = init_io_pipe_phv_out_data_56; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_57 = init_io_pipe_phv_out_data_57; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_58 = init_io_pipe_phv_out_data_58; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_59 = init_io_pipe_phv_out_data_59; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_60 = init_io_pipe_phv_out_data_60; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_61 = init_io_pipe_phv_out_data_61; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_62 = init_io_pipe_phv_out_data_62; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_63 = init_io_pipe_phv_out_data_63; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_64 = init_io_pipe_phv_out_data_64; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_65 = init_io_pipe_phv_out_data_65; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_66 = init_io_pipe_phv_out_data_66; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_67 = init_io_pipe_phv_out_data_67; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_68 = init_io_pipe_phv_out_data_68; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_69 = init_io_pipe_phv_out_data_69; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_70 = init_io_pipe_phv_out_data_70; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_71 = init_io_pipe_phv_out_data_71; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_72 = init_io_pipe_phv_out_data_72; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_73 = init_io_pipe_phv_out_data_73; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_74 = init_io_pipe_phv_out_data_74; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_75 = init_io_pipe_phv_out_data_75; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_76 = init_io_pipe_phv_out_data_76; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_77 = init_io_pipe_phv_out_data_77; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_78 = init_io_pipe_phv_out_data_78; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_79 = init_io_pipe_phv_out_data_79; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_80 = init_io_pipe_phv_out_data_80; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_81 = init_io_pipe_phv_out_data_81; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_82 = init_io_pipe_phv_out_data_82; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_83 = init_io_pipe_phv_out_data_83; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_84 = init_io_pipe_phv_out_data_84; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_85 = init_io_pipe_phv_out_data_85; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_86 = init_io_pipe_phv_out_data_86; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_87 = init_io_pipe_phv_out_data_87; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_88 = init_io_pipe_phv_out_data_88; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_89 = init_io_pipe_phv_out_data_89; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_90 = init_io_pipe_phv_out_data_90; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_91 = init_io_pipe_phv_out_data_91; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_92 = init_io_pipe_phv_out_data_92; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_93 = init_io_pipe_phv_out_data_93; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_94 = init_io_pipe_phv_out_data_94; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_95 = init_io_pipe_phv_out_data_95; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_96 = init_io_pipe_phv_out_data_96; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_97 = init_io_pipe_phv_out_data_97; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_98 = init_io_pipe_phv_out_data_98; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_99 = init_io_pipe_phv_out_data_99; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_100 = init_io_pipe_phv_out_data_100; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_101 = init_io_pipe_phv_out_data_101; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_102 = init_io_pipe_phv_out_data_102; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_103 = init_io_pipe_phv_out_data_103; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_104 = init_io_pipe_phv_out_data_104; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_105 = init_io_pipe_phv_out_data_105; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_106 = init_io_pipe_phv_out_data_106; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_107 = init_io_pipe_phv_out_data_107; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_108 = init_io_pipe_phv_out_data_108; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_109 = init_io_pipe_phv_out_data_109; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_110 = init_io_pipe_phv_out_data_110; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_111 = init_io_pipe_phv_out_data_111; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_112 = init_io_pipe_phv_out_data_112; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_113 = init_io_pipe_phv_out_data_113; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_114 = init_io_pipe_phv_out_data_114; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_115 = init_io_pipe_phv_out_data_115; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_116 = init_io_pipe_phv_out_data_116; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_117 = init_io_pipe_phv_out_data_117; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_118 = init_io_pipe_phv_out_data_118; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_119 = init_io_pipe_phv_out_data_119; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_120 = init_io_pipe_phv_out_data_120; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_121 = init_io_pipe_phv_out_data_121; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_122 = init_io_pipe_phv_out_data_122; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_123 = init_io_pipe_phv_out_data_123; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_124 = init_io_pipe_phv_out_data_124; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_125 = init_io_pipe_phv_out_data_125; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_126 = init_io_pipe_phv_out_data_126; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_127 = init_io_pipe_phv_out_data_127; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_data_128 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_14_io_pipe_phv_in_data_129 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_14_io_pipe_phv_in_data_130 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_14_io_pipe_phv_in_data_131 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_14_io_pipe_phv_in_data_132 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_14_io_pipe_phv_in_data_133 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_14_io_pipe_phv_in_data_134 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_14_io_pipe_phv_in_data_135 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_14_io_pipe_phv_in_data_136 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_14_io_pipe_phv_in_data_137 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_14_io_pipe_phv_in_data_138 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_14_io_pipe_phv_in_data_139 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_14_io_pipe_phv_in_data_140 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_14_io_pipe_phv_in_data_141 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_14_io_pipe_phv_in_data_142 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_14_io_pipe_phv_in_data_143 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_14_io_pipe_phv_in_data_144 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_14_io_pipe_phv_in_data_145 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_14_io_pipe_phv_in_data_146 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_14_io_pipe_phv_in_data_147 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_14_io_pipe_phv_in_data_148 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_14_io_pipe_phv_in_data_149 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_14_io_pipe_phv_in_data_150 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_14_io_pipe_phv_in_data_151 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_14_io_pipe_phv_in_data_152 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_14_io_pipe_phv_in_data_153 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_14_io_pipe_phv_in_data_154 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_14_io_pipe_phv_in_data_155 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_14_io_pipe_phv_in_data_156 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_14_io_pipe_phv_in_data_157 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_14_io_pipe_phv_in_data_158 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_14_io_pipe_phv_in_data_159 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_14_io_pipe_phv_in_header_0 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_14_io_pipe_phv_in_header_1 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_14_io_pipe_phv_in_header_2 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_14_io_pipe_phv_in_header_3 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_14_io_pipe_phv_in_header_4 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_14_io_pipe_phv_in_header_5 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_14_io_pipe_phv_in_header_6 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_14_io_pipe_phv_in_header_7 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_14_io_pipe_phv_in_header_8 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_14_io_pipe_phv_in_header_9 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_14_io_pipe_phv_in_header_10 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_14_io_pipe_phv_in_header_11 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_14_io_pipe_phv_in_header_12 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_14_io_pipe_phv_in_header_13 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_14_io_pipe_phv_in_header_14 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_14_io_pipe_phv_in_header_15 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_14_io_pipe_phv_in_parse_current_state = 8'h0; // @[ipsa.scala 94:65]
  assign proc_14_io_pipe_phv_in_parse_current_offset = 8'h0; // @[ipsa.scala 94:65]
  assign proc_14_io_pipe_phv_in_parse_transition_field = 16'h0; // @[ipsa.scala 94:65]
  assign proc_14_io_pipe_phv_in_next_processor_id = 4'h0; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_next_config_id = 1'h0; // @[ipsa.scala 94:65]
  assign proc_14_io_pipe_phv_in_is_valid_processor = 1'h0; // @[ipsa.scala 94:65]
  assign proc_14_io_pipe_phv_in_valid = init_io_pipe_phv_out_valid; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_14_io_pipe_phv_in_last = init_io_pipe_phv_out_last; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_clock = clock;
  assign proc_15_io_pipe_phv_in_data_0 = init_io_pipe_phv_out_data_0; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_1 = init_io_pipe_phv_out_data_1; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_2 = init_io_pipe_phv_out_data_2; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_3 = init_io_pipe_phv_out_data_3; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_4 = init_io_pipe_phv_out_data_4; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_5 = init_io_pipe_phv_out_data_5; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_6 = init_io_pipe_phv_out_data_6; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_7 = init_io_pipe_phv_out_data_7; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_8 = init_io_pipe_phv_out_data_8; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_9 = init_io_pipe_phv_out_data_9; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_10 = init_io_pipe_phv_out_data_10; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_11 = init_io_pipe_phv_out_data_11; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_12 = init_io_pipe_phv_out_data_12; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_13 = init_io_pipe_phv_out_data_13; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_14 = init_io_pipe_phv_out_data_14; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_15 = init_io_pipe_phv_out_data_15; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_16 = init_io_pipe_phv_out_data_16; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_17 = init_io_pipe_phv_out_data_17; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_18 = init_io_pipe_phv_out_data_18; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_19 = init_io_pipe_phv_out_data_19; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_20 = init_io_pipe_phv_out_data_20; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_21 = init_io_pipe_phv_out_data_21; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_22 = init_io_pipe_phv_out_data_22; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_23 = init_io_pipe_phv_out_data_23; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_24 = init_io_pipe_phv_out_data_24; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_25 = init_io_pipe_phv_out_data_25; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_26 = init_io_pipe_phv_out_data_26; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_27 = init_io_pipe_phv_out_data_27; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_28 = init_io_pipe_phv_out_data_28; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_29 = init_io_pipe_phv_out_data_29; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_30 = init_io_pipe_phv_out_data_30; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_31 = init_io_pipe_phv_out_data_31; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_32 = init_io_pipe_phv_out_data_32; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_33 = init_io_pipe_phv_out_data_33; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_34 = init_io_pipe_phv_out_data_34; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_35 = init_io_pipe_phv_out_data_35; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_36 = init_io_pipe_phv_out_data_36; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_37 = init_io_pipe_phv_out_data_37; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_38 = init_io_pipe_phv_out_data_38; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_39 = init_io_pipe_phv_out_data_39; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_40 = init_io_pipe_phv_out_data_40; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_41 = init_io_pipe_phv_out_data_41; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_42 = init_io_pipe_phv_out_data_42; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_43 = init_io_pipe_phv_out_data_43; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_44 = init_io_pipe_phv_out_data_44; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_45 = init_io_pipe_phv_out_data_45; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_46 = init_io_pipe_phv_out_data_46; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_47 = init_io_pipe_phv_out_data_47; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_48 = init_io_pipe_phv_out_data_48; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_49 = init_io_pipe_phv_out_data_49; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_50 = init_io_pipe_phv_out_data_50; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_51 = init_io_pipe_phv_out_data_51; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_52 = init_io_pipe_phv_out_data_52; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_53 = init_io_pipe_phv_out_data_53; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_54 = init_io_pipe_phv_out_data_54; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_55 = init_io_pipe_phv_out_data_55; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_56 = init_io_pipe_phv_out_data_56; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_57 = init_io_pipe_phv_out_data_57; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_58 = init_io_pipe_phv_out_data_58; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_59 = init_io_pipe_phv_out_data_59; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_60 = init_io_pipe_phv_out_data_60; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_61 = init_io_pipe_phv_out_data_61; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_62 = init_io_pipe_phv_out_data_62; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_63 = init_io_pipe_phv_out_data_63; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_64 = init_io_pipe_phv_out_data_64; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_65 = init_io_pipe_phv_out_data_65; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_66 = init_io_pipe_phv_out_data_66; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_67 = init_io_pipe_phv_out_data_67; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_68 = init_io_pipe_phv_out_data_68; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_69 = init_io_pipe_phv_out_data_69; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_70 = init_io_pipe_phv_out_data_70; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_71 = init_io_pipe_phv_out_data_71; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_72 = init_io_pipe_phv_out_data_72; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_73 = init_io_pipe_phv_out_data_73; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_74 = init_io_pipe_phv_out_data_74; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_75 = init_io_pipe_phv_out_data_75; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_76 = init_io_pipe_phv_out_data_76; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_77 = init_io_pipe_phv_out_data_77; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_78 = init_io_pipe_phv_out_data_78; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_79 = init_io_pipe_phv_out_data_79; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_80 = init_io_pipe_phv_out_data_80; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_81 = init_io_pipe_phv_out_data_81; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_82 = init_io_pipe_phv_out_data_82; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_83 = init_io_pipe_phv_out_data_83; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_84 = init_io_pipe_phv_out_data_84; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_85 = init_io_pipe_phv_out_data_85; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_86 = init_io_pipe_phv_out_data_86; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_87 = init_io_pipe_phv_out_data_87; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_88 = init_io_pipe_phv_out_data_88; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_89 = init_io_pipe_phv_out_data_89; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_90 = init_io_pipe_phv_out_data_90; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_91 = init_io_pipe_phv_out_data_91; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_92 = init_io_pipe_phv_out_data_92; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_93 = init_io_pipe_phv_out_data_93; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_94 = init_io_pipe_phv_out_data_94; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_95 = init_io_pipe_phv_out_data_95; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_96 = init_io_pipe_phv_out_data_96; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_97 = init_io_pipe_phv_out_data_97; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_98 = init_io_pipe_phv_out_data_98; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_99 = init_io_pipe_phv_out_data_99; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_100 = init_io_pipe_phv_out_data_100; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_101 = init_io_pipe_phv_out_data_101; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_102 = init_io_pipe_phv_out_data_102; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_103 = init_io_pipe_phv_out_data_103; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_104 = init_io_pipe_phv_out_data_104; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_105 = init_io_pipe_phv_out_data_105; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_106 = init_io_pipe_phv_out_data_106; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_107 = init_io_pipe_phv_out_data_107; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_108 = init_io_pipe_phv_out_data_108; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_109 = init_io_pipe_phv_out_data_109; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_110 = init_io_pipe_phv_out_data_110; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_111 = init_io_pipe_phv_out_data_111; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_112 = init_io_pipe_phv_out_data_112; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_113 = init_io_pipe_phv_out_data_113; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_114 = init_io_pipe_phv_out_data_114; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_115 = init_io_pipe_phv_out_data_115; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_116 = init_io_pipe_phv_out_data_116; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_117 = init_io_pipe_phv_out_data_117; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_118 = init_io_pipe_phv_out_data_118; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_119 = init_io_pipe_phv_out_data_119; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_120 = init_io_pipe_phv_out_data_120; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_121 = init_io_pipe_phv_out_data_121; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_122 = init_io_pipe_phv_out_data_122; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_123 = init_io_pipe_phv_out_data_123; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_124 = init_io_pipe_phv_out_data_124; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_125 = init_io_pipe_phv_out_data_125; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_126 = init_io_pipe_phv_out_data_126; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_127 = init_io_pipe_phv_out_data_127; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_data_128 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_15_io_pipe_phv_in_data_129 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_15_io_pipe_phv_in_data_130 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_15_io_pipe_phv_in_data_131 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_15_io_pipe_phv_in_data_132 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_15_io_pipe_phv_in_data_133 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_15_io_pipe_phv_in_data_134 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_15_io_pipe_phv_in_data_135 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_15_io_pipe_phv_in_data_136 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_15_io_pipe_phv_in_data_137 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_15_io_pipe_phv_in_data_138 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_15_io_pipe_phv_in_data_139 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_15_io_pipe_phv_in_data_140 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_15_io_pipe_phv_in_data_141 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_15_io_pipe_phv_in_data_142 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_15_io_pipe_phv_in_data_143 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_15_io_pipe_phv_in_data_144 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_15_io_pipe_phv_in_data_145 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_15_io_pipe_phv_in_data_146 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_15_io_pipe_phv_in_data_147 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_15_io_pipe_phv_in_data_148 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_15_io_pipe_phv_in_data_149 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_15_io_pipe_phv_in_data_150 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_15_io_pipe_phv_in_data_151 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_15_io_pipe_phv_in_data_152 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_15_io_pipe_phv_in_data_153 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_15_io_pipe_phv_in_data_154 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_15_io_pipe_phv_in_data_155 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_15_io_pipe_phv_in_data_156 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_15_io_pipe_phv_in_data_157 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_15_io_pipe_phv_in_data_158 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_15_io_pipe_phv_in_data_159 = 8'h0; // @[ipsa.scala 94:65]
  assign proc_15_io_pipe_phv_in_header_0 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_15_io_pipe_phv_in_header_1 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_15_io_pipe_phv_in_header_2 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_15_io_pipe_phv_in_header_3 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_15_io_pipe_phv_in_header_4 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_15_io_pipe_phv_in_header_5 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_15_io_pipe_phv_in_header_6 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_15_io_pipe_phv_in_header_7 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_15_io_pipe_phv_in_header_8 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_15_io_pipe_phv_in_header_9 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_15_io_pipe_phv_in_header_10 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_15_io_pipe_phv_in_header_11 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_15_io_pipe_phv_in_header_12 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_15_io_pipe_phv_in_header_13 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_15_io_pipe_phv_in_header_14 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_15_io_pipe_phv_in_header_15 = 16'h0; // @[ipsa.scala 94:65]
  assign proc_15_io_pipe_phv_in_parse_current_state = 8'h0; // @[ipsa.scala 94:65]
  assign proc_15_io_pipe_phv_in_parse_current_offset = 8'h0; // @[ipsa.scala 94:65]
  assign proc_15_io_pipe_phv_in_parse_transition_field = 16'h0; // @[ipsa.scala 94:65]
  assign proc_15_io_pipe_phv_in_next_processor_id = 4'h0; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_next_config_id = 1'h0; // @[ipsa.scala 94:65]
  assign proc_15_io_pipe_phv_in_is_valid_processor = 1'h0; // @[ipsa.scala 94:65]
  assign proc_15_io_pipe_phv_in_valid = init_io_pipe_phv_out_valid; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign proc_15_io_pipe_phv_in_last = init_io_pipe_phv_out_last; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  assign sram_cluster_0_clock = clock;
  assign sram_cluster_1_clock = clock;
  assign sram_cluster_2_clock = clock;
  assign sram_cluster_3_clock = clock;
  assign sram_cluster_4_clock = clock;
  assign sram_cluster_5_clock = clock;
  assign sram_cluster_6_clock = clock;
  assign sram_cluster_7_clock = clock;
  assign init_clock = clock;
  assign init_io_pipe_phv_in_data_0 = io_pipe_phv_in_data_0; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_1 = io_pipe_phv_in_data_1; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_2 = io_pipe_phv_in_data_2; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_3 = io_pipe_phv_in_data_3; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_4 = io_pipe_phv_in_data_4; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_5 = io_pipe_phv_in_data_5; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_6 = io_pipe_phv_in_data_6; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_7 = io_pipe_phv_in_data_7; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_8 = io_pipe_phv_in_data_8; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_9 = io_pipe_phv_in_data_9; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_10 = io_pipe_phv_in_data_10; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_11 = io_pipe_phv_in_data_11; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_12 = io_pipe_phv_in_data_12; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_13 = io_pipe_phv_in_data_13; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_14 = io_pipe_phv_in_data_14; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_15 = io_pipe_phv_in_data_15; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_16 = io_pipe_phv_in_data_16; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_17 = io_pipe_phv_in_data_17; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_18 = io_pipe_phv_in_data_18; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_19 = io_pipe_phv_in_data_19; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_20 = io_pipe_phv_in_data_20; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_21 = io_pipe_phv_in_data_21; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_22 = io_pipe_phv_in_data_22; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_23 = io_pipe_phv_in_data_23; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_24 = io_pipe_phv_in_data_24; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_25 = io_pipe_phv_in_data_25; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_26 = io_pipe_phv_in_data_26; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_27 = io_pipe_phv_in_data_27; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_28 = io_pipe_phv_in_data_28; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_29 = io_pipe_phv_in_data_29; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_30 = io_pipe_phv_in_data_30; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_31 = io_pipe_phv_in_data_31; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_32 = io_pipe_phv_in_data_32; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_33 = io_pipe_phv_in_data_33; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_34 = io_pipe_phv_in_data_34; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_35 = io_pipe_phv_in_data_35; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_36 = io_pipe_phv_in_data_36; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_37 = io_pipe_phv_in_data_37; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_38 = io_pipe_phv_in_data_38; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_39 = io_pipe_phv_in_data_39; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_40 = io_pipe_phv_in_data_40; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_41 = io_pipe_phv_in_data_41; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_42 = io_pipe_phv_in_data_42; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_43 = io_pipe_phv_in_data_43; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_44 = io_pipe_phv_in_data_44; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_45 = io_pipe_phv_in_data_45; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_46 = io_pipe_phv_in_data_46; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_47 = io_pipe_phv_in_data_47; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_48 = io_pipe_phv_in_data_48; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_49 = io_pipe_phv_in_data_49; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_50 = io_pipe_phv_in_data_50; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_51 = io_pipe_phv_in_data_51; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_52 = io_pipe_phv_in_data_52; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_53 = io_pipe_phv_in_data_53; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_54 = io_pipe_phv_in_data_54; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_55 = io_pipe_phv_in_data_55; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_56 = io_pipe_phv_in_data_56; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_57 = io_pipe_phv_in_data_57; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_58 = io_pipe_phv_in_data_58; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_59 = io_pipe_phv_in_data_59; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_60 = io_pipe_phv_in_data_60; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_61 = io_pipe_phv_in_data_61; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_62 = io_pipe_phv_in_data_62; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_63 = io_pipe_phv_in_data_63; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_64 = io_pipe_phv_in_data_64; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_65 = io_pipe_phv_in_data_65; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_66 = io_pipe_phv_in_data_66; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_67 = io_pipe_phv_in_data_67; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_68 = io_pipe_phv_in_data_68; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_69 = io_pipe_phv_in_data_69; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_70 = io_pipe_phv_in_data_70; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_71 = io_pipe_phv_in_data_71; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_72 = io_pipe_phv_in_data_72; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_73 = io_pipe_phv_in_data_73; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_74 = io_pipe_phv_in_data_74; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_75 = io_pipe_phv_in_data_75; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_76 = io_pipe_phv_in_data_76; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_77 = io_pipe_phv_in_data_77; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_78 = io_pipe_phv_in_data_78; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_79 = io_pipe_phv_in_data_79; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_80 = io_pipe_phv_in_data_80; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_81 = io_pipe_phv_in_data_81; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_82 = io_pipe_phv_in_data_82; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_83 = io_pipe_phv_in_data_83; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_84 = io_pipe_phv_in_data_84; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_85 = io_pipe_phv_in_data_85; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_86 = io_pipe_phv_in_data_86; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_87 = io_pipe_phv_in_data_87; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_88 = io_pipe_phv_in_data_88; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_89 = io_pipe_phv_in_data_89; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_90 = io_pipe_phv_in_data_90; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_91 = io_pipe_phv_in_data_91; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_92 = io_pipe_phv_in_data_92; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_93 = io_pipe_phv_in_data_93; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_94 = io_pipe_phv_in_data_94; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_95 = io_pipe_phv_in_data_95; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_96 = io_pipe_phv_in_data_96; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_97 = io_pipe_phv_in_data_97; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_98 = io_pipe_phv_in_data_98; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_99 = io_pipe_phv_in_data_99; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_100 = io_pipe_phv_in_data_100; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_101 = io_pipe_phv_in_data_101; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_102 = io_pipe_phv_in_data_102; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_103 = io_pipe_phv_in_data_103; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_104 = io_pipe_phv_in_data_104; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_105 = io_pipe_phv_in_data_105; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_106 = io_pipe_phv_in_data_106; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_107 = io_pipe_phv_in_data_107; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_108 = io_pipe_phv_in_data_108; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_109 = io_pipe_phv_in_data_109; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_110 = io_pipe_phv_in_data_110; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_111 = io_pipe_phv_in_data_111; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_112 = io_pipe_phv_in_data_112; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_113 = io_pipe_phv_in_data_113; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_114 = io_pipe_phv_in_data_114; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_115 = io_pipe_phv_in_data_115; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_116 = io_pipe_phv_in_data_116; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_117 = io_pipe_phv_in_data_117; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_118 = io_pipe_phv_in_data_118; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_119 = io_pipe_phv_in_data_119; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_120 = io_pipe_phv_in_data_120; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_121 = io_pipe_phv_in_data_121; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_122 = io_pipe_phv_in_data_122; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_123 = io_pipe_phv_in_data_123; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_124 = io_pipe_phv_in_data_124; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_125 = io_pipe_phv_in_data_125; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_126 = io_pipe_phv_in_data_126; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_127 = io_pipe_phv_in_data_127; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_valid = io_pipe_phv_in_valid; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_last = io_pipe_phv_in_last; // @[ipsa.scala 75:25]
  assign trans_0_clock = clock;
  assign trans_0_io_pipe_phv_in_data_0 = proc_0_io_pipe_phv_out_data_0; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_1 = proc_0_io_pipe_phv_out_data_1; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_2 = proc_0_io_pipe_phv_out_data_2; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_3 = proc_0_io_pipe_phv_out_data_3; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_4 = proc_0_io_pipe_phv_out_data_4; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_5 = proc_0_io_pipe_phv_out_data_5; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_6 = proc_0_io_pipe_phv_out_data_6; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_7 = proc_0_io_pipe_phv_out_data_7; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_8 = proc_0_io_pipe_phv_out_data_8; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_9 = proc_0_io_pipe_phv_out_data_9; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_10 = proc_0_io_pipe_phv_out_data_10; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_11 = proc_0_io_pipe_phv_out_data_11; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_12 = proc_0_io_pipe_phv_out_data_12; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_13 = proc_0_io_pipe_phv_out_data_13; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_14 = proc_0_io_pipe_phv_out_data_14; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_15 = proc_0_io_pipe_phv_out_data_15; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_16 = proc_0_io_pipe_phv_out_data_16; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_17 = proc_0_io_pipe_phv_out_data_17; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_18 = proc_0_io_pipe_phv_out_data_18; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_19 = proc_0_io_pipe_phv_out_data_19; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_20 = proc_0_io_pipe_phv_out_data_20; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_21 = proc_0_io_pipe_phv_out_data_21; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_22 = proc_0_io_pipe_phv_out_data_22; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_23 = proc_0_io_pipe_phv_out_data_23; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_24 = proc_0_io_pipe_phv_out_data_24; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_25 = proc_0_io_pipe_phv_out_data_25; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_26 = proc_0_io_pipe_phv_out_data_26; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_27 = proc_0_io_pipe_phv_out_data_27; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_28 = proc_0_io_pipe_phv_out_data_28; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_29 = proc_0_io_pipe_phv_out_data_29; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_30 = proc_0_io_pipe_phv_out_data_30; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_31 = proc_0_io_pipe_phv_out_data_31; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_32 = proc_0_io_pipe_phv_out_data_32; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_33 = proc_0_io_pipe_phv_out_data_33; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_34 = proc_0_io_pipe_phv_out_data_34; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_35 = proc_0_io_pipe_phv_out_data_35; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_36 = proc_0_io_pipe_phv_out_data_36; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_37 = proc_0_io_pipe_phv_out_data_37; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_38 = proc_0_io_pipe_phv_out_data_38; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_39 = proc_0_io_pipe_phv_out_data_39; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_40 = proc_0_io_pipe_phv_out_data_40; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_41 = proc_0_io_pipe_phv_out_data_41; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_42 = proc_0_io_pipe_phv_out_data_42; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_43 = proc_0_io_pipe_phv_out_data_43; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_44 = proc_0_io_pipe_phv_out_data_44; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_45 = proc_0_io_pipe_phv_out_data_45; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_46 = proc_0_io_pipe_phv_out_data_46; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_47 = proc_0_io_pipe_phv_out_data_47; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_48 = proc_0_io_pipe_phv_out_data_48; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_49 = proc_0_io_pipe_phv_out_data_49; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_50 = proc_0_io_pipe_phv_out_data_50; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_51 = proc_0_io_pipe_phv_out_data_51; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_52 = proc_0_io_pipe_phv_out_data_52; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_53 = proc_0_io_pipe_phv_out_data_53; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_54 = proc_0_io_pipe_phv_out_data_54; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_55 = proc_0_io_pipe_phv_out_data_55; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_56 = proc_0_io_pipe_phv_out_data_56; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_57 = proc_0_io_pipe_phv_out_data_57; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_58 = proc_0_io_pipe_phv_out_data_58; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_59 = proc_0_io_pipe_phv_out_data_59; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_60 = proc_0_io_pipe_phv_out_data_60; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_61 = proc_0_io_pipe_phv_out_data_61; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_62 = proc_0_io_pipe_phv_out_data_62; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_63 = proc_0_io_pipe_phv_out_data_63; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_64 = proc_0_io_pipe_phv_out_data_64; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_65 = proc_0_io_pipe_phv_out_data_65; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_66 = proc_0_io_pipe_phv_out_data_66; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_67 = proc_0_io_pipe_phv_out_data_67; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_68 = proc_0_io_pipe_phv_out_data_68; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_69 = proc_0_io_pipe_phv_out_data_69; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_70 = proc_0_io_pipe_phv_out_data_70; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_71 = proc_0_io_pipe_phv_out_data_71; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_72 = proc_0_io_pipe_phv_out_data_72; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_73 = proc_0_io_pipe_phv_out_data_73; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_74 = proc_0_io_pipe_phv_out_data_74; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_75 = proc_0_io_pipe_phv_out_data_75; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_76 = proc_0_io_pipe_phv_out_data_76; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_77 = proc_0_io_pipe_phv_out_data_77; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_78 = proc_0_io_pipe_phv_out_data_78; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_79 = proc_0_io_pipe_phv_out_data_79; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_80 = proc_0_io_pipe_phv_out_data_80; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_81 = proc_0_io_pipe_phv_out_data_81; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_82 = proc_0_io_pipe_phv_out_data_82; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_83 = proc_0_io_pipe_phv_out_data_83; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_84 = proc_0_io_pipe_phv_out_data_84; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_85 = proc_0_io_pipe_phv_out_data_85; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_86 = proc_0_io_pipe_phv_out_data_86; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_87 = proc_0_io_pipe_phv_out_data_87; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_88 = proc_0_io_pipe_phv_out_data_88; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_89 = proc_0_io_pipe_phv_out_data_89; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_90 = proc_0_io_pipe_phv_out_data_90; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_91 = proc_0_io_pipe_phv_out_data_91; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_92 = proc_0_io_pipe_phv_out_data_92; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_93 = proc_0_io_pipe_phv_out_data_93; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_94 = proc_0_io_pipe_phv_out_data_94; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_95 = proc_0_io_pipe_phv_out_data_95; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_96 = proc_0_io_pipe_phv_out_data_96; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_97 = proc_0_io_pipe_phv_out_data_97; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_98 = proc_0_io_pipe_phv_out_data_98; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_99 = proc_0_io_pipe_phv_out_data_99; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_100 = proc_0_io_pipe_phv_out_data_100; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_101 = proc_0_io_pipe_phv_out_data_101; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_102 = proc_0_io_pipe_phv_out_data_102; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_103 = proc_0_io_pipe_phv_out_data_103; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_104 = proc_0_io_pipe_phv_out_data_104; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_105 = proc_0_io_pipe_phv_out_data_105; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_106 = proc_0_io_pipe_phv_out_data_106; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_107 = proc_0_io_pipe_phv_out_data_107; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_108 = proc_0_io_pipe_phv_out_data_108; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_109 = proc_0_io_pipe_phv_out_data_109; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_110 = proc_0_io_pipe_phv_out_data_110; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_111 = proc_0_io_pipe_phv_out_data_111; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_112 = proc_0_io_pipe_phv_out_data_112; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_113 = proc_0_io_pipe_phv_out_data_113; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_114 = proc_0_io_pipe_phv_out_data_114; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_115 = proc_0_io_pipe_phv_out_data_115; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_116 = proc_0_io_pipe_phv_out_data_116; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_117 = proc_0_io_pipe_phv_out_data_117; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_118 = proc_0_io_pipe_phv_out_data_118; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_119 = proc_0_io_pipe_phv_out_data_119; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_120 = proc_0_io_pipe_phv_out_data_120; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_121 = proc_0_io_pipe_phv_out_data_121; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_122 = proc_0_io_pipe_phv_out_data_122; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_123 = proc_0_io_pipe_phv_out_data_123; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_124 = proc_0_io_pipe_phv_out_data_124; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_125 = proc_0_io_pipe_phv_out_data_125; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_126 = proc_0_io_pipe_phv_out_data_126; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_127 = proc_0_io_pipe_phv_out_data_127; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_128 = proc_0_io_pipe_phv_out_data_128; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_129 = proc_0_io_pipe_phv_out_data_129; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_130 = proc_0_io_pipe_phv_out_data_130; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_131 = proc_0_io_pipe_phv_out_data_131; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_132 = proc_0_io_pipe_phv_out_data_132; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_133 = proc_0_io_pipe_phv_out_data_133; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_134 = proc_0_io_pipe_phv_out_data_134; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_135 = proc_0_io_pipe_phv_out_data_135; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_136 = proc_0_io_pipe_phv_out_data_136; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_137 = proc_0_io_pipe_phv_out_data_137; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_138 = proc_0_io_pipe_phv_out_data_138; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_139 = proc_0_io_pipe_phv_out_data_139; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_140 = proc_0_io_pipe_phv_out_data_140; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_141 = proc_0_io_pipe_phv_out_data_141; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_142 = proc_0_io_pipe_phv_out_data_142; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_143 = proc_0_io_pipe_phv_out_data_143; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_144 = proc_0_io_pipe_phv_out_data_144; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_145 = proc_0_io_pipe_phv_out_data_145; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_146 = proc_0_io_pipe_phv_out_data_146; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_147 = proc_0_io_pipe_phv_out_data_147; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_148 = proc_0_io_pipe_phv_out_data_148; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_149 = proc_0_io_pipe_phv_out_data_149; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_150 = proc_0_io_pipe_phv_out_data_150; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_151 = proc_0_io_pipe_phv_out_data_151; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_152 = proc_0_io_pipe_phv_out_data_152; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_153 = proc_0_io_pipe_phv_out_data_153; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_154 = proc_0_io_pipe_phv_out_data_154; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_155 = proc_0_io_pipe_phv_out_data_155; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_156 = proc_0_io_pipe_phv_out_data_156; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_157 = proc_0_io_pipe_phv_out_data_157; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_158 = proc_0_io_pipe_phv_out_data_158; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_159 = proc_0_io_pipe_phv_out_data_159; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_header_0 = proc_0_io_pipe_phv_out_header_0; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_header_1 = proc_0_io_pipe_phv_out_header_1; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_header_2 = proc_0_io_pipe_phv_out_header_2; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_header_3 = proc_0_io_pipe_phv_out_header_3; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_header_4 = proc_0_io_pipe_phv_out_header_4; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_header_5 = proc_0_io_pipe_phv_out_header_5; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_header_6 = proc_0_io_pipe_phv_out_header_6; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_header_7 = proc_0_io_pipe_phv_out_header_7; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_header_8 = proc_0_io_pipe_phv_out_header_8; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_header_9 = proc_0_io_pipe_phv_out_header_9; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_header_10 = proc_0_io_pipe_phv_out_header_10; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_header_11 = proc_0_io_pipe_phv_out_header_11; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_header_12 = proc_0_io_pipe_phv_out_header_12; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_header_13 = proc_0_io_pipe_phv_out_header_13; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_header_14 = proc_0_io_pipe_phv_out_header_14; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_header_15 = proc_0_io_pipe_phv_out_header_15; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_parse_current_state = proc_0_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_parse_current_offset = proc_0_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_parse_transition_field = proc_0_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_next_processor_id = proc_0_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_next_config_id = proc_0_io_pipe_phv_out_next_config_id; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_valid = proc_0_io_pipe_phv_out_valid; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_last = proc_0_io_pipe_phv_out_last; // @[ipsa.scala 82:32]
  assign trans_0_io_next_proc_exist = 1'h0; // @[ipsa.scala 80:48]
  assign trans_1_clock = clock;
  assign trans_1_io_pipe_phv_in_data_0 = proc_1_io_pipe_phv_out_data_0; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_1 = proc_1_io_pipe_phv_out_data_1; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_2 = proc_1_io_pipe_phv_out_data_2; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_3 = proc_1_io_pipe_phv_out_data_3; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_4 = proc_1_io_pipe_phv_out_data_4; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_5 = proc_1_io_pipe_phv_out_data_5; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_6 = proc_1_io_pipe_phv_out_data_6; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_7 = proc_1_io_pipe_phv_out_data_7; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_8 = proc_1_io_pipe_phv_out_data_8; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_9 = proc_1_io_pipe_phv_out_data_9; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_10 = proc_1_io_pipe_phv_out_data_10; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_11 = proc_1_io_pipe_phv_out_data_11; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_12 = proc_1_io_pipe_phv_out_data_12; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_13 = proc_1_io_pipe_phv_out_data_13; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_14 = proc_1_io_pipe_phv_out_data_14; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_15 = proc_1_io_pipe_phv_out_data_15; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_16 = proc_1_io_pipe_phv_out_data_16; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_17 = proc_1_io_pipe_phv_out_data_17; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_18 = proc_1_io_pipe_phv_out_data_18; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_19 = proc_1_io_pipe_phv_out_data_19; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_20 = proc_1_io_pipe_phv_out_data_20; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_21 = proc_1_io_pipe_phv_out_data_21; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_22 = proc_1_io_pipe_phv_out_data_22; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_23 = proc_1_io_pipe_phv_out_data_23; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_24 = proc_1_io_pipe_phv_out_data_24; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_25 = proc_1_io_pipe_phv_out_data_25; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_26 = proc_1_io_pipe_phv_out_data_26; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_27 = proc_1_io_pipe_phv_out_data_27; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_28 = proc_1_io_pipe_phv_out_data_28; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_29 = proc_1_io_pipe_phv_out_data_29; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_30 = proc_1_io_pipe_phv_out_data_30; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_31 = proc_1_io_pipe_phv_out_data_31; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_32 = proc_1_io_pipe_phv_out_data_32; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_33 = proc_1_io_pipe_phv_out_data_33; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_34 = proc_1_io_pipe_phv_out_data_34; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_35 = proc_1_io_pipe_phv_out_data_35; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_36 = proc_1_io_pipe_phv_out_data_36; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_37 = proc_1_io_pipe_phv_out_data_37; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_38 = proc_1_io_pipe_phv_out_data_38; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_39 = proc_1_io_pipe_phv_out_data_39; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_40 = proc_1_io_pipe_phv_out_data_40; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_41 = proc_1_io_pipe_phv_out_data_41; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_42 = proc_1_io_pipe_phv_out_data_42; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_43 = proc_1_io_pipe_phv_out_data_43; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_44 = proc_1_io_pipe_phv_out_data_44; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_45 = proc_1_io_pipe_phv_out_data_45; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_46 = proc_1_io_pipe_phv_out_data_46; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_47 = proc_1_io_pipe_phv_out_data_47; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_48 = proc_1_io_pipe_phv_out_data_48; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_49 = proc_1_io_pipe_phv_out_data_49; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_50 = proc_1_io_pipe_phv_out_data_50; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_51 = proc_1_io_pipe_phv_out_data_51; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_52 = proc_1_io_pipe_phv_out_data_52; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_53 = proc_1_io_pipe_phv_out_data_53; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_54 = proc_1_io_pipe_phv_out_data_54; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_55 = proc_1_io_pipe_phv_out_data_55; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_56 = proc_1_io_pipe_phv_out_data_56; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_57 = proc_1_io_pipe_phv_out_data_57; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_58 = proc_1_io_pipe_phv_out_data_58; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_59 = proc_1_io_pipe_phv_out_data_59; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_60 = proc_1_io_pipe_phv_out_data_60; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_61 = proc_1_io_pipe_phv_out_data_61; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_62 = proc_1_io_pipe_phv_out_data_62; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_63 = proc_1_io_pipe_phv_out_data_63; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_64 = proc_1_io_pipe_phv_out_data_64; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_65 = proc_1_io_pipe_phv_out_data_65; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_66 = proc_1_io_pipe_phv_out_data_66; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_67 = proc_1_io_pipe_phv_out_data_67; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_68 = proc_1_io_pipe_phv_out_data_68; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_69 = proc_1_io_pipe_phv_out_data_69; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_70 = proc_1_io_pipe_phv_out_data_70; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_71 = proc_1_io_pipe_phv_out_data_71; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_72 = proc_1_io_pipe_phv_out_data_72; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_73 = proc_1_io_pipe_phv_out_data_73; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_74 = proc_1_io_pipe_phv_out_data_74; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_75 = proc_1_io_pipe_phv_out_data_75; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_76 = proc_1_io_pipe_phv_out_data_76; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_77 = proc_1_io_pipe_phv_out_data_77; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_78 = proc_1_io_pipe_phv_out_data_78; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_79 = proc_1_io_pipe_phv_out_data_79; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_80 = proc_1_io_pipe_phv_out_data_80; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_81 = proc_1_io_pipe_phv_out_data_81; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_82 = proc_1_io_pipe_phv_out_data_82; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_83 = proc_1_io_pipe_phv_out_data_83; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_84 = proc_1_io_pipe_phv_out_data_84; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_85 = proc_1_io_pipe_phv_out_data_85; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_86 = proc_1_io_pipe_phv_out_data_86; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_87 = proc_1_io_pipe_phv_out_data_87; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_88 = proc_1_io_pipe_phv_out_data_88; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_89 = proc_1_io_pipe_phv_out_data_89; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_90 = proc_1_io_pipe_phv_out_data_90; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_91 = proc_1_io_pipe_phv_out_data_91; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_92 = proc_1_io_pipe_phv_out_data_92; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_93 = proc_1_io_pipe_phv_out_data_93; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_94 = proc_1_io_pipe_phv_out_data_94; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_95 = proc_1_io_pipe_phv_out_data_95; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_96 = proc_1_io_pipe_phv_out_data_96; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_97 = proc_1_io_pipe_phv_out_data_97; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_98 = proc_1_io_pipe_phv_out_data_98; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_99 = proc_1_io_pipe_phv_out_data_99; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_100 = proc_1_io_pipe_phv_out_data_100; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_101 = proc_1_io_pipe_phv_out_data_101; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_102 = proc_1_io_pipe_phv_out_data_102; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_103 = proc_1_io_pipe_phv_out_data_103; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_104 = proc_1_io_pipe_phv_out_data_104; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_105 = proc_1_io_pipe_phv_out_data_105; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_106 = proc_1_io_pipe_phv_out_data_106; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_107 = proc_1_io_pipe_phv_out_data_107; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_108 = proc_1_io_pipe_phv_out_data_108; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_109 = proc_1_io_pipe_phv_out_data_109; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_110 = proc_1_io_pipe_phv_out_data_110; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_111 = proc_1_io_pipe_phv_out_data_111; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_112 = proc_1_io_pipe_phv_out_data_112; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_113 = proc_1_io_pipe_phv_out_data_113; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_114 = proc_1_io_pipe_phv_out_data_114; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_115 = proc_1_io_pipe_phv_out_data_115; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_116 = proc_1_io_pipe_phv_out_data_116; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_117 = proc_1_io_pipe_phv_out_data_117; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_118 = proc_1_io_pipe_phv_out_data_118; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_119 = proc_1_io_pipe_phv_out_data_119; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_120 = proc_1_io_pipe_phv_out_data_120; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_121 = proc_1_io_pipe_phv_out_data_121; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_122 = proc_1_io_pipe_phv_out_data_122; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_123 = proc_1_io_pipe_phv_out_data_123; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_124 = proc_1_io_pipe_phv_out_data_124; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_125 = proc_1_io_pipe_phv_out_data_125; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_126 = proc_1_io_pipe_phv_out_data_126; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_127 = proc_1_io_pipe_phv_out_data_127; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_128 = proc_1_io_pipe_phv_out_data_128; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_129 = proc_1_io_pipe_phv_out_data_129; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_130 = proc_1_io_pipe_phv_out_data_130; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_131 = proc_1_io_pipe_phv_out_data_131; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_132 = proc_1_io_pipe_phv_out_data_132; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_133 = proc_1_io_pipe_phv_out_data_133; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_134 = proc_1_io_pipe_phv_out_data_134; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_135 = proc_1_io_pipe_phv_out_data_135; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_136 = proc_1_io_pipe_phv_out_data_136; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_137 = proc_1_io_pipe_phv_out_data_137; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_138 = proc_1_io_pipe_phv_out_data_138; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_139 = proc_1_io_pipe_phv_out_data_139; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_140 = proc_1_io_pipe_phv_out_data_140; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_141 = proc_1_io_pipe_phv_out_data_141; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_142 = proc_1_io_pipe_phv_out_data_142; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_143 = proc_1_io_pipe_phv_out_data_143; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_144 = proc_1_io_pipe_phv_out_data_144; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_145 = proc_1_io_pipe_phv_out_data_145; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_146 = proc_1_io_pipe_phv_out_data_146; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_147 = proc_1_io_pipe_phv_out_data_147; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_148 = proc_1_io_pipe_phv_out_data_148; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_149 = proc_1_io_pipe_phv_out_data_149; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_150 = proc_1_io_pipe_phv_out_data_150; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_151 = proc_1_io_pipe_phv_out_data_151; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_152 = proc_1_io_pipe_phv_out_data_152; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_153 = proc_1_io_pipe_phv_out_data_153; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_154 = proc_1_io_pipe_phv_out_data_154; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_155 = proc_1_io_pipe_phv_out_data_155; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_156 = proc_1_io_pipe_phv_out_data_156; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_157 = proc_1_io_pipe_phv_out_data_157; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_158 = proc_1_io_pipe_phv_out_data_158; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_159 = proc_1_io_pipe_phv_out_data_159; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_header_0 = proc_1_io_pipe_phv_out_header_0; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_header_1 = proc_1_io_pipe_phv_out_header_1; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_header_2 = proc_1_io_pipe_phv_out_header_2; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_header_3 = proc_1_io_pipe_phv_out_header_3; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_header_4 = proc_1_io_pipe_phv_out_header_4; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_header_5 = proc_1_io_pipe_phv_out_header_5; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_header_6 = proc_1_io_pipe_phv_out_header_6; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_header_7 = proc_1_io_pipe_phv_out_header_7; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_header_8 = proc_1_io_pipe_phv_out_header_8; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_header_9 = proc_1_io_pipe_phv_out_header_9; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_header_10 = proc_1_io_pipe_phv_out_header_10; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_header_11 = proc_1_io_pipe_phv_out_header_11; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_header_12 = proc_1_io_pipe_phv_out_header_12; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_header_13 = proc_1_io_pipe_phv_out_header_13; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_header_14 = proc_1_io_pipe_phv_out_header_14; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_header_15 = proc_1_io_pipe_phv_out_header_15; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_parse_current_state = proc_1_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_parse_current_offset = proc_1_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_parse_transition_field = proc_1_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_next_processor_id = proc_1_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_next_config_id = proc_1_io_pipe_phv_out_next_config_id; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_valid = proc_1_io_pipe_phv_out_valid; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_last = proc_1_io_pipe_phv_out_last; // @[ipsa.scala 82:32]
  assign trans_1_io_next_proc_exist = 1'h1; // @[ipsa.scala 80:48]
  assign trans_2_clock = clock;
  assign trans_2_io_pipe_phv_in_data_0 = proc_2_io_pipe_phv_out_data_0; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_1 = proc_2_io_pipe_phv_out_data_1; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_2 = proc_2_io_pipe_phv_out_data_2; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_3 = proc_2_io_pipe_phv_out_data_3; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_4 = proc_2_io_pipe_phv_out_data_4; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_5 = proc_2_io_pipe_phv_out_data_5; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_6 = proc_2_io_pipe_phv_out_data_6; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_7 = proc_2_io_pipe_phv_out_data_7; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_8 = proc_2_io_pipe_phv_out_data_8; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_9 = proc_2_io_pipe_phv_out_data_9; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_10 = proc_2_io_pipe_phv_out_data_10; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_11 = proc_2_io_pipe_phv_out_data_11; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_12 = proc_2_io_pipe_phv_out_data_12; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_13 = proc_2_io_pipe_phv_out_data_13; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_14 = proc_2_io_pipe_phv_out_data_14; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_15 = proc_2_io_pipe_phv_out_data_15; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_16 = proc_2_io_pipe_phv_out_data_16; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_17 = proc_2_io_pipe_phv_out_data_17; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_18 = proc_2_io_pipe_phv_out_data_18; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_19 = proc_2_io_pipe_phv_out_data_19; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_20 = proc_2_io_pipe_phv_out_data_20; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_21 = proc_2_io_pipe_phv_out_data_21; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_22 = proc_2_io_pipe_phv_out_data_22; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_23 = proc_2_io_pipe_phv_out_data_23; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_24 = proc_2_io_pipe_phv_out_data_24; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_25 = proc_2_io_pipe_phv_out_data_25; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_26 = proc_2_io_pipe_phv_out_data_26; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_27 = proc_2_io_pipe_phv_out_data_27; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_28 = proc_2_io_pipe_phv_out_data_28; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_29 = proc_2_io_pipe_phv_out_data_29; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_30 = proc_2_io_pipe_phv_out_data_30; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_31 = proc_2_io_pipe_phv_out_data_31; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_32 = proc_2_io_pipe_phv_out_data_32; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_33 = proc_2_io_pipe_phv_out_data_33; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_34 = proc_2_io_pipe_phv_out_data_34; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_35 = proc_2_io_pipe_phv_out_data_35; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_36 = proc_2_io_pipe_phv_out_data_36; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_37 = proc_2_io_pipe_phv_out_data_37; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_38 = proc_2_io_pipe_phv_out_data_38; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_39 = proc_2_io_pipe_phv_out_data_39; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_40 = proc_2_io_pipe_phv_out_data_40; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_41 = proc_2_io_pipe_phv_out_data_41; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_42 = proc_2_io_pipe_phv_out_data_42; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_43 = proc_2_io_pipe_phv_out_data_43; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_44 = proc_2_io_pipe_phv_out_data_44; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_45 = proc_2_io_pipe_phv_out_data_45; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_46 = proc_2_io_pipe_phv_out_data_46; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_47 = proc_2_io_pipe_phv_out_data_47; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_48 = proc_2_io_pipe_phv_out_data_48; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_49 = proc_2_io_pipe_phv_out_data_49; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_50 = proc_2_io_pipe_phv_out_data_50; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_51 = proc_2_io_pipe_phv_out_data_51; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_52 = proc_2_io_pipe_phv_out_data_52; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_53 = proc_2_io_pipe_phv_out_data_53; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_54 = proc_2_io_pipe_phv_out_data_54; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_55 = proc_2_io_pipe_phv_out_data_55; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_56 = proc_2_io_pipe_phv_out_data_56; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_57 = proc_2_io_pipe_phv_out_data_57; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_58 = proc_2_io_pipe_phv_out_data_58; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_59 = proc_2_io_pipe_phv_out_data_59; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_60 = proc_2_io_pipe_phv_out_data_60; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_61 = proc_2_io_pipe_phv_out_data_61; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_62 = proc_2_io_pipe_phv_out_data_62; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_63 = proc_2_io_pipe_phv_out_data_63; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_64 = proc_2_io_pipe_phv_out_data_64; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_65 = proc_2_io_pipe_phv_out_data_65; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_66 = proc_2_io_pipe_phv_out_data_66; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_67 = proc_2_io_pipe_phv_out_data_67; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_68 = proc_2_io_pipe_phv_out_data_68; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_69 = proc_2_io_pipe_phv_out_data_69; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_70 = proc_2_io_pipe_phv_out_data_70; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_71 = proc_2_io_pipe_phv_out_data_71; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_72 = proc_2_io_pipe_phv_out_data_72; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_73 = proc_2_io_pipe_phv_out_data_73; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_74 = proc_2_io_pipe_phv_out_data_74; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_75 = proc_2_io_pipe_phv_out_data_75; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_76 = proc_2_io_pipe_phv_out_data_76; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_77 = proc_2_io_pipe_phv_out_data_77; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_78 = proc_2_io_pipe_phv_out_data_78; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_79 = proc_2_io_pipe_phv_out_data_79; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_80 = proc_2_io_pipe_phv_out_data_80; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_81 = proc_2_io_pipe_phv_out_data_81; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_82 = proc_2_io_pipe_phv_out_data_82; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_83 = proc_2_io_pipe_phv_out_data_83; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_84 = proc_2_io_pipe_phv_out_data_84; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_85 = proc_2_io_pipe_phv_out_data_85; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_86 = proc_2_io_pipe_phv_out_data_86; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_87 = proc_2_io_pipe_phv_out_data_87; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_88 = proc_2_io_pipe_phv_out_data_88; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_89 = proc_2_io_pipe_phv_out_data_89; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_90 = proc_2_io_pipe_phv_out_data_90; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_91 = proc_2_io_pipe_phv_out_data_91; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_92 = proc_2_io_pipe_phv_out_data_92; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_93 = proc_2_io_pipe_phv_out_data_93; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_94 = proc_2_io_pipe_phv_out_data_94; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_95 = proc_2_io_pipe_phv_out_data_95; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_96 = proc_2_io_pipe_phv_out_data_96; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_97 = proc_2_io_pipe_phv_out_data_97; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_98 = proc_2_io_pipe_phv_out_data_98; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_99 = proc_2_io_pipe_phv_out_data_99; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_100 = proc_2_io_pipe_phv_out_data_100; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_101 = proc_2_io_pipe_phv_out_data_101; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_102 = proc_2_io_pipe_phv_out_data_102; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_103 = proc_2_io_pipe_phv_out_data_103; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_104 = proc_2_io_pipe_phv_out_data_104; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_105 = proc_2_io_pipe_phv_out_data_105; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_106 = proc_2_io_pipe_phv_out_data_106; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_107 = proc_2_io_pipe_phv_out_data_107; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_108 = proc_2_io_pipe_phv_out_data_108; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_109 = proc_2_io_pipe_phv_out_data_109; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_110 = proc_2_io_pipe_phv_out_data_110; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_111 = proc_2_io_pipe_phv_out_data_111; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_112 = proc_2_io_pipe_phv_out_data_112; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_113 = proc_2_io_pipe_phv_out_data_113; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_114 = proc_2_io_pipe_phv_out_data_114; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_115 = proc_2_io_pipe_phv_out_data_115; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_116 = proc_2_io_pipe_phv_out_data_116; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_117 = proc_2_io_pipe_phv_out_data_117; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_118 = proc_2_io_pipe_phv_out_data_118; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_119 = proc_2_io_pipe_phv_out_data_119; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_120 = proc_2_io_pipe_phv_out_data_120; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_121 = proc_2_io_pipe_phv_out_data_121; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_122 = proc_2_io_pipe_phv_out_data_122; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_123 = proc_2_io_pipe_phv_out_data_123; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_124 = proc_2_io_pipe_phv_out_data_124; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_125 = proc_2_io_pipe_phv_out_data_125; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_126 = proc_2_io_pipe_phv_out_data_126; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_127 = proc_2_io_pipe_phv_out_data_127; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_128 = proc_2_io_pipe_phv_out_data_128; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_129 = proc_2_io_pipe_phv_out_data_129; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_130 = proc_2_io_pipe_phv_out_data_130; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_131 = proc_2_io_pipe_phv_out_data_131; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_132 = proc_2_io_pipe_phv_out_data_132; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_133 = proc_2_io_pipe_phv_out_data_133; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_134 = proc_2_io_pipe_phv_out_data_134; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_135 = proc_2_io_pipe_phv_out_data_135; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_136 = proc_2_io_pipe_phv_out_data_136; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_137 = proc_2_io_pipe_phv_out_data_137; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_138 = proc_2_io_pipe_phv_out_data_138; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_139 = proc_2_io_pipe_phv_out_data_139; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_140 = proc_2_io_pipe_phv_out_data_140; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_141 = proc_2_io_pipe_phv_out_data_141; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_142 = proc_2_io_pipe_phv_out_data_142; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_143 = proc_2_io_pipe_phv_out_data_143; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_144 = proc_2_io_pipe_phv_out_data_144; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_145 = proc_2_io_pipe_phv_out_data_145; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_146 = proc_2_io_pipe_phv_out_data_146; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_147 = proc_2_io_pipe_phv_out_data_147; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_148 = proc_2_io_pipe_phv_out_data_148; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_149 = proc_2_io_pipe_phv_out_data_149; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_150 = proc_2_io_pipe_phv_out_data_150; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_151 = proc_2_io_pipe_phv_out_data_151; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_152 = proc_2_io_pipe_phv_out_data_152; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_153 = proc_2_io_pipe_phv_out_data_153; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_154 = proc_2_io_pipe_phv_out_data_154; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_155 = proc_2_io_pipe_phv_out_data_155; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_156 = proc_2_io_pipe_phv_out_data_156; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_157 = proc_2_io_pipe_phv_out_data_157; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_158 = proc_2_io_pipe_phv_out_data_158; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_159 = proc_2_io_pipe_phv_out_data_159; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_header_0 = proc_2_io_pipe_phv_out_header_0; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_header_1 = proc_2_io_pipe_phv_out_header_1; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_header_2 = proc_2_io_pipe_phv_out_header_2; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_header_3 = proc_2_io_pipe_phv_out_header_3; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_header_4 = proc_2_io_pipe_phv_out_header_4; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_header_5 = proc_2_io_pipe_phv_out_header_5; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_header_6 = proc_2_io_pipe_phv_out_header_6; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_header_7 = proc_2_io_pipe_phv_out_header_7; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_header_8 = proc_2_io_pipe_phv_out_header_8; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_header_9 = proc_2_io_pipe_phv_out_header_9; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_header_10 = proc_2_io_pipe_phv_out_header_10; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_header_11 = proc_2_io_pipe_phv_out_header_11; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_header_12 = proc_2_io_pipe_phv_out_header_12; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_header_13 = proc_2_io_pipe_phv_out_header_13; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_header_14 = proc_2_io_pipe_phv_out_header_14; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_header_15 = proc_2_io_pipe_phv_out_header_15; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_parse_current_state = proc_2_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_parse_current_offset = proc_2_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_parse_transition_field = proc_2_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_next_processor_id = proc_2_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_next_config_id = proc_2_io_pipe_phv_out_next_config_id; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_valid = proc_2_io_pipe_phv_out_valid; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_last = proc_2_io_pipe_phv_out_last; // @[ipsa.scala 82:32]
  assign trans_2_io_next_proc_exist = 1'h1; // @[ipsa.scala 80:48]
  assign trans_3_clock = clock;
  assign trans_3_io_pipe_phv_in_data_0 = proc_3_io_pipe_phv_out_data_0; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_1 = proc_3_io_pipe_phv_out_data_1; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_2 = proc_3_io_pipe_phv_out_data_2; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_3 = proc_3_io_pipe_phv_out_data_3; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_4 = proc_3_io_pipe_phv_out_data_4; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_5 = proc_3_io_pipe_phv_out_data_5; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_6 = proc_3_io_pipe_phv_out_data_6; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_7 = proc_3_io_pipe_phv_out_data_7; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_8 = proc_3_io_pipe_phv_out_data_8; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_9 = proc_3_io_pipe_phv_out_data_9; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_10 = proc_3_io_pipe_phv_out_data_10; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_11 = proc_3_io_pipe_phv_out_data_11; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_12 = proc_3_io_pipe_phv_out_data_12; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_13 = proc_3_io_pipe_phv_out_data_13; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_14 = proc_3_io_pipe_phv_out_data_14; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_15 = proc_3_io_pipe_phv_out_data_15; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_16 = proc_3_io_pipe_phv_out_data_16; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_17 = proc_3_io_pipe_phv_out_data_17; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_18 = proc_3_io_pipe_phv_out_data_18; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_19 = proc_3_io_pipe_phv_out_data_19; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_20 = proc_3_io_pipe_phv_out_data_20; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_21 = proc_3_io_pipe_phv_out_data_21; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_22 = proc_3_io_pipe_phv_out_data_22; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_23 = proc_3_io_pipe_phv_out_data_23; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_24 = proc_3_io_pipe_phv_out_data_24; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_25 = proc_3_io_pipe_phv_out_data_25; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_26 = proc_3_io_pipe_phv_out_data_26; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_27 = proc_3_io_pipe_phv_out_data_27; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_28 = proc_3_io_pipe_phv_out_data_28; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_29 = proc_3_io_pipe_phv_out_data_29; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_30 = proc_3_io_pipe_phv_out_data_30; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_31 = proc_3_io_pipe_phv_out_data_31; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_32 = proc_3_io_pipe_phv_out_data_32; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_33 = proc_3_io_pipe_phv_out_data_33; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_34 = proc_3_io_pipe_phv_out_data_34; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_35 = proc_3_io_pipe_phv_out_data_35; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_36 = proc_3_io_pipe_phv_out_data_36; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_37 = proc_3_io_pipe_phv_out_data_37; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_38 = proc_3_io_pipe_phv_out_data_38; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_39 = proc_3_io_pipe_phv_out_data_39; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_40 = proc_3_io_pipe_phv_out_data_40; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_41 = proc_3_io_pipe_phv_out_data_41; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_42 = proc_3_io_pipe_phv_out_data_42; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_43 = proc_3_io_pipe_phv_out_data_43; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_44 = proc_3_io_pipe_phv_out_data_44; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_45 = proc_3_io_pipe_phv_out_data_45; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_46 = proc_3_io_pipe_phv_out_data_46; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_47 = proc_3_io_pipe_phv_out_data_47; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_48 = proc_3_io_pipe_phv_out_data_48; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_49 = proc_3_io_pipe_phv_out_data_49; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_50 = proc_3_io_pipe_phv_out_data_50; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_51 = proc_3_io_pipe_phv_out_data_51; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_52 = proc_3_io_pipe_phv_out_data_52; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_53 = proc_3_io_pipe_phv_out_data_53; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_54 = proc_3_io_pipe_phv_out_data_54; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_55 = proc_3_io_pipe_phv_out_data_55; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_56 = proc_3_io_pipe_phv_out_data_56; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_57 = proc_3_io_pipe_phv_out_data_57; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_58 = proc_3_io_pipe_phv_out_data_58; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_59 = proc_3_io_pipe_phv_out_data_59; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_60 = proc_3_io_pipe_phv_out_data_60; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_61 = proc_3_io_pipe_phv_out_data_61; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_62 = proc_3_io_pipe_phv_out_data_62; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_63 = proc_3_io_pipe_phv_out_data_63; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_64 = proc_3_io_pipe_phv_out_data_64; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_65 = proc_3_io_pipe_phv_out_data_65; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_66 = proc_3_io_pipe_phv_out_data_66; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_67 = proc_3_io_pipe_phv_out_data_67; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_68 = proc_3_io_pipe_phv_out_data_68; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_69 = proc_3_io_pipe_phv_out_data_69; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_70 = proc_3_io_pipe_phv_out_data_70; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_71 = proc_3_io_pipe_phv_out_data_71; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_72 = proc_3_io_pipe_phv_out_data_72; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_73 = proc_3_io_pipe_phv_out_data_73; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_74 = proc_3_io_pipe_phv_out_data_74; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_75 = proc_3_io_pipe_phv_out_data_75; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_76 = proc_3_io_pipe_phv_out_data_76; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_77 = proc_3_io_pipe_phv_out_data_77; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_78 = proc_3_io_pipe_phv_out_data_78; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_79 = proc_3_io_pipe_phv_out_data_79; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_80 = proc_3_io_pipe_phv_out_data_80; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_81 = proc_3_io_pipe_phv_out_data_81; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_82 = proc_3_io_pipe_phv_out_data_82; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_83 = proc_3_io_pipe_phv_out_data_83; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_84 = proc_3_io_pipe_phv_out_data_84; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_85 = proc_3_io_pipe_phv_out_data_85; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_86 = proc_3_io_pipe_phv_out_data_86; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_87 = proc_3_io_pipe_phv_out_data_87; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_88 = proc_3_io_pipe_phv_out_data_88; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_89 = proc_3_io_pipe_phv_out_data_89; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_90 = proc_3_io_pipe_phv_out_data_90; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_91 = proc_3_io_pipe_phv_out_data_91; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_92 = proc_3_io_pipe_phv_out_data_92; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_93 = proc_3_io_pipe_phv_out_data_93; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_94 = proc_3_io_pipe_phv_out_data_94; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_95 = proc_3_io_pipe_phv_out_data_95; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_96 = proc_3_io_pipe_phv_out_data_96; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_97 = proc_3_io_pipe_phv_out_data_97; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_98 = proc_3_io_pipe_phv_out_data_98; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_99 = proc_3_io_pipe_phv_out_data_99; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_100 = proc_3_io_pipe_phv_out_data_100; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_101 = proc_3_io_pipe_phv_out_data_101; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_102 = proc_3_io_pipe_phv_out_data_102; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_103 = proc_3_io_pipe_phv_out_data_103; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_104 = proc_3_io_pipe_phv_out_data_104; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_105 = proc_3_io_pipe_phv_out_data_105; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_106 = proc_3_io_pipe_phv_out_data_106; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_107 = proc_3_io_pipe_phv_out_data_107; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_108 = proc_3_io_pipe_phv_out_data_108; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_109 = proc_3_io_pipe_phv_out_data_109; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_110 = proc_3_io_pipe_phv_out_data_110; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_111 = proc_3_io_pipe_phv_out_data_111; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_112 = proc_3_io_pipe_phv_out_data_112; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_113 = proc_3_io_pipe_phv_out_data_113; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_114 = proc_3_io_pipe_phv_out_data_114; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_115 = proc_3_io_pipe_phv_out_data_115; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_116 = proc_3_io_pipe_phv_out_data_116; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_117 = proc_3_io_pipe_phv_out_data_117; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_118 = proc_3_io_pipe_phv_out_data_118; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_119 = proc_3_io_pipe_phv_out_data_119; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_120 = proc_3_io_pipe_phv_out_data_120; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_121 = proc_3_io_pipe_phv_out_data_121; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_122 = proc_3_io_pipe_phv_out_data_122; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_123 = proc_3_io_pipe_phv_out_data_123; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_124 = proc_3_io_pipe_phv_out_data_124; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_125 = proc_3_io_pipe_phv_out_data_125; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_126 = proc_3_io_pipe_phv_out_data_126; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_127 = proc_3_io_pipe_phv_out_data_127; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_128 = proc_3_io_pipe_phv_out_data_128; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_129 = proc_3_io_pipe_phv_out_data_129; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_130 = proc_3_io_pipe_phv_out_data_130; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_131 = proc_3_io_pipe_phv_out_data_131; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_132 = proc_3_io_pipe_phv_out_data_132; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_133 = proc_3_io_pipe_phv_out_data_133; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_134 = proc_3_io_pipe_phv_out_data_134; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_135 = proc_3_io_pipe_phv_out_data_135; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_136 = proc_3_io_pipe_phv_out_data_136; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_137 = proc_3_io_pipe_phv_out_data_137; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_138 = proc_3_io_pipe_phv_out_data_138; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_139 = proc_3_io_pipe_phv_out_data_139; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_140 = proc_3_io_pipe_phv_out_data_140; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_141 = proc_3_io_pipe_phv_out_data_141; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_142 = proc_3_io_pipe_phv_out_data_142; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_143 = proc_3_io_pipe_phv_out_data_143; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_144 = proc_3_io_pipe_phv_out_data_144; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_145 = proc_3_io_pipe_phv_out_data_145; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_146 = proc_3_io_pipe_phv_out_data_146; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_147 = proc_3_io_pipe_phv_out_data_147; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_148 = proc_3_io_pipe_phv_out_data_148; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_149 = proc_3_io_pipe_phv_out_data_149; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_150 = proc_3_io_pipe_phv_out_data_150; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_151 = proc_3_io_pipe_phv_out_data_151; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_152 = proc_3_io_pipe_phv_out_data_152; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_153 = proc_3_io_pipe_phv_out_data_153; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_154 = proc_3_io_pipe_phv_out_data_154; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_155 = proc_3_io_pipe_phv_out_data_155; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_156 = proc_3_io_pipe_phv_out_data_156; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_157 = proc_3_io_pipe_phv_out_data_157; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_158 = proc_3_io_pipe_phv_out_data_158; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_159 = proc_3_io_pipe_phv_out_data_159; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_header_0 = proc_3_io_pipe_phv_out_header_0; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_header_1 = proc_3_io_pipe_phv_out_header_1; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_header_2 = proc_3_io_pipe_phv_out_header_2; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_header_3 = proc_3_io_pipe_phv_out_header_3; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_header_4 = proc_3_io_pipe_phv_out_header_4; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_header_5 = proc_3_io_pipe_phv_out_header_5; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_header_6 = proc_3_io_pipe_phv_out_header_6; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_header_7 = proc_3_io_pipe_phv_out_header_7; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_header_8 = proc_3_io_pipe_phv_out_header_8; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_header_9 = proc_3_io_pipe_phv_out_header_9; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_header_10 = proc_3_io_pipe_phv_out_header_10; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_header_11 = proc_3_io_pipe_phv_out_header_11; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_header_12 = proc_3_io_pipe_phv_out_header_12; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_header_13 = proc_3_io_pipe_phv_out_header_13; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_header_14 = proc_3_io_pipe_phv_out_header_14; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_header_15 = proc_3_io_pipe_phv_out_header_15; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_parse_current_state = proc_3_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_parse_current_offset = proc_3_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_parse_transition_field = proc_3_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_next_processor_id = proc_3_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_next_config_id = proc_3_io_pipe_phv_out_next_config_id; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_valid = proc_3_io_pipe_phv_out_valid; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_last = proc_3_io_pipe_phv_out_last; // @[ipsa.scala 82:32]
  assign trans_3_io_next_proc_exist = 1'h1; // @[ipsa.scala 80:48]
  assign trans_4_clock = clock;
  assign trans_4_io_pipe_phv_in_data_0 = proc_4_io_pipe_phv_out_data_0; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_1 = proc_4_io_pipe_phv_out_data_1; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_2 = proc_4_io_pipe_phv_out_data_2; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_3 = proc_4_io_pipe_phv_out_data_3; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_4 = proc_4_io_pipe_phv_out_data_4; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_5 = proc_4_io_pipe_phv_out_data_5; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_6 = proc_4_io_pipe_phv_out_data_6; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_7 = proc_4_io_pipe_phv_out_data_7; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_8 = proc_4_io_pipe_phv_out_data_8; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_9 = proc_4_io_pipe_phv_out_data_9; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_10 = proc_4_io_pipe_phv_out_data_10; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_11 = proc_4_io_pipe_phv_out_data_11; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_12 = proc_4_io_pipe_phv_out_data_12; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_13 = proc_4_io_pipe_phv_out_data_13; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_14 = proc_4_io_pipe_phv_out_data_14; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_15 = proc_4_io_pipe_phv_out_data_15; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_16 = proc_4_io_pipe_phv_out_data_16; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_17 = proc_4_io_pipe_phv_out_data_17; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_18 = proc_4_io_pipe_phv_out_data_18; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_19 = proc_4_io_pipe_phv_out_data_19; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_20 = proc_4_io_pipe_phv_out_data_20; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_21 = proc_4_io_pipe_phv_out_data_21; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_22 = proc_4_io_pipe_phv_out_data_22; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_23 = proc_4_io_pipe_phv_out_data_23; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_24 = proc_4_io_pipe_phv_out_data_24; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_25 = proc_4_io_pipe_phv_out_data_25; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_26 = proc_4_io_pipe_phv_out_data_26; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_27 = proc_4_io_pipe_phv_out_data_27; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_28 = proc_4_io_pipe_phv_out_data_28; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_29 = proc_4_io_pipe_phv_out_data_29; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_30 = proc_4_io_pipe_phv_out_data_30; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_31 = proc_4_io_pipe_phv_out_data_31; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_32 = proc_4_io_pipe_phv_out_data_32; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_33 = proc_4_io_pipe_phv_out_data_33; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_34 = proc_4_io_pipe_phv_out_data_34; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_35 = proc_4_io_pipe_phv_out_data_35; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_36 = proc_4_io_pipe_phv_out_data_36; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_37 = proc_4_io_pipe_phv_out_data_37; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_38 = proc_4_io_pipe_phv_out_data_38; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_39 = proc_4_io_pipe_phv_out_data_39; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_40 = proc_4_io_pipe_phv_out_data_40; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_41 = proc_4_io_pipe_phv_out_data_41; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_42 = proc_4_io_pipe_phv_out_data_42; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_43 = proc_4_io_pipe_phv_out_data_43; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_44 = proc_4_io_pipe_phv_out_data_44; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_45 = proc_4_io_pipe_phv_out_data_45; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_46 = proc_4_io_pipe_phv_out_data_46; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_47 = proc_4_io_pipe_phv_out_data_47; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_48 = proc_4_io_pipe_phv_out_data_48; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_49 = proc_4_io_pipe_phv_out_data_49; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_50 = proc_4_io_pipe_phv_out_data_50; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_51 = proc_4_io_pipe_phv_out_data_51; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_52 = proc_4_io_pipe_phv_out_data_52; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_53 = proc_4_io_pipe_phv_out_data_53; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_54 = proc_4_io_pipe_phv_out_data_54; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_55 = proc_4_io_pipe_phv_out_data_55; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_56 = proc_4_io_pipe_phv_out_data_56; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_57 = proc_4_io_pipe_phv_out_data_57; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_58 = proc_4_io_pipe_phv_out_data_58; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_59 = proc_4_io_pipe_phv_out_data_59; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_60 = proc_4_io_pipe_phv_out_data_60; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_61 = proc_4_io_pipe_phv_out_data_61; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_62 = proc_4_io_pipe_phv_out_data_62; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_63 = proc_4_io_pipe_phv_out_data_63; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_64 = proc_4_io_pipe_phv_out_data_64; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_65 = proc_4_io_pipe_phv_out_data_65; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_66 = proc_4_io_pipe_phv_out_data_66; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_67 = proc_4_io_pipe_phv_out_data_67; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_68 = proc_4_io_pipe_phv_out_data_68; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_69 = proc_4_io_pipe_phv_out_data_69; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_70 = proc_4_io_pipe_phv_out_data_70; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_71 = proc_4_io_pipe_phv_out_data_71; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_72 = proc_4_io_pipe_phv_out_data_72; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_73 = proc_4_io_pipe_phv_out_data_73; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_74 = proc_4_io_pipe_phv_out_data_74; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_75 = proc_4_io_pipe_phv_out_data_75; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_76 = proc_4_io_pipe_phv_out_data_76; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_77 = proc_4_io_pipe_phv_out_data_77; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_78 = proc_4_io_pipe_phv_out_data_78; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_79 = proc_4_io_pipe_phv_out_data_79; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_80 = proc_4_io_pipe_phv_out_data_80; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_81 = proc_4_io_pipe_phv_out_data_81; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_82 = proc_4_io_pipe_phv_out_data_82; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_83 = proc_4_io_pipe_phv_out_data_83; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_84 = proc_4_io_pipe_phv_out_data_84; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_85 = proc_4_io_pipe_phv_out_data_85; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_86 = proc_4_io_pipe_phv_out_data_86; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_87 = proc_4_io_pipe_phv_out_data_87; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_88 = proc_4_io_pipe_phv_out_data_88; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_89 = proc_4_io_pipe_phv_out_data_89; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_90 = proc_4_io_pipe_phv_out_data_90; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_91 = proc_4_io_pipe_phv_out_data_91; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_92 = proc_4_io_pipe_phv_out_data_92; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_93 = proc_4_io_pipe_phv_out_data_93; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_94 = proc_4_io_pipe_phv_out_data_94; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_95 = proc_4_io_pipe_phv_out_data_95; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_96 = proc_4_io_pipe_phv_out_data_96; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_97 = proc_4_io_pipe_phv_out_data_97; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_98 = proc_4_io_pipe_phv_out_data_98; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_99 = proc_4_io_pipe_phv_out_data_99; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_100 = proc_4_io_pipe_phv_out_data_100; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_101 = proc_4_io_pipe_phv_out_data_101; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_102 = proc_4_io_pipe_phv_out_data_102; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_103 = proc_4_io_pipe_phv_out_data_103; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_104 = proc_4_io_pipe_phv_out_data_104; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_105 = proc_4_io_pipe_phv_out_data_105; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_106 = proc_4_io_pipe_phv_out_data_106; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_107 = proc_4_io_pipe_phv_out_data_107; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_108 = proc_4_io_pipe_phv_out_data_108; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_109 = proc_4_io_pipe_phv_out_data_109; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_110 = proc_4_io_pipe_phv_out_data_110; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_111 = proc_4_io_pipe_phv_out_data_111; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_112 = proc_4_io_pipe_phv_out_data_112; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_113 = proc_4_io_pipe_phv_out_data_113; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_114 = proc_4_io_pipe_phv_out_data_114; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_115 = proc_4_io_pipe_phv_out_data_115; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_116 = proc_4_io_pipe_phv_out_data_116; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_117 = proc_4_io_pipe_phv_out_data_117; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_118 = proc_4_io_pipe_phv_out_data_118; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_119 = proc_4_io_pipe_phv_out_data_119; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_120 = proc_4_io_pipe_phv_out_data_120; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_121 = proc_4_io_pipe_phv_out_data_121; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_122 = proc_4_io_pipe_phv_out_data_122; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_123 = proc_4_io_pipe_phv_out_data_123; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_124 = proc_4_io_pipe_phv_out_data_124; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_125 = proc_4_io_pipe_phv_out_data_125; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_126 = proc_4_io_pipe_phv_out_data_126; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_127 = proc_4_io_pipe_phv_out_data_127; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_128 = proc_4_io_pipe_phv_out_data_128; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_129 = proc_4_io_pipe_phv_out_data_129; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_130 = proc_4_io_pipe_phv_out_data_130; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_131 = proc_4_io_pipe_phv_out_data_131; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_132 = proc_4_io_pipe_phv_out_data_132; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_133 = proc_4_io_pipe_phv_out_data_133; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_134 = proc_4_io_pipe_phv_out_data_134; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_135 = proc_4_io_pipe_phv_out_data_135; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_136 = proc_4_io_pipe_phv_out_data_136; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_137 = proc_4_io_pipe_phv_out_data_137; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_138 = proc_4_io_pipe_phv_out_data_138; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_139 = proc_4_io_pipe_phv_out_data_139; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_140 = proc_4_io_pipe_phv_out_data_140; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_141 = proc_4_io_pipe_phv_out_data_141; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_142 = proc_4_io_pipe_phv_out_data_142; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_143 = proc_4_io_pipe_phv_out_data_143; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_144 = proc_4_io_pipe_phv_out_data_144; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_145 = proc_4_io_pipe_phv_out_data_145; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_146 = proc_4_io_pipe_phv_out_data_146; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_147 = proc_4_io_pipe_phv_out_data_147; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_148 = proc_4_io_pipe_phv_out_data_148; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_149 = proc_4_io_pipe_phv_out_data_149; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_150 = proc_4_io_pipe_phv_out_data_150; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_151 = proc_4_io_pipe_phv_out_data_151; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_152 = proc_4_io_pipe_phv_out_data_152; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_153 = proc_4_io_pipe_phv_out_data_153; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_154 = proc_4_io_pipe_phv_out_data_154; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_155 = proc_4_io_pipe_phv_out_data_155; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_156 = proc_4_io_pipe_phv_out_data_156; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_157 = proc_4_io_pipe_phv_out_data_157; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_158 = proc_4_io_pipe_phv_out_data_158; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_data_159 = proc_4_io_pipe_phv_out_data_159; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_header_0 = proc_4_io_pipe_phv_out_header_0; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_header_1 = proc_4_io_pipe_phv_out_header_1; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_header_2 = proc_4_io_pipe_phv_out_header_2; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_header_3 = proc_4_io_pipe_phv_out_header_3; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_header_4 = proc_4_io_pipe_phv_out_header_4; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_header_5 = proc_4_io_pipe_phv_out_header_5; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_header_6 = proc_4_io_pipe_phv_out_header_6; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_header_7 = proc_4_io_pipe_phv_out_header_7; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_header_8 = proc_4_io_pipe_phv_out_header_8; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_header_9 = proc_4_io_pipe_phv_out_header_9; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_header_10 = proc_4_io_pipe_phv_out_header_10; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_header_11 = proc_4_io_pipe_phv_out_header_11; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_header_12 = proc_4_io_pipe_phv_out_header_12; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_header_13 = proc_4_io_pipe_phv_out_header_13; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_header_14 = proc_4_io_pipe_phv_out_header_14; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_header_15 = proc_4_io_pipe_phv_out_header_15; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_parse_current_state = proc_4_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_parse_current_offset = proc_4_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_parse_transition_field = proc_4_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_next_processor_id = proc_4_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_next_config_id = proc_4_io_pipe_phv_out_next_config_id; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_valid = proc_4_io_pipe_phv_out_valid; // @[ipsa.scala 82:32]
  assign trans_4_io_pipe_phv_in_last = proc_4_io_pipe_phv_out_last; // @[ipsa.scala 82:32]
  assign trans_4_io_next_proc_exist = 1'h1; // @[ipsa.scala 80:48]
  assign trans_5_clock = clock;
  assign trans_5_io_pipe_phv_in_data_0 = proc_5_io_pipe_phv_out_data_0; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_1 = proc_5_io_pipe_phv_out_data_1; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_2 = proc_5_io_pipe_phv_out_data_2; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_3 = proc_5_io_pipe_phv_out_data_3; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_4 = proc_5_io_pipe_phv_out_data_4; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_5 = proc_5_io_pipe_phv_out_data_5; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_6 = proc_5_io_pipe_phv_out_data_6; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_7 = proc_5_io_pipe_phv_out_data_7; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_8 = proc_5_io_pipe_phv_out_data_8; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_9 = proc_5_io_pipe_phv_out_data_9; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_10 = proc_5_io_pipe_phv_out_data_10; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_11 = proc_5_io_pipe_phv_out_data_11; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_12 = proc_5_io_pipe_phv_out_data_12; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_13 = proc_5_io_pipe_phv_out_data_13; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_14 = proc_5_io_pipe_phv_out_data_14; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_15 = proc_5_io_pipe_phv_out_data_15; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_16 = proc_5_io_pipe_phv_out_data_16; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_17 = proc_5_io_pipe_phv_out_data_17; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_18 = proc_5_io_pipe_phv_out_data_18; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_19 = proc_5_io_pipe_phv_out_data_19; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_20 = proc_5_io_pipe_phv_out_data_20; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_21 = proc_5_io_pipe_phv_out_data_21; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_22 = proc_5_io_pipe_phv_out_data_22; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_23 = proc_5_io_pipe_phv_out_data_23; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_24 = proc_5_io_pipe_phv_out_data_24; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_25 = proc_5_io_pipe_phv_out_data_25; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_26 = proc_5_io_pipe_phv_out_data_26; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_27 = proc_5_io_pipe_phv_out_data_27; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_28 = proc_5_io_pipe_phv_out_data_28; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_29 = proc_5_io_pipe_phv_out_data_29; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_30 = proc_5_io_pipe_phv_out_data_30; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_31 = proc_5_io_pipe_phv_out_data_31; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_32 = proc_5_io_pipe_phv_out_data_32; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_33 = proc_5_io_pipe_phv_out_data_33; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_34 = proc_5_io_pipe_phv_out_data_34; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_35 = proc_5_io_pipe_phv_out_data_35; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_36 = proc_5_io_pipe_phv_out_data_36; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_37 = proc_5_io_pipe_phv_out_data_37; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_38 = proc_5_io_pipe_phv_out_data_38; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_39 = proc_5_io_pipe_phv_out_data_39; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_40 = proc_5_io_pipe_phv_out_data_40; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_41 = proc_5_io_pipe_phv_out_data_41; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_42 = proc_5_io_pipe_phv_out_data_42; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_43 = proc_5_io_pipe_phv_out_data_43; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_44 = proc_5_io_pipe_phv_out_data_44; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_45 = proc_5_io_pipe_phv_out_data_45; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_46 = proc_5_io_pipe_phv_out_data_46; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_47 = proc_5_io_pipe_phv_out_data_47; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_48 = proc_5_io_pipe_phv_out_data_48; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_49 = proc_5_io_pipe_phv_out_data_49; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_50 = proc_5_io_pipe_phv_out_data_50; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_51 = proc_5_io_pipe_phv_out_data_51; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_52 = proc_5_io_pipe_phv_out_data_52; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_53 = proc_5_io_pipe_phv_out_data_53; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_54 = proc_5_io_pipe_phv_out_data_54; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_55 = proc_5_io_pipe_phv_out_data_55; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_56 = proc_5_io_pipe_phv_out_data_56; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_57 = proc_5_io_pipe_phv_out_data_57; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_58 = proc_5_io_pipe_phv_out_data_58; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_59 = proc_5_io_pipe_phv_out_data_59; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_60 = proc_5_io_pipe_phv_out_data_60; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_61 = proc_5_io_pipe_phv_out_data_61; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_62 = proc_5_io_pipe_phv_out_data_62; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_63 = proc_5_io_pipe_phv_out_data_63; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_64 = proc_5_io_pipe_phv_out_data_64; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_65 = proc_5_io_pipe_phv_out_data_65; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_66 = proc_5_io_pipe_phv_out_data_66; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_67 = proc_5_io_pipe_phv_out_data_67; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_68 = proc_5_io_pipe_phv_out_data_68; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_69 = proc_5_io_pipe_phv_out_data_69; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_70 = proc_5_io_pipe_phv_out_data_70; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_71 = proc_5_io_pipe_phv_out_data_71; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_72 = proc_5_io_pipe_phv_out_data_72; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_73 = proc_5_io_pipe_phv_out_data_73; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_74 = proc_5_io_pipe_phv_out_data_74; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_75 = proc_5_io_pipe_phv_out_data_75; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_76 = proc_5_io_pipe_phv_out_data_76; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_77 = proc_5_io_pipe_phv_out_data_77; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_78 = proc_5_io_pipe_phv_out_data_78; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_79 = proc_5_io_pipe_phv_out_data_79; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_80 = proc_5_io_pipe_phv_out_data_80; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_81 = proc_5_io_pipe_phv_out_data_81; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_82 = proc_5_io_pipe_phv_out_data_82; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_83 = proc_5_io_pipe_phv_out_data_83; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_84 = proc_5_io_pipe_phv_out_data_84; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_85 = proc_5_io_pipe_phv_out_data_85; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_86 = proc_5_io_pipe_phv_out_data_86; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_87 = proc_5_io_pipe_phv_out_data_87; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_88 = proc_5_io_pipe_phv_out_data_88; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_89 = proc_5_io_pipe_phv_out_data_89; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_90 = proc_5_io_pipe_phv_out_data_90; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_91 = proc_5_io_pipe_phv_out_data_91; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_92 = proc_5_io_pipe_phv_out_data_92; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_93 = proc_5_io_pipe_phv_out_data_93; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_94 = proc_5_io_pipe_phv_out_data_94; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_95 = proc_5_io_pipe_phv_out_data_95; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_96 = proc_5_io_pipe_phv_out_data_96; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_97 = proc_5_io_pipe_phv_out_data_97; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_98 = proc_5_io_pipe_phv_out_data_98; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_99 = proc_5_io_pipe_phv_out_data_99; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_100 = proc_5_io_pipe_phv_out_data_100; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_101 = proc_5_io_pipe_phv_out_data_101; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_102 = proc_5_io_pipe_phv_out_data_102; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_103 = proc_5_io_pipe_phv_out_data_103; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_104 = proc_5_io_pipe_phv_out_data_104; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_105 = proc_5_io_pipe_phv_out_data_105; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_106 = proc_5_io_pipe_phv_out_data_106; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_107 = proc_5_io_pipe_phv_out_data_107; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_108 = proc_5_io_pipe_phv_out_data_108; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_109 = proc_5_io_pipe_phv_out_data_109; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_110 = proc_5_io_pipe_phv_out_data_110; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_111 = proc_5_io_pipe_phv_out_data_111; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_112 = proc_5_io_pipe_phv_out_data_112; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_113 = proc_5_io_pipe_phv_out_data_113; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_114 = proc_5_io_pipe_phv_out_data_114; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_115 = proc_5_io_pipe_phv_out_data_115; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_116 = proc_5_io_pipe_phv_out_data_116; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_117 = proc_5_io_pipe_phv_out_data_117; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_118 = proc_5_io_pipe_phv_out_data_118; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_119 = proc_5_io_pipe_phv_out_data_119; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_120 = proc_5_io_pipe_phv_out_data_120; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_121 = proc_5_io_pipe_phv_out_data_121; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_122 = proc_5_io_pipe_phv_out_data_122; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_123 = proc_5_io_pipe_phv_out_data_123; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_124 = proc_5_io_pipe_phv_out_data_124; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_125 = proc_5_io_pipe_phv_out_data_125; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_126 = proc_5_io_pipe_phv_out_data_126; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_127 = proc_5_io_pipe_phv_out_data_127; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_128 = proc_5_io_pipe_phv_out_data_128; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_129 = proc_5_io_pipe_phv_out_data_129; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_130 = proc_5_io_pipe_phv_out_data_130; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_131 = proc_5_io_pipe_phv_out_data_131; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_132 = proc_5_io_pipe_phv_out_data_132; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_133 = proc_5_io_pipe_phv_out_data_133; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_134 = proc_5_io_pipe_phv_out_data_134; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_135 = proc_5_io_pipe_phv_out_data_135; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_136 = proc_5_io_pipe_phv_out_data_136; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_137 = proc_5_io_pipe_phv_out_data_137; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_138 = proc_5_io_pipe_phv_out_data_138; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_139 = proc_5_io_pipe_phv_out_data_139; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_140 = proc_5_io_pipe_phv_out_data_140; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_141 = proc_5_io_pipe_phv_out_data_141; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_142 = proc_5_io_pipe_phv_out_data_142; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_143 = proc_5_io_pipe_phv_out_data_143; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_144 = proc_5_io_pipe_phv_out_data_144; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_145 = proc_5_io_pipe_phv_out_data_145; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_146 = proc_5_io_pipe_phv_out_data_146; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_147 = proc_5_io_pipe_phv_out_data_147; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_148 = proc_5_io_pipe_phv_out_data_148; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_149 = proc_5_io_pipe_phv_out_data_149; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_150 = proc_5_io_pipe_phv_out_data_150; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_151 = proc_5_io_pipe_phv_out_data_151; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_152 = proc_5_io_pipe_phv_out_data_152; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_153 = proc_5_io_pipe_phv_out_data_153; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_154 = proc_5_io_pipe_phv_out_data_154; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_155 = proc_5_io_pipe_phv_out_data_155; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_156 = proc_5_io_pipe_phv_out_data_156; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_157 = proc_5_io_pipe_phv_out_data_157; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_158 = proc_5_io_pipe_phv_out_data_158; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_data_159 = proc_5_io_pipe_phv_out_data_159; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_header_0 = proc_5_io_pipe_phv_out_header_0; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_header_1 = proc_5_io_pipe_phv_out_header_1; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_header_2 = proc_5_io_pipe_phv_out_header_2; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_header_3 = proc_5_io_pipe_phv_out_header_3; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_header_4 = proc_5_io_pipe_phv_out_header_4; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_header_5 = proc_5_io_pipe_phv_out_header_5; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_header_6 = proc_5_io_pipe_phv_out_header_6; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_header_7 = proc_5_io_pipe_phv_out_header_7; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_header_8 = proc_5_io_pipe_phv_out_header_8; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_header_9 = proc_5_io_pipe_phv_out_header_9; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_header_10 = proc_5_io_pipe_phv_out_header_10; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_header_11 = proc_5_io_pipe_phv_out_header_11; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_header_12 = proc_5_io_pipe_phv_out_header_12; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_header_13 = proc_5_io_pipe_phv_out_header_13; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_header_14 = proc_5_io_pipe_phv_out_header_14; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_header_15 = proc_5_io_pipe_phv_out_header_15; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_parse_current_state = proc_5_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_parse_current_offset = proc_5_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_parse_transition_field = proc_5_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_next_processor_id = proc_5_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_next_config_id = proc_5_io_pipe_phv_out_next_config_id; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_valid = proc_5_io_pipe_phv_out_valid; // @[ipsa.scala 82:32]
  assign trans_5_io_pipe_phv_in_last = proc_5_io_pipe_phv_out_last; // @[ipsa.scala 82:32]
  assign trans_5_io_next_proc_exist = 1'h1; // @[ipsa.scala 80:48]
  assign trans_6_clock = clock;
  assign trans_6_io_pipe_phv_in_data_0 = proc_6_io_pipe_phv_out_data_0; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_1 = proc_6_io_pipe_phv_out_data_1; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_2 = proc_6_io_pipe_phv_out_data_2; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_3 = proc_6_io_pipe_phv_out_data_3; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_4 = proc_6_io_pipe_phv_out_data_4; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_5 = proc_6_io_pipe_phv_out_data_5; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_6 = proc_6_io_pipe_phv_out_data_6; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_7 = proc_6_io_pipe_phv_out_data_7; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_8 = proc_6_io_pipe_phv_out_data_8; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_9 = proc_6_io_pipe_phv_out_data_9; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_10 = proc_6_io_pipe_phv_out_data_10; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_11 = proc_6_io_pipe_phv_out_data_11; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_12 = proc_6_io_pipe_phv_out_data_12; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_13 = proc_6_io_pipe_phv_out_data_13; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_14 = proc_6_io_pipe_phv_out_data_14; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_15 = proc_6_io_pipe_phv_out_data_15; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_16 = proc_6_io_pipe_phv_out_data_16; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_17 = proc_6_io_pipe_phv_out_data_17; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_18 = proc_6_io_pipe_phv_out_data_18; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_19 = proc_6_io_pipe_phv_out_data_19; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_20 = proc_6_io_pipe_phv_out_data_20; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_21 = proc_6_io_pipe_phv_out_data_21; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_22 = proc_6_io_pipe_phv_out_data_22; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_23 = proc_6_io_pipe_phv_out_data_23; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_24 = proc_6_io_pipe_phv_out_data_24; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_25 = proc_6_io_pipe_phv_out_data_25; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_26 = proc_6_io_pipe_phv_out_data_26; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_27 = proc_6_io_pipe_phv_out_data_27; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_28 = proc_6_io_pipe_phv_out_data_28; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_29 = proc_6_io_pipe_phv_out_data_29; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_30 = proc_6_io_pipe_phv_out_data_30; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_31 = proc_6_io_pipe_phv_out_data_31; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_32 = proc_6_io_pipe_phv_out_data_32; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_33 = proc_6_io_pipe_phv_out_data_33; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_34 = proc_6_io_pipe_phv_out_data_34; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_35 = proc_6_io_pipe_phv_out_data_35; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_36 = proc_6_io_pipe_phv_out_data_36; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_37 = proc_6_io_pipe_phv_out_data_37; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_38 = proc_6_io_pipe_phv_out_data_38; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_39 = proc_6_io_pipe_phv_out_data_39; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_40 = proc_6_io_pipe_phv_out_data_40; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_41 = proc_6_io_pipe_phv_out_data_41; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_42 = proc_6_io_pipe_phv_out_data_42; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_43 = proc_6_io_pipe_phv_out_data_43; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_44 = proc_6_io_pipe_phv_out_data_44; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_45 = proc_6_io_pipe_phv_out_data_45; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_46 = proc_6_io_pipe_phv_out_data_46; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_47 = proc_6_io_pipe_phv_out_data_47; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_48 = proc_6_io_pipe_phv_out_data_48; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_49 = proc_6_io_pipe_phv_out_data_49; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_50 = proc_6_io_pipe_phv_out_data_50; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_51 = proc_6_io_pipe_phv_out_data_51; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_52 = proc_6_io_pipe_phv_out_data_52; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_53 = proc_6_io_pipe_phv_out_data_53; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_54 = proc_6_io_pipe_phv_out_data_54; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_55 = proc_6_io_pipe_phv_out_data_55; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_56 = proc_6_io_pipe_phv_out_data_56; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_57 = proc_6_io_pipe_phv_out_data_57; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_58 = proc_6_io_pipe_phv_out_data_58; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_59 = proc_6_io_pipe_phv_out_data_59; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_60 = proc_6_io_pipe_phv_out_data_60; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_61 = proc_6_io_pipe_phv_out_data_61; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_62 = proc_6_io_pipe_phv_out_data_62; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_63 = proc_6_io_pipe_phv_out_data_63; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_64 = proc_6_io_pipe_phv_out_data_64; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_65 = proc_6_io_pipe_phv_out_data_65; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_66 = proc_6_io_pipe_phv_out_data_66; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_67 = proc_6_io_pipe_phv_out_data_67; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_68 = proc_6_io_pipe_phv_out_data_68; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_69 = proc_6_io_pipe_phv_out_data_69; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_70 = proc_6_io_pipe_phv_out_data_70; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_71 = proc_6_io_pipe_phv_out_data_71; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_72 = proc_6_io_pipe_phv_out_data_72; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_73 = proc_6_io_pipe_phv_out_data_73; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_74 = proc_6_io_pipe_phv_out_data_74; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_75 = proc_6_io_pipe_phv_out_data_75; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_76 = proc_6_io_pipe_phv_out_data_76; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_77 = proc_6_io_pipe_phv_out_data_77; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_78 = proc_6_io_pipe_phv_out_data_78; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_79 = proc_6_io_pipe_phv_out_data_79; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_80 = proc_6_io_pipe_phv_out_data_80; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_81 = proc_6_io_pipe_phv_out_data_81; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_82 = proc_6_io_pipe_phv_out_data_82; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_83 = proc_6_io_pipe_phv_out_data_83; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_84 = proc_6_io_pipe_phv_out_data_84; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_85 = proc_6_io_pipe_phv_out_data_85; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_86 = proc_6_io_pipe_phv_out_data_86; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_87 = proc_6_io_pipe_phv_out_data_87; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_88 = proc_6_io_pipe_phv_out_data_88; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_89 = proc_6_io_pipe_phv_out_data_89; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_90 = proc_6_io_pipe_phv_out_data_90; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_91 = proc_6_io_pipe_phv_out_data_91; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_92 = proc_6_io_pipe_phv_out_data_92; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_93 = proc_6_io_pipe_phv_out_data_93; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_94 = proc_6_io_pipe_phv_out_data_94; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_95 = proc_6_io_pipe_phv_out_data_95; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_96 = proc_6_io_pipe_phv_out_data_96; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_97 = proc_6_io_pipe_phv_out_data_97; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_98 = proc_6_io_pipe_phv_out_data_98; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_99 = proc_6_io_pipe_phv_out_data_99; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_100 = proc_6_io_pipe_phv_out_data_100; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_101 = proc_6_io_pipe_phv_out_data_101; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_102 = proc_6_io_pipe_phv_out_data_102; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_103 = proc_6_io_pipe_phv_out_data_103; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_104 = proc_6_io_pipe_phv_out_data_104; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_105 = proc_6_io_pipe_phv_out_data_105; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_106 = proc_6_io_pipe_phv_out_data_106; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_107 = proc_6_io_pipe_phv_out_data_107; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_108 = proc_6_io_pipe_phv_out_data_108; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_109 = proc_6_io_pipe_phv_out_data_109; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_110 = proc_6_io_pipe_phv_out_data_110; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_111 = proc_6_io_pipe_phv_out_data_111; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_112 = proc_6_io_pipe_phv_out_data_112; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_113 = proc_6_io_pipe_phv_out_data_113; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_114 = proc_6_io_pipe_phv_out_data_114; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_115 = proc_6_io_pipe_phv_out_data_115; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_116 = proc_6_io_pipe_phv_out_data_116; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_117 = proc_6_io_pipe_phv_out_data_117; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_118 = proc_6_io_pipe_phv_out_data_118; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_119 = proc_6_io_pipe_phv_out_data_119; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_120 = proc_6_io_pipe_phv_out_data_120; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_121 = proc_6_io_pipe_phv_out_data_121; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_122 = proc_6_io_pipe_phv_out_data_122; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_123 = proc_6_io_pipe_phv_out_data_123; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_124 = proc_6_io_pipe_phv_out_data_124; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_125 = proc_6_io_pipe_phv_out_data_125; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_126 = proc_6_io_pipe_phv_out_data_126; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_127 = proc_6_io_pipe_phv_out_data_127; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_128 = proc_6_io_pipe_phv_out_data_128; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_129 = proc_6_io_pipe_phv_out_data_129; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_130 = proc_6_io_pipe_phv_out_data_130; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_131 = proc_6_io_pipe_phv_out_data_131; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_132 = proc_6_io_pipe_phv_out_data_132; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_133 = proc_6_io_pipe_phv_out_data_133; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_134 = proc_6_io_pipe_phv_out_data_134; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_135 = proc_6_io_pipe_phv_out_data_135; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_136 = proc_6_io_pipe_phv_out_data_136; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_137 = proc_6_io_pipe_phv_out_data_137; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_138 = proc_6_io_pipe_phv_out_data_138; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_139 = proc_6_io_pipe_phv_out_data_139; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_140 = proc_6_io_pipe_phv_out_data_140; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_141 = proc_6_io_pipe_phv_out_data_141; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_142 = proc_6_io_pipe_phv_out_data_142; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_143 = proc_6_io_pipe_phv_out_data_143; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_144 = proc_6_io_pipe_phv_out_data_144; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_145 = proc_6_io_pipe_phv_out_data_145; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_146 = proc_6_io_pipe_phv_out_data_146; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_147 = proc_6_io_pipe_phv_out_data_147; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_148 = proc_6_io_pipe_phv_out_data_148; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_149 = proc_6_io_pipe_phv_out_data_149; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_150 = proc_6_io_pipe_phv_out_data_150; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_151 = proc_6_io_pipe_phv_out_data_151; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_152 = proc_6_io_pipe_phv_out_data_152; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_153 = proc_6_io_pipe_phv_out_data_153; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_154 = proc_6_io_pipe_phv_out_data_154; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_155 = proc_6_io_pipe_phv_out_data_155; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_156 = proc_6_io_pipe_phv_out_data_156; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_157 = proc_6_io_pipe_phv_out_data_157; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_158 = proc_6_io_pipe_phv_out_data_158; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_data_159 = proc_6_io_pipe_phv_out_data_159; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_header_0 = proc_6_io_pipe_phv_out_header_0; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_header_1 = proc_6_io_pipe_phv_out_header_1; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_header_2 = proc_6_io_pipe_phv_out_header_2; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_header_3 = proc_6_io_pipe_phv_out_header_3; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_header_4 = proc_6_io_pipe_phv_out_header_4; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_header_5 = proc_6_io_pipe_phv_out_header_5; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_header_6 = proc_6_io_pipe_phv_out_header_6; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_header_7 = proc_6_io_pipe_phv_out_header_7; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_header_8 = proc_6_io_pipe_phv_out_header_8; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_header_9 = proc_6_io_pipe_phv_out_header_9; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_header_10 = proc_6_io_pipe_phv_out_header_10; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_header_11 = proc_6_io_pipe_phv_out_header_11; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_header_12 = proc_6_io_pipe_phv_out_header_12; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_header_13 = proc_6_io_pipe_phv_out_header_13; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_header_14 = proc_6_io_pipe_phv_out_header_14; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_header_15 = proc_6_io_pipe_phv_out_header_15; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_parse_current_state = proc_6_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_parse_current_offset = proc_6_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_parse_transition_field = proc_6_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_next_processor_id = proc_6_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_next_config_id = proc_6_io_pipe_phv_out_next_config_id; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_valid = proc_6_io_pipe_phv_out_valid; // @[ipsa.scala 82:32]
  assign trans_6_io_pipe_phv_in_last = proc_6_io_pipe_phv_out_last; // @[ipsa.scala 82:32]
  assign trans_6_io_next_proc_exist = 1'h1; // @[ipsa.scala 80:48]
  assign trans_7_clock = clock;
  assign trans_7_io_pipe_phv_in_data_0 = proc_7_io_pipe_phv_out_data_0; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_1 = proc_7_io_pipe_phv_out_data_1; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_2 = proc_7_io_pipe_phv_out_data_2; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_3 = proc_7_io_pipe_phv_out_data_3; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_4 = proc_7_io_pipe_phv_out_data_4; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_5 = proc_7_io_pipe_phv_out_data_5; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_6 = proc_7_io_pipe_phv_out_data_6; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_7 = proc_7_io_pipe_phv_out_data_7; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_8 = proc_7_io_pipe_phv_out_data_8; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_9 = proc_7_io_pipe_phv_out_data_9; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_10 = proc_7_io_pipe_phv_out_data_10; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_11 = proc_7_io_pipe_phv_out_data_11; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_12 = proc_7_io_pipe_phv_out_data_12; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_13 = proc_7_io_pipe_phv_out_data_13; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_14 = proc_7_io_pipe_phv_out_data_14; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_15 = proc_7_io_pipe_phv_out_data_15; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_16 = proc_7_io_pipe_phv_out_data_16; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_17 = proc_7_io_pipe_phv_out_data_17; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_18 = proc_7_io_pipe_phv_out_data_18; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_19 = proc_7_io_pipe_phv_out_data_19; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_20 = proc_7_io_pipe_phv_out_data_20; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_21 = proc_7_io_pipe_phv_out_data_21; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_22 = proc_7_io_pipe_phv_out_data_22; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_23 = proc_7_io_pipe_phv_out_data_23; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_24 = proc_7_io_pipe_phv_out_data_24; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_25 = proc_7_io_pipe_phv_out_data_25; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_26 = proc_7_io_pipe_phv_out_data_26; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_27 = proc_7_io_pipe_phv_out_data_27; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_28 = proc_7_io_pipe_phv_out_data_28; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_29 = proc_7_io_pipe_phv_out_data_29; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_30 = proc_7_io_pipe_phv_out_data_30; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_31 = proc_7_io_pipe_phv_out_data_31; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_32 = proc_7_io_pipe_phv_out_data_32; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_33 = proc_7_io_pipe_phv_out_data_33; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_34 = proc_7_io_pipe_phv_out_data_34; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_35 = proc_7_io_pipe_phv_out_data_35; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_36 = proc_7_io_pipe_phv_out_data_36; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_37 = proc_7_io_pipe_phv_out_data_37; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_38 = proc_7_io_pipe_phv_out_data_38; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_39 = proc_7_io_pipe_phv_out_data_39; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_40 = proc_7_io_pipe_phv_out_data_40; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_41 = proc_7_io_pipe_phv_out_data_41; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_42 = proc_7_io_pipe_phv_out_data_42; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_43 = proc_7_io_pipe_phv_out_data_43; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_44 = proc_7_io_pipe_phv_out_data_44; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_45 = proc_7_io_pipe_phv_out_data_45; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_46 = proc_7_io_pipe_phv_out_data_46; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_47 = proc_7_io_pipe_phv_out_data_47; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_48 = proc_7_io_pipe_phv_out_data_48; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_49 = proc_7_io_pipe_phv_out_data_49; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_50 = proc_7_io_pipe_phv_out_data_50; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_51 = proc_7_io_pipe_phv_out_data_51; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_52 = proc_7_io_pipe_phv_out_data_52; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_53 = proc_7_io_pipe_phv_out_data_53; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_54 = proc_7_io_pipe_phv_out_data_54; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_55 = proc_7_io_pipe_phv_out_data_55; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_56 = proc_7_io_pipe_phv_out_data_56; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_57 = proc_7_io_pipe_phv_out_data_57; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_58 = proc_7_io_pipe_phv_out_data_58; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_59 = proc_7_io_pipe_phv_out_data_59; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_60 = proc_7_io_pipe_phv_out_data_60; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_61 = proc_7_io_pipe_phv_out_data_61; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_62 = proc_7_io_pipe_phv_out_data_62; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_63 = proc_7_io_pipe_phv_out_data_63; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_64 = proc_7_io_pipe_phv_out_data_64; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_65 = proc_7_io_pipe_phv_out_data_65; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_66 = proc_7_io_pipe_phv_out_data_66; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_67 = proc_7_io_pipe_phv_out_data_67; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_68 = proc_7_io_pipe_phv_out_data_68; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_69 = proc_7_io_pipe_phv_out_data_69; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_70 = proc_7_io_pipe_phv_out_data_70; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_71 = proc_7_io_pipe_phv_out_data_71; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_72 = proc_7_io_pipe_phv_out_data_72; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_73 = proc_7_io_pipe_phv_out_data_73; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_74 = proc_7_io_pipe_phv_out_data_74; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_75 = proc_7_io_pipe_phv_out_data_75; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_76 = proc_7_io_pipe_phv_out_data_76; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_77 = proc_7_io_pipe_phv_out_data_77; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_78 = proc_7_io_pipe_phv_out_data_78; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_79 = proc_7_io_pipe_phv_out_data_79; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_80 = proc_7_io_pipe_phv_out_data_80; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_81 = proc_7_io_pipe_phv_out_data_81; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_82 = proc_7_io_pipe_phv_out_data_82; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_83 = proc_7_io_pipe_phv_out_data_83; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_84 = proc_7_io_pipe_phv_out_data_84; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_85 = proc_7_io_pipe_phv_out_data_85; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_86 = proc_7_io_pipe_phv_out_data_86; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_87 = proc_7_io_pipe_phv_out_data_87; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_88 = proc_7_io_pipe_phv_out_data_88; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_89 = proc_7_io_pipe_phv_out_data_89; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_90 = proc_7_io_pipe_phv_out_data_90; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_91 = proc_7_io_pipe_phv_out_data_91; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_92 = proc_7_io_pipe_phv_out_data_92; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_93 = proc_7_io_pipe_phv_out_data_93; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_94 = proc_7_io_pipe_phv_out_data_94; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_95 = proc_7_io_pipe_phv_out_data_95; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_96 = proc_7_io_pipe_phv_out_data_96; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_97 = proc_7_io_pipe_phv_out_data_97; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_98 = proc_7_io_pipe_phv_out_data_98; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_99 = proc_7_io_pipe_phv_out_data_99; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_100 = proc_7_io_pipe_phv_out_data_100; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_101 = proc_7_io_pipe_phv_out_data_101; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_102 = proc_7_io_pipe_phv_out_data_102; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_103 = proc_7_io_pipe_phv_out_data_103; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_104 = proc_7_io_pipe_phv_out_data_104; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_105 = proc_7_io_pipe_phv_out_data_105; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_106 = proc_7_io_pipe_phv_out_data_106; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_107 = proc_7_io_pipe_phv_out_data_107; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_108 = proc_7_io_pipe_phv_out_data_108; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_109 = proc_7_io_pipe_phv_out_data_109; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_110 = proc_7_io_pipe_phv_out_data_110; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_111 = proc_7_io_pipe_phv_out_data_111; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_112 = proc_7_io_pipe_phv_out_data_112; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_113 = proc_7_io_pipe_phv_out_data_113; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_114 = proc_7_io_pipe_phv_out_data_114; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_115 = proc_7_io_pipe_phv_out_data_115; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_116 = proc_7_io_pipe_phv_out_data_116; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_117 = proc_7_io_pipe_phv_out_data_117; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_118 = proc_7_io_pipe_phv_out_data_118; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_119 = proc_7_io_pipe_phv_out_data_119; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_120 = proc_7_io_pipe_phv_out_data_120; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_121 = proc_7_io_pipe_phv_out_data_121; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_122 = proc_7_io_pipe_phv_out_data_122; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_123 = proc_7_io_pipe_phv_out_data_123; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_124 = proc_7_io_pipe_phv_out_data_124; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_125 = proc_7_io_pipe_phv_out_data_125; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_126 = proc_7_io_pipe_phv_out_data_126; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_127 = proc_7_io_pipe_phv_out_data_127; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_128 = proc_7_io_pipe_phv_out_data_128; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_129 = proc_7_io_pipe_phv_out_data_129; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_130 = proc_7_io_pipe_phv_out_data_130; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_131 = proc_7_io_pipe_phv_out_data_131; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_132 = proc_7_io_pipe_phv_out_data_132; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_133 = proc_7_io_pipe_phv_out_data_133; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_134 = proc_7_io_pipe_phv_out_data_134; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_135 = proc_7_io_pipe_phv_out_data_135; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_136 = proc_7_io_pipe_phv_out_data_136; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_137 = proc_7_io_pipe_phv_out_data_137; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_138 = proc_7_io_pipe_phv_out_data_138; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_139 = proc_7_io_pipe_phv_out_data_139; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_140 = proc_7_io_pipe_phv_out_data_140; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_141 = proc_7_io_pipe_phv_out_data_141; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_142 = proc_7_io_pipe_phv_out_data_142; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_143 = proc_7_io_pipe_phv_out_data_143; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_144 = proc_7_io_pipe_phv_out_data_144; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_145 = proc_7_io_pipe_phv_out_data_145; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_146 = proc_7_io_pipe_phv_out_data_146; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_147 = proc_7_io_pipe_phv_out_data_147; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_148 = proc_7_io_pipe_phv_out_data_148; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_149 = proc_7_io_pipe_phv_out_data_149; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_150 = proc_7_io_pipe_phv_out_data_150; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_151 = proc_7_io_pipe_phv_out_data_151; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_152 = proc_7_io_pipe_phv_out_data_152; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_153 = proc_7_io_pipe_phv_out_data_153; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_154 = proc_7_io_pipe_phv_out_data_154; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_155 = proc_7_io_pipe_phv_out_data_155; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_156 = proc_7_io_pipe_phv_out_data_156; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_157 = proc_7_io_pipe_phv_out_data_157; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_158 = proc_7_io_pipe_phv_out_data_158; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_data_159 = proc_7_io_pipe_phv_out_data_159; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_header_0 = proc_7_io_pipe_phv_out_header_0; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_header_1 = proc_7_io_pipe_phv_out_header_1; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_header_2 = proc_7_io_pipe_phv_out_header_2; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_header_3 = proc_7_io_pipe_phv_out_header_3; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_header_4 = proc_7_io_pipe_phv_out_header_4; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_header_5 = proc_7_io_pipe_phv_out_header_5; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_header_6 = proc_7_io_pipe_phv_out_header_6; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_header_7 = proc_7_io_pipe_phv_out_header_7; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_header_8 = proc_7_io_pipe_phv_out_header_8; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_header_9 = proc_7_io_pipe_phv_out_header_9; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_header_10 = proc_7_io_pipe_phv_out_header_10; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_header_11 = proc_7_io_pipe_phv_out_header_11; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_header_12 = proc_7_io_pipe_phv_out_header_12; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_header_13 = proc_7_io_pipe_phv_out_header_13; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_header_14 = proc_7_io_pipe_phv_out_header_14; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_header_15 = proc_7_io_pipe_phv_out_header_15; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_parse_current_state = proc_7_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_parse_current_offset = proc_7_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_parse_transition_field = proc_7_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_next_processor_id = proc_7_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_next_config_id = proc_7_io_pipe_phv_out_next_config_id; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_valid = proc_7_io_pipe_phv_out_valid; // @[ipsa.scala 82:32]
  assign trans_7_io_pipe_phv_in_last = proc_7_io_pipe_phv_out_last; // @[ipsa.scala 82:32]
  assign trans_7_io_next_proc_exist = 1'h1; // @[ipsa.scala 80:48]
  assign trans_8_clock = clock;
  assign trans_8_io_pipe_phv_in_data_0 = proc_8_io_pipe_phv_out_data_0; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_1 = proc_8_io_pipe_phv_out_data_1; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_2 = proc_8_io_pipe_phv_out_data_2; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_3 = proc_8_io_pipe_phv_out_data_3; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_4 = proc_8_io_pipe_phv_out_data_4; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_5 = proc_8_io_pipe_phv_out_data_5; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_6 = proc_8_io_pipe_phv_out_data_6; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_7 = proc_8_io_pipe_phv_out_data_7; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_8 = proc_8_io_pipe_phv_out_data_8; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_9 = proc_8_io_pipe_phv_out_data_9; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_10 = proc_8_io_pipe_phv_out_data_10; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_11 = proc_8_io_pipe_phv_out_data_11; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_12 = proc_8_io_pipe_phv_out_data_12; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_13 = proc_8_io_pipe_phv_out_data_13; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_14 = proc_8_io_pipe_phv_out_data_14; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_15 = proc_8_io_pipe_phv_out_data_15; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_16 = proc_8_io_pipe_phv_out_data_16; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_17 = proc_8_io_pipe_phv_out_data_17; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_18 = proc_8_io_pipe_phv_out_data_18; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_19 = proc_8_io_pipe_phv_out_data_19; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_20 = proc_8_io_pipe_phv_out_data_20; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_21 = proc_8_io_pipe_phv_out_data_21; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_22 = proc_8_io_pipe_phv_out_data_22; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_23 = proc_8_io_pipe_phv_out_data_23; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_24 = proc_8_io_pipe_phv_out_data_24; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_25 = proc_8_io_pipe_phv_out_data_25; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_26 = proc_8_io_pipe_phv_out_data_26; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_27 = proc_8_io_pipe_phv_out_data_27; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_28 = proc_8_io_pipe_phv_out_data_28; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_29 = proc_8_io_pipe_phv_out_data_29; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_30 = proc_8_io_pipe_phv_out_data_30; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_31 = proc_8_io_pipe_phv_out_data_31; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_32 = proc_8_io_pipe_phv_out_data_32; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_33 = proc_8_io_pipe_phv_out_data_33; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_34 = proc_8_io_pipe_phv_out_data_34; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_35 = proc_8_io_pipe_phv_out_data_35; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_36 = proc_8_io_pipe_phv_out_data_36; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_37 = proc_8_io_pipe_phv_out_data_37; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_38 = proc_8_io_pipe_phv_out_data_38; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_39 = proc_8_io_pipe_phv_out_data_39; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_40 = proc_8_io_pipe_phv_out_data_40; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_41 = proc_8_io_pipe_phv_out_data_41; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_42 = proc_8_io_pipe_phv_out_data_42; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_43 = proc_8_io_pipe_phv_out_data_43; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_44 = proc_8_io_pipe_phv_out_data_44; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_45 = proc_8_io_pipe_phv_out_data_45; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_46 = proc_8_io_pipe_phv_out_data_46; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_47 = proc_8_io_pipe_phv_out_data_47; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_48 = proc_8_io_pipe_phv_out_data_48; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_49 = proc_8_io_pipe_phv_out_data_49; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_50 = proc_8_io_pipe_phv_out_data_50; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_51 = proc_8_io_pipe_phv_out_data_51; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_52 = proc_8_io_pipe_phv_out_data_52; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_53 = proc_8_io_pipe_phv_out_data_53; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_54 = proc_8_io_pipe_phv_out_data_54; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_55 = proc_8_io_pipe_phv_out_data_55; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_56 = proc_8_io_pipe_phv_out_data_56; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_57 = proc_8_io_pipe_phv_out_data_57; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_58 = proc_8_io_pipe_phv_out_data_58; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_59 = proc_8_io_pipe_phv_out_data_59; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_60 = proc_8_io_pipe_phv_out_data_60; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_61 = proc_8_io_pipe_phv_out_data_61; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_62 = proc_8_io_pipe_phv_out_data_62; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_63 = proc_8_io_pipe_phv_out_data_63; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_64 = proc_8_io_pipe_phv_out_data_64; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_65 = proc_8_io_pipe_phv_out_data_65; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_66 = proc_8_io_pipe_phv_out_data_66; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_67 = proc_8_io_pipe_phv_out_data_67; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_68 = proc_8_io_pipe_phv_out_data_68; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_69 = proc_8_io_pipe_phv_out_data_69; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_70 = proc_8_io_pipe_phv_out_data_70; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_71 = proc_8_io_pipe_phv_out_data_71; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_72 = proc_8_io_pipe_phv_out_data_72; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_73 = proc_8_io_pipe_phv_out_data_73; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_74 = proc_8_io_pipe_phv_out_data_74; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_75 = proc_8_io_pipe_phv_out_data_75; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_76 = proc_8_io_pipe_phv_out_data_76; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_77 = proc_8_io_pipe_phv_out_data_77; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_78 = proc_8_io_pipe_phv_out_data_78; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_79 = proc_8_io_pipe_phv_out_data_79; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_80 = proc_8_io_pipe_phv_out_data_80; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_81 = proc_8_io_pipe_phv_out_data_81; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_82 = proc_8_io_pipe_phv_out_data_82; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_83 = proc_8_io_pipe_phv_out_data_83; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_84 = proc_8_io_pipe_phv_out_data_84; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_85 = proc_8_io_pipe_phv_out_data_85; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_86 = proc_8_io_pipe_phv_out_data_86; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_87 = proc_8_io_pipe_phv_out_data_87; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_88 = proc_8_io_pipe_phv_out_data_88; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_89 = proc_8_io_pipe_phv_out_data_89; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_90 = proc_8_io_pipe_phv_out_data_90; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_91 = proc_8_io_pipe_phv_out_data_91; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_92 = proc_8_io_pipe_phv_out_data_92; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_93 = proc_8_io_pipe_phv_out_data_93; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_94 = proc_8_io_pipe_phv_out_data_94; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_95 = proc_8_io_pipe_phv_out_data_95; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_96 = proc_8_io_pipe_phv_out_data_96; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_97 = proc_8_io_pipe_phv_out_data_97; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_98 = proc_8_io_pipe_phv_out_data_98; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_99 = proc_8_io_pipe_phv_out_data_99; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_100 = proc_8_io_pipe_phv_out_data_100; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_101 = proc_8_io_pipe_phv_out_data_101; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_102 = proc_8_io_pipe_phv_out_data_102; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_103 = proc_8_io_pipe_phv_out_data_103; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_104 = proc_8_io_pipe_phv_out_data_104; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_105 = proc_8_io_pipe_phv_out_data_105; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_106 = proc_8_io_pipe_phv_out_data_106; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_107 = proc_8_io_pipe_phv_out_data_107; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_108 = proc_8_io_pipe_phv_out_data_108; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_109 = proc_8_io_pipe_phv_out_data_109; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_110 = proc_8_io_pipe_phv_out_data_110; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_111 = proc_8_io_pipe_phv_out_data_111; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_112 = proc_8_io_pipe_phv_out_data_112; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_113 = proc_8_io_pipe_phv_out_data_113; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_114 = proc_8_io_pipe_phv_out_data_114; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_115 = proc_8_io_pipe_phv_out_data_115; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_116 = proc_8_io_pipe_phv_out_data_116; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_117 = proc_8_io_pipe_phv_out_data_117; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_118 = proc_8_io_pipe_phv_out_data_118; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_119 = proc_8_io_pipe_phv_out_data_119; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_120 = proc_8_io_pipe_phv_out_data_120; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_121 = proc_8_io_pipe_phv_out_data_121; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_122 = proc_8_io_pipe_phv_out_data_122; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_123 = proc_8_io_pipe_phv_out_data_123; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_124 = proc_8_io_pipe_phv_out_data_124; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_125 = proc_8_io_pipe_phv_out_data_125; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_126 = proc_8_io_pipe_phv_out_data_126; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_127 = proc_8_io_pipe_phv_out_data_127; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_128 = proc_8_io_pipe_phv_out_data_128; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_129 = proc_8_io_pipe_phv_out_data_129; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_130 = proc_8_io_pipe_phv_out_data_130; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_131 = proc_8_io_pipe_phv_out_data_131; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_132 = proc_8_io_pipe_phv_out_data_132; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_133 = proc_8_io_pipe_phv_out_data_133; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_134 = proc_8_io_pipe_phv_out_data_134; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_135 = proc_8_io_pipe_phv_out_data_135; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_136 = proc_8_io_pipe_phv_out_data_136; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_137 = proc_8_io_pipe_phv_out_data_137; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_138 = proc_8_io_pipe_phv_out_data_138; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_139 = proc_8_io_pipe_phv_out_data_139; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_140 = proc_8_io_pipe_phv_out_data_140; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_141 = proc_8_io_pipe_phv_out_data_141; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_142 = proc_8_io_pipe_phv_out_data_142; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_143 = proc_8_io_pipe_phv_out_data_143; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_144 = proc_8_io_pipe_phv_out_data_144; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_145 = proc_8_io_pipe_phv_out_data_145; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_146 = proc_8_io_pipe_phv_out_data_146; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_147 = proc_8_io_pipe_phv_out_data_147; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_148 = proc_8_io_pipe_phv_out_data_148; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_149 = proc_8_io_pipe_phv_out_data_149; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_150 = proc_8_io_pipe_phv_out_data_150; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_151 = proc_8_io_pipe_phv_out_data_151; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_152 = proc_8_io_pipe_phv_out_data_152; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_153 = proc_8_io_pipe_phv_out_data_153; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_154 = proc_8_io_pipe_phv_out_data_154; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_155 = proc_8_io_pipe_phv_out_data_155; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_156 = proc_8_io_pipe_phv_out_data_156; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_157 = proc_8_io_pipe_phv_out_data_157; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_158 = proc_8_io_pipe_phv_out_data_158; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_data_159 = proc_8_io_pipe_phv_out_data_159; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_header_0 = proc_8_io_pipe_phv_out_header_0; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_header_1 = proc_8_io_pipe_phv_out_header_1; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_header_2 = proc_8_io_pipe_phv_out_header_2; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_header_3 = proc_8_io_pipe_phv_out_header_3; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_header_4 = proc_8_io_pipe_phv_out_header_4; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_header_5 = proc_8_io_pipe_phv_out_header_5; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_header_6 = proc_8_io_pipe_phv_out_header_6; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_header_7 = proc_8_io_pipe_phv_out_header_7; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_header_8 = proc_8_io_pipe_phv_out_header_8; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_header_9 = proc_8_io_pipe_phv_out_header_9; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_header_10 = proc_8_io_pipe_phv_out_header_10; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_header_11 = proc_8_io_pipe_phv_out_header_11; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_header_12 = proc_8_io_pipe_phv_out_header_12; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_header_13 = proc_8_io_pipe_phv_out_header_13; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_header_14 = proc_8_io_pipe_phv_out_header_14; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_header_15 = proc_8_io_pipe_phv_out_header_15; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_parse_current_state = proc_8_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_parse_current_offset = proc_8_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_parse_transition_field = proc_8_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_next_processor_id = proc_8_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_next_config_id = proc_8_io_pipe_phv_out_next_config_id; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_valid = proc_8_io_pipe_phv_out_valid; // @[ipsa.scala 82:32]
  assign trans_8_io_pipe_phv_in_last = proc_8_io_pipe_phv_out_last; // @[ipsa.scala 82:32]
  assign trans_8_io_next_proc_exist = 1'h1; // @[ipsa.scala 80:48]
  assign trans_9_clock = clock;
  assign trans_9_io_pipe_phv_in_data_0 = proc_9_io_pipe_phv_out_data_0; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_1 = proc_9_io_pipe_phv_out_data_1; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_2 = proc_9_io_pipe_phv_out_data_2; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_3 = proc_9_io_pipe_phv_out_data_3; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_4 = proc_9_io_pipe_phv_out_data_4; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_5 = proc_9_io_pipe_phv_out_data_5; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_6 = proc_9_io_pipe_phv_out_data_6; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_7 = proc_9_io_pipe_phv_out_data_7; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_8 = proc_9_io_pipe_phv_out_data_8; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_9 = proc_9_io_pipe_phv_out_data_9; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_10 = proc_9_io_pipe_phv_out_data_10; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_11 = proc_9_io_pipe_phv_out_data_11; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_12 = proc_9_io_pipe_phv_out_data_12; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_13 = proc_9_io_pipe_phv_out_data_13; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_14 = proc_9_io_pipe_phv_out_data_14; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_15 = proc_9_io_pipe_phv_out_data_15; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_16 = proc_9_io_pipe_phv_out_data_16; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_17 = proc_9_io_pipe_phv_out_data_17; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_18 = proc_9_io_pipe_phv_out_data_18; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_19 = proc_9_io_pipe_phv_out_data_19; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_20 = proc_9_io_pipe_phv_out_data_20; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_21 = proc_9_io_pipe_phv_out_data_21; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_22 = proc_9_io_pipe_phv_out_data_22; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_23 = proc_9_io_pipe_phv_out_data_23; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_24 = proc_9_io_pipe_phv_out_data_24; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_25 = proc_9_io_pipe_phv_out_data_25; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_26 = proc_9_io_pipe_phv_out_data_26; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_27 = proc_9_io_pipe_phv_out_data_27; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_28 = proc_9_io_pipe_phv_out_data_28; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_29 = proc_9_io_pipe_phv_out_data_29; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_30 = proc_9_io_pipe_phv_out_data_30; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_31 = proc_9_io_pipe_phv_out_data_31; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_32 = proc_9_io_pipe_phv_out_data_32; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_33 = proc_9_io_pipe_phv_out_data_33; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_34 = proc_9_io_pipe_phv_out_data_34; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_35 = proc_9_io_pipe_phv_out_data_35; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_36 = proc_9_io_pipe_phv_out_data_36; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_37 = proc_9_io_pipe_phv_out_data_37; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_38 = proc_9_io_pipe_phv_out_data_38; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_39 = proc_9_io_pipe_phv_out_data_39; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_40 = proc_9_io_pipe_phv_out_data_40; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_41 = proc_9_io_pipe_phv_out_data_41; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_42 = proc_9_io_pipe_phv_out_data_42; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_43 = proc_9_io_pipe_phv_out_data_43; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_44 = proc_9_io_pipe_phv_out_data_44; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_45 = proc_9_io_pipe_phv_out_data_45; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_46 = proc_9_io_pipe_phv_out_data_46; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_47 = proc_9_io_pipe_phv_out_data_47; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_48 = proc_9_io_pipe_phv_out_data_48; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_49 = proc_9_io_pipe_phv_out_data_49; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_50 = proc_9_io_pipe_phv_out_data_50; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_51 = proc_9_io_pipe_phv_out_data_51; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_52 = proc_9_io_pipe_phv_out_data_52; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_53 = proc_9_io_pipe_phv_out_data_53; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_54 = proc_9_io_pipe_phv_out_data_54; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_55 = proc_9_io_pipe_phv_out_data_55; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_56 = proc_9_io_pipe_phv_out_data_56; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_57 = proc_9_io_pipe_phv_out_data_57; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_58 = proc_9_io_pipe_phv_out_data_58; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_59 = proc_9_io_pipe_phv_out_data_59; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_60 = proc_9_io_pipe_phv_out_data_60; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_61 = proc_9_io_pipe_phv_out_data_61; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_62 = proc_9_io_pipe_phv_out_data_62; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_63 = proc_9_io_pipe_phv_out_data_63; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_64 = proc_9_io_pipe_phv_out_data_64; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_65 = proc_9_io_pipe_phv_out_data_65; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_66 = proc_9_io_pipe_phv_out_data_66; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_67 = proc_9_io_pipe_phv_out_data_67; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_68 = proc_9_io_pipe_phv_out_data_68; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_69 = proc_9_io_pipe_phv_out_data_69; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_70 = proc_9_io_pipe_phv_out_data_70; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_71 = proc_9_io_pipe_phv_out_data_71; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_72 = proc_9_io_pipe_phv_out_data_72; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_73 = proc_9_io_pipe_phv_out_data_73; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_74 = proc_9_io_pipe_phv_out_data_74; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_75 = proc_9_io_pipe_phv_out_data_75; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_76 = proc_9_io_pipe_phv_out_data_76; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_77 = proc_9_io_pipe_phv_out_data_77; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_78 = proc_9_io_pipe_phv_out_data_78; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_79 = proc_9_io_pipe_phv_out_data_79; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_80 = proc_9_io_pipe_phv_out_data_80; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_81 = proc_9_io_pipe_phv_out_data_81; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_82 = proc_9_io_pipe_phv_out_data_82; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_83 = proc_9_io_pipe_phv_out_data_83; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_84 = proc_9_io_pipe_phv_out_data_84; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_85 = proc_9_io_pipe_phv_out_data_85; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_86 = proc_9_io_pipe_phv_out_data_86; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_87 = proc_9_io_pipe_phv_out_data_87; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_88 = proc_9_io_pipe_phv_out_data_88; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_89 = proc_9_io_pipe_phv_out_data_89; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_90 = proc_9_io_pipe_phv_out_data_90; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_91 = proc_9_io_pipe_phv_out_data_91; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_92 = proc_9_io_pipe_phv_out_data_92; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_93 = proc_9_io_pipe_phv_out_data_93; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_94 = proc_9_io_pipe_phv_out_data_94; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_95 = proc_9_io_pipe_phv_out_data_95; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_96 = proc_9_io_pipe_phv_out_data_96; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_97 = proc_9_io_pipe_phv_out_data_97; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_98 = proc_9_io_pipe_phv_out_data_98; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_99 = proc_9_io_pipe_phv_out_data_99; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_100 = proc_9_io_pipe_phv_out_data_100; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_101 = proc_9_io_pipe_phv_out_data_101; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_102 = proc_9_io_pipe_phv_out_data_102; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_103 = proc_9_io_pipe_phv_out_data_103; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_104 = proc_9_io_pipe_phv_out_data_104; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_105 = proc_9_io_pipe_phv_out_data_105; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_106 = proc_9_io_pipe_phv_out_data_106; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_107 = proc_9_io_pipe_phv_out_data_107; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_108 = proc_9_io_pipe_phv_out_data_108; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_109 = proc_9_io_pipe_phv_out_data_109; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_110 = proc_9_io_pipe_phv_out_data_110; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_111 = proc_9_io_pipe_phv_out_data_111; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_112 = proc_9_io_pipe_phv_out_data_112; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_113 = proc_9_io_pipe_phv_out_data_113; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_114 = proc_9_io_pipe_phv_out_data_114; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_115 = proc_9_io_pipe_phv_out_data_115; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_116 = proc_9_io_pipe_phv_out_data_116; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_117 = proc_9_io_pipe_phv_out_data_117; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_118 = proc_9_io_pipe_phv_out_data_118; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_119 = proc_9_io_pipe_phv_out_data_119; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_120 = proc_9_io_pipe_phv_out_data_120; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_121 = proc_9_io_pipe_phv_out_data_121; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_122 = proc_9_io_pipe_phv_out_data_122; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_123 = proc_9_io_pipe_phv_out_data_123; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_124 = proc_9_io_pipe_phv_out_data_124; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_125 = proc_9_io_pipe_phv_out_data_125; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_126 = proc_9_io_pipe_phv_out_data_126; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_127 = proc_9_io_pipe_phv_out_data_127; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_128 = proc_9_io_pipe_phv_out_data_128; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_129 = proc_9_io_pipe_phv_out_data_129; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_130 = proc_9_io_pipe_phv_out_data_130; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_131 = proc_9_io_pipe_phv_out_data_131; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_132 = proc_9_io_pipe_phv_out_data_132; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_133 = proc_9_io_pipe_phv_out_data_133; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_134 = proc_9_io_pipe_phv_out_data_134; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_135 = proc_9_io_pipe_phv_out_data_135; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_136 = proc_9_io_pipe_phv_out_data_136; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_137 = proc_9_io_pipe_phv_out_data_137; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_138 = proc_9_io_pipe_phv_out_data_138; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_139 = proc_9_io_pipe_phv_out_data_139; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_140 = proc_9_io_pipe_phv_out_data_140; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_141 = proc_9_io_pipe_phv_out_data_141; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_142 = proc_9_io_pipe_phv_out_data_142; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_143 = proc_9_io_pipe_phv_out_data_143; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_144 = proc_9_io_pipe_phv_out_data_144; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_145 = proc_9_io_pipe_phv_out_data_145; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_146 = proc_9_io_pipe_phv_out_data_146; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_147 = proc_9_io_pipe_phv_out_data_147; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_148 = proc_9_io_pipe_phv_out_data_148; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_149 = proc_9_io_pipe_phv_out_data_149; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_150 = proc_9_io_pipe_phv_out_data_150; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_151 = proc_9_io_pipe_phv_out_data_151; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_152 = proc_9_io_pipe_phv_out_data_152; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_153 = proc_9_io_pipe_phv_out_data_153; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_154 = proc_9_io_pipe_phv_out_data_154; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_155 = proc_9_io_pipe_phv_out_data_155; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_156 = proc_9_io_pipe_phv_out_data_156; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_157 = proc_9_io_pipe_phv_out_data_157; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_158 = proc_9_io_pipe_phv_out_data_158; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_data_159 = proc_9_io_pipe_phv_out_data_159; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_header_0 = proc_9_io_pipe_phv_out_header_0; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_header_1 = proc_9_io_pipe_phv_out_header_1; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_header_2 = proc_9_io_pipe_phv_out_header_2; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_header_3 = proc_9_io_pipe_phv_out_header_3; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_header_4 = proc_9_io_pipe_phv_out_header_4; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_header_5 = proc_9_io_pipe_phv_out_header_5; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_header_6 = proc_9_io_pipe_phv_out_header_6; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_header_7 = proc_9_io_pipe_phv_out_header_7; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_header_8 = proc_9_io_pipe_phv_out_header_8; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_header_9 = proc_9_io_pipe_phv_out_header_9; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_header_10 = proc_9_io_pipe_phv_out_header_10; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_header_11 = proc_9_io_pipe_phv_out_header_11; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_header_12 = proc_9_io_pipe_phv_out_header_12; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_header_13 = proc_9_io_pipe_phv_out_header_13; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_header_14 = proc_9_io_pipe_phv_out_header_14; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_header_15 = proc_9_io_pipe_phv_out_header_15; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_parse_current_state = proc_9_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_parse_current_offset = proc_9_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_parse_transition_field = proc_9_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_next_processor_id = proc_9_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_next_config_id = proc_9_io_pipe_phv_out_next_config_id; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_valid = proc_9_io_pipe_phv_out_valid; // @[ipsa.scala 82:32]
  assign trans_9_io_pipe_phv_in_last = proc_9_io_pipe_phv_out_last; // @[ipsa.scala 82:32]
  assign trans_9_io_next_proc_exist = 1'h1; // @[ipsa.scala 80:48]
  assign trans_10_clock = clock;
  assign trans_10_io_pipe_phv_in_data_0 = proc_10_io_pipe_phv_out_data_0; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_1 = proc_10_io_pipe_phv_out_data_1; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_2 = proc_10_io_pipe_phv_out_data_2; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_3 = proc_10_io_pipe_phv_out_data_3; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_4 = proc_10_io_pipe_phv_out_data_4; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_5 = proc_10_io_pipe_phv_out_data_5; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_6 = proc_10_io_pipe_phv_out_data_6; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_7 = proc_10_io_pipe_phv_out_data_7; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_8 = proc_10_io_pipe_phv_out_data_8; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_9 = proc_10_io_pipe_phv_out_data_9; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_10 = proc_10_io_pipe_phv_out_data_10; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_11 = proc_10_io_pipe_phv_out_data_11; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_12 = proc_10_io_pipe_phv_out_data_12; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_13 = proc_10_io_pipe_phv_out_data_13; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_14 = proc_10_io_pipe_phv_out_data_14; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_15 = proc_10_io_pipe_phv_out_data_15; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_16 = proc_10_io_pipe_phv_out_data_16; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_17 = proc_10_io_pipe_phv_out_data_17; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_18 = proc_10_io_pipe_phv_out_data_18; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_19 = proc_10_io_pipe_phv_out_data_19; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_20 = proc_10_io_pipe_phv_out_data_20; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_21 = proc_10_io_pipe_phv_out_data_21; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_22 = proc_10_io_pipe_phv_out_data_22; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_23 = proc_10_io_pipe_phv_out_data_23; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_24 = proc_10_io_pipe_phv_out_data_24; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_25 = proc_10_io_pipe_phv_out_data_25; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_26 = proc_10_io_pipe_phv_out_data_26; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_27 = proc_10_io_pipe_phv_out_data_27; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_28 = proc_10_io_pipe_phv_out_data_28; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_29 = proc_10_io_pipe_phv_out_data_29; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_30 = proc_10_io_pipe_phv_out_data_30; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_31 = proc_10_io_pipe_phv_out_data_31; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_32 = proc_10_io_pipe_phv_out_data_32; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_33 = proc_10_io_pipe_phv_out_data_33; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_34 = proc_10_io_pipe_phv_out_data_34; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_35 = proc_10_io_pipe_phv_out_data_35; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_36 = proc_10_io_pipe_phv_out_data_36; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_37 = proc_10_io_pipe_phv_out_data_37; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_38 = proc_10_io_pipe_phv_out_data_38; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_39 = proc_10_io_pipe_phv_out_data_39; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_40 = proc_10_io_pipe_phv_out_data_40; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_41 = proc_10_io_pipe_phv_out_data_41; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_42 = proc_10_io_pipe_phv_out_data_42; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_43 = proc_10_io_pipe_phv_out_data_43; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_44 = proc_10_io_pipe_phv_out_data_44; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_45 = proc_10_io_pipe_phv_out_data_45; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_46 = proc_10_io_pipe_phv_out_data_46; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_47 = proc_10_io_pipe_phv_out_data_47; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_48 = proc_10_io_pipe_phv_out_data_48; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_49 = proc_10_io_pipe_phv_out_data_49; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_50 = proc_10_io_pipe_phv_out_data_50; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_51 = proc_10_io_pipe_phv_out_data_51; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_52 = proc_10_io_pipe_phv_out_data_52; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_53 = proc_10_io_pipe_phv_out_data_53; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_54 = proc_10_io_pipe_phv_out_data_54; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_55 = proc_10_io_pipe_phv_out_data_55; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_56 = proc_10_io_pipe_phv_out_data_56; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_57 = proc_10_io_pipe_phv_out_data_57; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_58 = proc_10_io_pipe_phv_out_data_58; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_59 = proc_10_io_pipe_phv_out_data_59; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_60 = proc_10_io_pipe_phv_out_data_60; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_61 = proc_10_io_pipe_phv_out_data_61; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_62 = proc_10_io_pipe_phv_out_data_62; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_63 = proc_10_io_pipe_phv_out_data_63; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_64 = proc_10_io_pipe_phv_out_data_64; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_65 = proc_10_io_pipe_phv_out_data_65; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_66 = proc_10_io_pipe_phv_out_data_66; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_67 = proc_10_io_pipe_phv_out_data_67; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_68 = proc_10_io_pipe_phv_out_data_68; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_69 = proc_10_io_pipe_phv_out_data_69; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_70 = proc_10_io_pipe_phv_out_data_70; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_71 = proc_10_io_pipe_phv_out_data_71; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_72 = proc_10_io_pipe_phv_out_data_72; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_73 = proc_10_io_pipe_phv_out_data_73; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_74 = proc_10_io_pipe_phv_out_data_74; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_75 = proc_10_io_pipe_phv_out_data_75; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_76 = proc_10_io_pipe_phv_out_data_76; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_77 = proc_10_io_pipe_phv_out_data_77; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_78 = proc_10_io_pipe_phv_out_data_78; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_79 = proc_10_io_pipe_phv_out_data_79; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_80 = proc_10_io_pipe_phv_out_data_80; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_81 = proc_10_io_pipe_phv_out_data_81; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_82 = proc_10_io_pipe_phv_out_data_82; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_83 = proc_10_io_pipe_phv_out_data_83; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_84 = proc_10_io_pipe_phv_out_data_84; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_85 = proc_10_io_pipe_phv_out_data_85; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_86 = proc_10_io_pipe_phv_out_data_86; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_87 = proc_10_io_pipe_phv_out_data_87; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_88 = proc_10_io_pipe_phv_out_data_88; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_89 = proc_10_io_pipe_phv_out_data_89; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_90 = proc_10_io_pipe_phv_out_data_90; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_91 = proc_10_io_pipe_phv_out_data_91; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_92 = proc_10_io_pipe_phv_out_data_92; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_93 = proc_10_io_pipe_phv_out_data_93; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_94 = proc_10_io_pipe_phv_out_data_94; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_95 = proc_10_io_pipe_phv_out_data_95; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_96 = proc_10_io_pipe_phv_out_data_96; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_97 = proc_10_io_pipe_phv_out_data_97; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_98 = proc_10_io_pipe_phv_out_data_98; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_99 = proc_10_io_pipe_phv_out_data_99; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_100 = proc_10_io_pipe_phv_out_data_100; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_101 = proc_10_io_pipe_phv_out_data_101; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_102 = proc_10_io_pipe_phv_out_data_102; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_103 = proc_10_io_pipe_phv_out_data_103; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_104 = proc_10_io_pipe_phv_out_data_104; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_105 = proc_10_io_pipe_phv_out_data_105; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_106 = proc_10_io_pipe_phv_out_data_106; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_107 = proc_10_io_pipe_phv_out_data_107; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_108 = proc_10_io_pipe_phv_out_data_108; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_109 = proc_10_io_pipe_phv_out_data_109; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_110 = proc_10_io_pipe_phv_out_data_110; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_111 = proc_10_io_pipe_phv_out_data_111; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_112 = proc_10_io_pipe_phv_out_data_112; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_113 = proc_10_io_pipe_phv_out_data_113; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_114 = proc_10_io_pipe_phv_out_data_114; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_115 = proc_10_io_pipe_phv_out_data_115; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_116 = proc_10_io_pipe_phv_out_data_116; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_117 = proc_10_io_pipe_phv_out_data_117; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_118 = proc_10_io_pipe_phv_out_data_118; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_119 = proc_10_io_pipe_phv_out_data_119; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_120 = proc_10_io_pipe_phv_out_data_120; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_121 = proc_10_io_pipe_phv_out_data_121; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_122 = proc_10_io_pipe_phv_out_data_122; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_123 = proc_10_io_pipe_phv_out_data_123; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_124 = proc_10_io_pipe_phv_out_data_124; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_125 = proc_10_io_pipe_phv_out_data_125; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_126 = proc_10_io_pipe_phv_out_data_126; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_127 = proc_10_io_pipe_phv_out_data_127; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_128 = proc_10_io_pipe_phv_out_data_128; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_129 = proc_10_io_pipe_phv_out_data_129; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_130 = proc_10_io_pipe_phv_out_data_130; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_131 = proc_10_io_pipe_phv_out_data_131; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_132 = proc_10_io_pipe_phv_out_data_132; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_133 = proc_10_io_pipe_phv_out_data_133; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_134 = proc_10_io_pipe_phv_out_data_134; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_135 = proc_10_io_pipe_phv_out_data_135; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_136 = proc_10_io_pipe_phv_out_data_136; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_137 = proc_10_io_pipe_phv_out_data_137; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_138 = proc_10_io_pipe_phv_out_data_138; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_139 = proc_10_io_pipe_phv_out_data_139; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_140 = proc_10_io_pipe_phv_out_data_140; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_141 = proc_10_io_pipe_phv_out_data_141; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_142 = proc_10_io_pipe_phv_out_data_142; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_143 = proc_10_io_pipe_phv_out_data_143; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_144 = proc_10_io_pipe_phv_out_data_144; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_145 = proc_10_io_pipe_phv_out_data_145; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_146 = proc_10_io_pipe_phv_out_data_146; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_147 = proc_10_io_pipe_phv_out_data_147; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_148 = proc_10_io_pipe_phv_out_data_148; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_149 = proc_10_io_pipe_phv_out_data_149; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_150 = proc_10_io_pipe_phv_out_data_150; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_151 = proc_10_io_pipe_phv_out_data_151; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_152 = proc_10_io_pipe_phv_out_data_152; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_153 = proc_10_io_pipe_phv_out_data_153; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_154 = proc_10_io_pipe_phv_out_data_154; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_155 = proc_10_io_pipe_phv_out_data_155; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_156 = proc_10_io_pipe_phv_out_data_156; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_157 = proc_10_io_pipe_phv_out_data_157; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_158 = proc_10_io_pipe_phv_out_data_158; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_data_159 = proc_10_io_pipe_phv_out_data_159; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_header_0 = proc_10_io_pipe_phv_out_header_0; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_header_1 = proc_10_io_pipe_phv_out_header_1; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_header_2 = proc_10_io_pipe_phv_out_header_2; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_header_3 = proc_10_io_pipe_phv_out_header_3; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_header_4 = proc_10_io_pipe_phv_out_header_4; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_header_5 = proc_10_io_pipe_phv_out_header_5; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_header_6 = proc_10_io_pipe_phv_out_header_6; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_header_7 = proc_10_io_pipe_phv_out_header_7; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_header_8 = proc_10_io_pipe_phv_out_header_8; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_header_9 = proc_10_io_pipe_phv_out_header_9; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_header_10 = proc_10_io_pipe_phv_out_header_10; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_header_11 = proc_10_io_pipe_phv_out_header_11; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_header_12 = proc_10_io_pipe_phv_out_header_12; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_header_13 = proc_10_io_pipe_phv_out_header_13; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_header_14 = proc_10_io_pipe_phv_out_header_14; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_header_15 = proc_10_io_pipe_phv_out_header_15; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_parse_current_state = proc_10_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_parse_current_offset = proc_10_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_parse_transition_field = proc_10_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_next_processor_id = proc_10_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_next_config_id = proc_10_io_pipe_phv_out_next_config_id; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_valid = proc_10_io_pipe_phv_out_valid; // @[ipsa.scala 82:32]
  assign trans_10_io_pipe_phv_in_last = proc_10_io_pipe_phv_out_last; // @[ipsa.scala 82:32]
  assign trans_10_io_next_proc_exist = 1'h1; // @[ipsa.scala 80:48]
  assign trans_11_clock = clock;
  assign trans_11_io_pipe_phv_in_data_0 = proc_11_io_pipe_phv_out_data_0; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_1 = proc_11_io_pipe_phv_out_data_1; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_2 = proc_11_io_pipe_phv_out_data_2; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_3 = proc_11_io_pipe_phv_out_data_3; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_4 = proc_11_io_pipe_phv_out_data_4; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_5 = proc_11_io_pipe_phv_out_data_5; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_6 = proc_11_io_pipe_phv_out_data_6; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_7 = proc_11_io_pipe_phv_out_data_7; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_8 = proc_11_io_pipe_phv_out_data_8; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_9 = proc_11_io_pipe_phv_out_data_9; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_10 = proc_11_io_pipe_phv_out_data_10; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_11 = proc_11_io_pipe_phv_out_data_11; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_12 = proc_11_io_pipe_phv_out_data_12; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_13 = proc_11_io_pipe_phv_out_data_13; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_14 = proc_11_io_pipe_phv_out_data_14; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_15 = proc_11_io_pipe_phv_out_data_15; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_16 = proc_11_io_pipe_phv_out_data_16; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_17 = proc_11_io_pipe_phv_out_data_17; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_18 = proc_11_io_pipe_phv_out_data_18; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_19 = proc_11_io_pipe_phv_out_data_19; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_20 = proc_11_io_pipe_phv_out_data_20; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_21 = proc_11_io_pipe_phv_out_data_21; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_22 = proc_11_io_pipe_phv_out_data_22; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_23 = proc_11_io_pipe_phv_out_data_23; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_24 = proc_11_io_pipe_phv_out_data_24; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_25 = proc_11_io_pipe_phv_out_data_25; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_26 = proc_11_io_pipe_phv_out_data_26; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_27 = proc_11_io_pipe_phv_out_data_27; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_28 = proc_11_io_pipe_phv_out_data_28; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_29 = proc_11_io_pipe_phv_out_data_29; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_30 = proc_11_io_pipe_phv_out_data_30; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_31 = proc_11_io_pipe_phv_out_data_31; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_32 = proc_11_io_pipe_phv_out_data_32; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_33 = proc_11_io_pipe_phv_out_data_33; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_34 = proc_11_io_pipe_phv_out_data_34; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_35 = proc_11_io_pipe_phv_out_data_35; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_36 = proc_11_io_pipe_phv_out_data_36; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_37 = proc_11_io_pipe_phv_out_data_37; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_38 = proc_11_io_pipe_phv_out_data_38; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_39 = proc_11_io_pipe_phv_out_data_39; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_40 = proc_11_io_pipe_phv_out_data_40; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_41 = proc_11_io_pipe_phv_out_data_41; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_42 = proc_11_io_pipe_phv_out_data_42; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_43 = proc_11_io_pipe_phv_out_data_43; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_44 = proc_11_io_pipe_phv_out_data_44; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_45 = proc_11_io_pipe_phv_out_data_45; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_46 = proc_11_io_pipe_phv_out_data_46; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_47 = proc_11_io_pipe_phv_out_data_47; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_48 = proc_11_io_pipe_phv_out_data_48; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_49 = proc_11_io_pipe_phv_out_data_49; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_50 = proc_11_io_pipe_phv_out_data_50; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_51 = proc_11_io_pipe_phv_out_data_51; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_52 = proc_11_io_pipe_phv_out_data_52; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_53 = proc_11_io_pipe_phv_out_data_53; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_54 = proc_11_io_pipe_phv_out_data_54; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_55 = proc_11_io_pipe_phv_out_data_55; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_56 = proc_11_io_pipe_phv_out_data_56; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_57 = proc_11_io_pipe_phv_out_data_57; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_58 = proc_11_io_pipe_phv_out_data_58; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_59 = proc_11_io_pipe_phv_out_data_59; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_60 = proc_11_io_pipe_phv_out_data_60; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_61 = proc_11_io_pipe_phv_out_data_61; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_62 = proc_11_io_pipe_phv_out_data_62; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_63 = proc_11_io_pipe_phv_out_data_63; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_64 = proc_11_io_pipe_phv_out_data_64; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_65 = proc_11_io_pipe_phv_out_data_65; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_66 = proc_11_io_pipe_phv_out_data_66; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_67 = proc_11_io_pipe_phv_out_data_67; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_68 = proc_11_io_pipe_phv_out_data_68; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_69 = proc_11_io_pipe_phv_out_data_69; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_70 = proc_11_io_pipe_phv_out_data_70; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_71 = proc_11_io_pipe_phv_out_data_71; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_72 = proc_11_io_pipe_phv_out_data_72; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_73 = proc_11_io_pipe_phv_out_data_73; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_74 = proc_11_io_pipe_phv_out_data_74; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_75 = proc_11_io_pipe_phv_out_data_75; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_76 = proc_11_io_pipe_phv_out_data_76; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_77 = proc_11_io_pipe_phv_out_data_77; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_78 = proc_11_io_pipe_phv_out_data_78; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_79 = proc_11_io_pipe_phv_out_data_79; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_80 = proc_11_io_pipe_phv_out_data_80; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_81 = proc_11_io_pipe_phv_out_data_81; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_82 = proc_11_io_pipe_phv_out_data_82; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_83 = proc_11_io_pipe_phv_out_data_83; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_84 = proc_11_io_pipe_phv_out_data_84; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_85 = proc_11_io_pipe_phv_out_data_85; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_86 = proc_11_io_pipe_phv_out_data_86; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_87 = proc_11_io_pipe_phv_out_data_87; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_88 = proc_11_io_pipe_phv_out_data_88; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_89 = proc_11_io_pipe_phv_out_data_89; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_90 = proc_11_io_pipe_phv_out_data_90; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_91 = proc_11_io_pipe_phv_out_data_91; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_92 = proc_11_io_pipe_phv_out_data_92; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_93 = proc_11_io_pipe_phv_out_data_93; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_94 = proc_11_io_pipe_phv_out_data_94; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_95 = proc_11_io_pipe_phv_out_data_95; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_96 = proc_11_io_pipe_phv_out_data_96; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_97 = proc_11_io_pipe_phv_out_data_97; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_98 = proc_11_io_pipe_phv_out_data_98; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_99 = proc_11_io_pipe_phv_out_data_99; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_100 = proc_11_io_pipe_phv_out_data_100; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_101 = proc_11_io_pipe_phv_out_data_101; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_102 = proc_11_io_pipe_phv_out_data_102; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_103 = proc_11_io_pipe_phv_out_data_103; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_104 = proc_11_io_pipe_phv_out_data_104; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_105 = proc_11_io_pipe_phv_out_data_105; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_106 = proc_11_io_pipe_phv_out_data_106; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_107 = proc_11_io_pipe_phv_out_data_107; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_108 = proc_11_io_pipe_phv_out_data_108; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_109 = proc_11_io_pipe_phv_out_data_109; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_110 = proc_11_io_pipe_phv_out_data_110; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_111 = proc_11_io_pipe_phv_out_data_111; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_112 = proc_11_io_pipe_phv_out_data_112; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_113 = proc_11_io_pipe_phv_out_data_113; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_114 = proc_11_io_pipe_phv_out_data_114; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_115 = proc_11_io_pipe_phv_out_data_115; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_116 = proc_11_io_pipe_phv_out_data_116; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_117 = proc_11_io_pipe_phv_out_data_117; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_118 = proc_11_io_pipe_phv_out_data_118; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_119 = proc_11_io_pipe_phv_out_data_119; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_120 = proc_11_io_pipe_phv_out_data_120; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_121 = proc_11_io_pipe_phv_out_data_121; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_122 = proc_11_io_pipe_phv_out_data_122; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_123 = proc_11_io_pipe_phv_out_data_123; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_124 = proc_11_io_pipe_phv_out_data_124; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_125 = proc_11_io_pipe_phv_out_data_125; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_126 = proc_11_io_pipe_phv_out_data_126; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_127 = proc_11_io_pipe_phv_out_data_127; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_128 = proc_11_io_pipe_phv_out_data_128; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_129 = proc_11_io_pipe_phv_out_data_129; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_130 = proc_11_io_pipe_phv_out_data_130; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_131 = proc_11_io_pipe_phv_out_data_131; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_132 = proc_11_io_pipe_phv_out_data_132; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_133 = proc_11_io_pipe_phv_out_data_133; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_134 = proc_11_io_pipe_phv_out_data_134; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_135 = proc_11_io_pipe_phv_out_data_135; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_136 = proc_11_io_pipe_phv_out_data_136; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_137 = proc_11_io_pipe_phv_out_data_137; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_138 = proc_11_io_pipe_phv_out_data_138; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_139 = proc_11_io_pipe_phv_out_data_139; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_140 = proc_11_io_pipe_phv_out_data_140; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_141 = proc_11_io_pipe_phv_out_data_141; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_142 = proc_11_io_pipe_phv_out_data_142; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_143 = proc_11_io_pipe_phv_out_data_143; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_144 = proc_11_io_pipe_phv_out_data_144; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_145 = proc_11_io_pipe_phv_out_data_145; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_146 = proc_11_io_pipe_phv_out_data_146; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_147 = proc_11_io_pipe_phv_out_data_147; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_148 = proc_11_io_pipe_phv_out_data_148; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_149 = proc_11_io_pipe_phv_out_data_149; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_150 = proc_11_io_pipe_phv_out_data_150; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_151 = proc_11_io_pipe_phv_out_data_151; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_152 = proc_11_io_pipe_phv_out_data_152; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_153 = proc_11_io_pipe_phv_out_data_153; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_154 = proc_11_io_pipe_phv_out_data_154; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_155 = proc_11_io_pipe_phv_out_data_155; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_156 = proc_11_io_pipe_phv_out_data_156; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_157 = proc_11_io_pipe_phv_out_data_157; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_158 = proc_11_io_pipe_phv_out_data_158; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_data_159 = proc_11_io_pipe_phv_out_data_159; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_header_0 = proc_11_io_pipe_phv_out_header_0; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_header_1 = proc_11_io_pipe_phv_out_header_1; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_header_2 = proc_11_io_pipe_phv_out_header_2; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_header_3 = proc_11_io_pipe_phv_out_header_3; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_header_4 = proc_11_io_pipe_phv_out_header_4; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_header_5 = proc_11_io_pipe_phv_out_header_5; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_header_6 = proc_11_io_pipe_phv_out_header_6; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_header_7 = proc_11_io_pipe_phv_out_header_7; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_header_8 = proc_11_io_pipe_phv_out_header_8; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_header_9 = proc_11_io_pipe_phv_out_header_9; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_header_10 = proc_11_io_pipe_phv_out_header_10; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_header_11 = proc_11_io_pipe_phv_out_header_11; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_header_12 = proc_11_io_pipe_phv_out_header_12; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_header_13 = proc_11_io_pipe_phv_out_header_13; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_header_14 = proc_11_io_pipe_phv_out_header_14; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_header_15 = proc_11_io_pipe_phv_out_header_15; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_parse_current_state = proc_11_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_parse_current_offset = proc_11_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_parse_transition_field = proc_11_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_next_processor_id = proc_11_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_next_config_id = proc_11_io_pipe_phv_out_next_config_id; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_valid = proc_11_io_pipe_phv_out_valid; // @[ipsa.scala 82:32]
  assign trans_11_io_pipe_phv_in_last = proc_11_io_pipe_phv_out_last; // @[ipsa.scala 82:32]
  assign trans_11_io_next_proc_exist = 1'h1; // @[ipsa.scala 80:48]
  assign trans_12_clock = clock;
  assign trans_12_io_pipe_phv_in_data_0 = proc_12_io_pipe_phv_out_data_0; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_1 = proc_12_io_pipe_phv_out_data_1; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_2 = proc_12_io_pipe_phv_out_data_2; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_3 = proc_12_io_pipe_phv_out_data_3; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_4 = proc_12_io_pipe_phv_out_data_4; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_5 = proc_12_io_pipe_phv_out_data_5; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_6 = proc_12_io_pipe_phv_out_data_6; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_7 = proc_12_io_pipe_phv_out_data_7; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_8 = proc_12_io_pipe_phv_out_data_8; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_9 = proc_12_io_pipe_phv_out_data_9; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_10 = proc_12_io_pipe_phv_out_data_10; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_11 = proc_12_io_pipe_phv_out_data_11; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_12 = proc_12_io_pipe_phv_out_data_12; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_13 = proc_12_io_pipe_phv_out_data_13; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_14 = proc_12_io_pipe_phv_out_data_14; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_15 = proc_12_io_pipe_phv_out_data_15; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_16 = proc_12_io_pipe_phv_out_data_16; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_17 = proc_12_io_pipe_phv_out_data_17; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_18 = proc_12_io_pipe_phv_out_data_18; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_19 = proc_12_io_pipe_phv_out_data_19; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_20 = proc_12_io_pipe_phv_out_data_20; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_21 = proc_12_io_pipe_phv_out_data_21; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_22 = proc_12_io_pipe_phv_out_data_22; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_23 = proc_12_io_pipe_phv_out_data_23; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_24 = proc_12_io_pipe_phv_out_data_24; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_25 = proc_12_io_pipe_phv_out_data_25; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_26 = proc_12_io_pipe_phv_out_data_26; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_27 = proc_12_io_pipe_phv_out_data_27; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_28 = proc_12_io_pipe_phv_out_data_28; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_29 = proc_12_io_pipe_phv_out_data_29; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_30 = proc_12_io_pipe_phv_out_data_30; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_31 = proc_12_io_pipe_phv_out_data_31; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_32 = proc_12_io_pipe_phv_out_data_32; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_33 = proc_12_io_pipe_phv_out_data_33; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_34 = proc_12_io_pipe_phv_out_data_34; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_35 = proc_12_io_pipe_phv_out_data_35; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_36 = proc_12_io_pipe_phv_out_data_36; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_37 = proc_12_io_pipe_phv_out_data_37; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_38 = proc_12_io_pipe_phv_out_data_38; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_39 = proc_12_io_pipe_phv_out_data_39; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_40 = proc_12_io_pipe_phv_out_data_40; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_41 = proc_12_io_pipe_phv_out_data_41; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_42 = proc_12_io_pipe_phv_out_data_42; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_43 = proc_12_io_pipe_phv_out_data_43; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_44 = proc_12_io_pipe_phv_out_data_44; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_45 = proc_12_io_pipe_phv_out_data_45; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_46 = proc_12_io_pipe_phv_out_data_46; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_47 = proc_12_io_pipe_phv_out_data_47; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_48 = proc_12_io_pipe_phv_out_data_48; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_49 = proc_12_io_pipe_phv_out_data_49; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_50 = proc_12_io_pipe_phv_out_data_50; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_51 = proc_12_io_pipe_phv_out_data_51; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_52 = proc_12_io_pipe_phv_out_data_52; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_53 = proc_12_io_pipe_phv_out_data_53; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_54 = proc_12_io_pipe_phv_out_data_54; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_55 = proc_12_io_pipe_phv_out_data_55; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_56 = proc_12_io_pipe_phv_out_data_56; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_57 = proc_12_io_pipe_phv_out_data_57; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_58 = proc_12_io_pipe_phv_out_data_58; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_59 = proc_12_io_pipe_phv_out_data_59; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_60 = proc_12_io_pipe_phv_out_data_60; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_61 = proc_12_io_pipe_phv_out_data_61; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_62 = proc_12_io_pipe_phv_out_data_62; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_63 = proc_12_io_pipe_phv_out_data_63; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_64 = proc_12_io_pipe_phv_out_data_64; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_65 = proc_12_io_pipe_phv_out_data_65; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_66 = proc_12_io_pipe_phv_out_data_66; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_67 = proc_12_io_pipe_phv_out_data_67; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_68 = proc_12_io_pipe_phv_out_data_68; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_69 = proc_12_io_pipe_phv_out_data_69; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_70 = proc_12_io_pipe_phv_out_data_70; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_71 = proc_12_io_pipe_phv_out_data_71; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_72 = proc_12_io_pipe_phv_out_data_72; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_73 = proc_12_io_pipe_phv_out_data_73; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_74 = proc_12_io_pipe_phv_out_data_74; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_75 = proc_12_io_pipe_phv_out_data_75; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_76 = proc_12_io_pipe_phv_out_data_76; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_77 = proc_12_io_pipe_phv_out_data_77; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_78 = proc_12_io_pipe_phv_out_data_78; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_79 = proc_12_io_pipe_phv_out_data_79; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_80 = proc_12_io_pipe_phv_out_data_80; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_81 = proc_12_io_pipe_phv_out_data_81; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_82 = proc_12_io_pipe_phv_out_data_82; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_83 = proc_12_io_pipe_phv_out_data_83; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_84 = proc_12_io_pipe_phv_out_data_84; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_85 = proc_12_io_pipe_phv_out_data_85; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_86 = proc_12_io_pipe_phv_out_data_86; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_87 = proc_12_io_pipe_phv_out_data_87; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_88 = proc_12_io_pipe_phv_out_data_88; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_89 = proc_12_io_pipe_phv_out_data_89; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_90 = proc_12_io_pipe_phv_out_data_90; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_91 = proc_12_io_pipe_phv_out_data_91; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_92 = proc_12_io_pipe_phv_out_data_92; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_93 = proc_12_io_pipe_phv_out_data_93; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_94 = proc_12_io_pipe_phv_out_data_94; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_95 = proc_12_io_pipe_phv_out_data_95; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_96 = proc_12_io_pipe_phv_out_data_96; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_97 = proc_12_io_pipe_phv_out_data_97; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_98 = proc_12_io_pipe_phv_out_data_98; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_99 = proc_12_io_pipe_phv_out_data_99; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_100 = proc_12_io_pipe_phv_out_data_100; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_101 = proc_12_io_pipe_phv_out_data_101; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_102 = proc_12_io_pipe_phv_out_data_102; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_103 = proc_12_io_pipe_phv_out_data_103; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_104 = proc_12_io_pipe_phv_out_data_104; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_105 = proc_12_io_pipe_phv_out_data_105; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_106 = proc_12_io_pipe_phv_out_data_106; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_107 = proc_12_io_pipe_phv_out_data_107; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_108 = proc_12_io_pipe_phv_out_data_108; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_109 = proc_12_io_pipe_phv_out_data_109; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_110 = proc_12_io_pipe_phv_out_data_110; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_111 = proc_12_io_pipe_phv_out_data_111; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_112 = proc_12_io_pipe_phv_out_data_112; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_113 = proc_12_io_pipe_phv_out_data_113; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_114 = proc_12_io_pipe_phv_out_data_114; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_115 = proc_12_io_pipe_phv_out_data_115; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_116 = proc_12_io_pipe_phv_out_data_116; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_117 = proc_12_io_pipe_phv_out_data_117; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_118 = proc_12_io_pipe_phv_out_data_118; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_119 = proc_12_io_pipe_phv_out_data_119; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_120 = proc_12_io_pipe_phv_out_data_120; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_121 = proc_12_io_pipe_phv_out_data_121; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_122 = proc_12_io_pipe_phv_out_data_122; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_123 = proc_12_io_pipe_phv_out_data_123; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_124 = proc_12_io_pipe_phv_out_data_124; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_125 = proc_12_io_pipe_phv_out_data_125; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_126 = proc_12_io_pipe_phv_out_data_126; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_127 = proc_12_io_pipe_phv_out_data_127; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_128 = proc_12_io_pipe_phv_out_data_128; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_129 = proc_12_io_pipe_phv_out_data_129; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_130 = proc_12_io_pipe_phv_out_data_130; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_131 = proc_12_io_pipe_phv_out_data_131; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_132 = proc_12_io_pipe_phv_out_data_132; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_133 = proc_12_io_pipe_phv_out_data_133; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_134 = proc_12_io_pipe_phv_out_data_134; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_135 = proc_12_io_pipe_phv_out_data_135; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_136 = proc_12_io_pipe_phv_out_data_136; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_137 = proc_12_io_pipe_phv_out_data_137; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_138 = proc_12_io_pipe_phv_out_data_138; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_139 = proc_12_io_pipe_phv_out_data_139; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_140 = proc_12_io_pipe_phv_out_data_140; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_141 = proc_12_io_pipe_phv_out_data_141; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_142 = proc_12_io_pipe_phv_out_data_142; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_143 = proc_12_io_pipe_phv_out_data_143; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_144 = proc_12_io_pipe_phv_out_data_144; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_145 = proc_12_io_pipe_phv_out_data_145; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_146 = proc_12_io_pipe_phv_out_data_146; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_147 = proc_12_io_pipe_phv_out_data_147; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_148 = proc_12_io_pipe_phv_out_data_148; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_149 = proc_12_io_pipe_phv_out_data_149; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_150 = proc_12_io_pipe_phv_out_data_150; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_151 = proc_12_io_pipe_phv_out_data_151; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_152 = proc_12_io_pipe_phv_out_data_152; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_153 = proc_12_io_pipe_phv_out_data_153; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_154 = proc_12_io_pipe_phv_out_data_154; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_155 = proc_12_io_pipe_phv_out_data_155; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_156 = proc_12_io_pipe_phv_out_data_156; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_157 = proc_12_io_pipe_phv_out_data_157; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_158 = proc_12_io_pipe_phv_out_data_158; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_data_159 = proc_12_io_pipe_phv_out_data_159; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_header_0 = proc_12_io_pipe_phv_out_header_0; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_header_1 = proc_12_io_pipe_phv_out_header_1; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_header_2 = proc_12_io_pipe_phv_out_header_2; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_header_3 = proc_12_io_pipe_phv_out_header_3; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_header_4 = proc_12_io_pipe_phv_out_header_4; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_header_5 = proc_12_io_pipe_phv_out_header_5; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_header_6 = proc_12_io_pipe_phv_out_header_6; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_header_7 = proc_12_io_pipe_phv_out_header_7; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_header_8 = proc_12_io_pipe_phv_out_header_8; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_header_9 = proc_12_io_pipe_phv_out_header_9; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_header_10 = proc_12_io_pipe_phv_out_header_10; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_header_11 = proc_12_io_pipe_phv_out_header_11; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_header_12 = proc_12_io_pipe_phv_out_header_12; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_header_13 = proc_12_io_pipe_phv_out_header_13; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_header_14 = proc_12_io_pipe_phv_out_header_14; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_header_15 = proc_12_io_pipe_phv_out_header_15; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_parse_current_state = proc_12_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_parse_current_offset = proc_12_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_parse_transition_field = proc_12_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_next_processor_id = proc_12_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_next_config_id = proc_12_io_pipe_phv_out_next_config_id; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_valid = proc_12_io_pipe_phv_out_valid; // @[ipsa.scala 82:32]
  assign trans_12_io_pipe_phv_in_last = proc_12_io_pipe_phv_out_last; // @[ipsa.scala 82:32]
  assign trans_12_io_next_proc_exist = 1'h1; // @[ipsa.scala 80:48]
  assign trans_13_clock = clock;
  assign trans_13_io_pipe_phv_in_data_0 = proc_13_io_pipe_phv_out_data_0; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_1 = proc_13_io_pipe_phv_out_data_1; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_2 = proc_13_io_pipe_phv_out_data_2; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_3 = proc_13_io_pipe_phv_out_data_3; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_4 = proc_13_io_pipe_phv_out_data_4; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_5 = proc_13_io_pipe_phv_out_data_5; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_6 = proc_13_io_pipe_phv_out_data_6; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_7 = proc_13_io_pipe_phv_out_data_7; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_8 = proc_13_io_pipe_phv_out_data_8; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_9 = proc_13_io_pipe_phv_out_data_9; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_10 = proc_13_io_pipe_phv_out_data_10; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_11 = proc_13_io_pipe_phv_out_data_11; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_12 = proc_13_io_pipe_phv_out_data_12; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_13 = proc_13_io_pipe_phv_out_data_13; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_14 = proc_13_io_pipe_phv_out_data_14; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_15 = proc_13_io_pipe_phv_out_data_15; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_16 = proc_13_io_pipe_phv_out_data_16; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_17 = proc_13_io_pipe_phv_out_data_17; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_18 = proc_13_io_pipe_phv_out_data_18; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_19 = proc_13_io_pipe_phv_out_data_19; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_20 = proc_13_io_pipe_phv_out_data_20; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_21 = proc_13_io_pipe_phv_out_data_21; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_22 = proc_13_io_pipe_phv_out_data_22; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_23 = proc_13_io_pipe_phv_out_data_23; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_24 = proc_13_io_pipe_phv_out_data_24; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_25 = proc_13_io_pipe_phv_out_data_25; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_26 = proc_13_io_pipe_phv_out_data_26; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_27 = proc_13_io_pipe_phv_out_data_27; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_28 = proc_13_io_pipe_phv_out_data_28; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_29 = proc_13_io_pipe_phv_out_data_29; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_30 = proc_13_io_pipe_phv_out_data_30; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_31 = proc_13_io_pipe_phv_out_data_31; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_32 = proc_13_io_pipe_phv_out_data_32; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_33 = proc_13_io_pipe_phv_out_data_33; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_34 = proc_13_io_pipe_phv_out_data_34; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_35 = proc_13_io_pipe_phv_out_data_35; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_36 = proc_13_io_pipe_phv_out_data_36; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_37 = proc_13_io_pipe_phv_out_data_37; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_38 = proc_13_io_pipe_phv_out_data_38; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_39 = proc_13_io_pipe_phv_out_data_39; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_40 = proc_13_io_pipe_phv_out_data_40; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_41 = proc_13_io_pipe_phv_out_data_41; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_42 = proc_13_io_pipe_phv_out_data_42; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_43 = proc_13_io_pipe_phv_out_data_43; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_44 = proc_13_io_pipe_phv_out_data_44; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_45 = proc_13_io_pipe_phv_out_data_45; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_46 = proc_13_io_pipe_phv_out_data_46; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_47 = proc_13_io_pipe_phv_out_data_47; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_48 = proc_13_io_pipe_phv_out_data_48; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_49 = proc_13_io_pipe_phv_out_data_49; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_50 = proc_13_io_pipe_phv_out_data_50; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_51 = proc_13_io_pipe_phv_out_data_51; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_52 = proc_13_io_pipe_phv_out_data_52; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_53 = proc_13_io_pipe_phv_out_data_53; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_54 = proc_13_io_pipe_phv_out_data_54; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_55 = proc_13_io_pipe_phv_out_data_55; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_56 = proc_13_io_pipe_phv_out_data_56; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_57 = proc_13_io_pipe_phv_out_data_57; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_58 = proc_13_io_pipe_phv_out_data_58; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_59 = proc_13_io_pipe_phv_out_data_59; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_60 = proc_13_io_pipe_phv_out_data_60; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_61 = proc_13_io_pipe_phv_out_data_61; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_62 = proc_13_io_pipe_phv_out_data_62; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_63 = proc_13_io_pipe_phv_out_data_63; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_64 = proc_13_io_pipe_phv_out_data_64; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_65 = proc_13_io_pipe_phv_out_data_65; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_66 = proc_13_io_pipe_phv_out_data_66; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_67 = proc_13_io_pipe_phv_out_data_67; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_68 = proc_13_io_pipe_phv_out_data_68; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_69 = proc_13_io_pipe_phv_out_data_69; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_70 = proc_13_io_pipe_phv_out_data_70; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_71 = proc_13_io_pipe_phv_out_data_71; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_72 = proc_13_io_pipe_phv_out_data_72; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_73 = proc_13_io_pipe_phv_out_data_73; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_74 = proc_13_io_pipe_phv_out_data_74; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_75 = proc_13_io_pipe_phv_out_data_75; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_76 = proc_13_io_pipe_phv_out_data_76; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_77 = proc_13_io_pipe_phv_out_data_77; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_78 = proc_13_io_pipe_phv_out_data_78; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_79 = proc_13_io_pipe_phv_out_data_79; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_80 = proc_13_io_pipe_phv_out_data_80; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_81 = proc_13_io_pipe_phv_out_data_81; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_82 = proc_13_io_pipe_phv_out_data_82; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_83 = proc_13_io_pipe_phv_out_data_83; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_84 = proc_13_io_pipe_phv_out_data_84; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_85 = proc_13_io_pipe_phv_out_data_85; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_86 = proc_13_io_pipe_phv_out_data_86; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_87 = proc_13_io_pipe_phv_out_data_87; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_88 = proc_13_io_pipe_phv_out_data_88; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_89 = proc_13_io_pipe_phv_out_data_89; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_90 = proc_13_io_pipe_phv_out_data_90; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_91 = proc_13_io_pipe_phv_out_data_91; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_92 = proc_13_io_pipe_phv_out_data_92; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_93 = proc_13_io_pipe_phv_out_data_93; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_94 = proc_13_io_pipe_phv_out_data_94; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_95 = proc_13_io_pipe_phv_out_data_95; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_96 = proc_13_io_pipe_phv_out_data_96; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_97 = proc_13_io_pipe_phv_out_data_97; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_98 = proc_13_io_pipe_phv_out_data_98; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_99 = proc_13_io_pipe_phv_out_data_99; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_100 = proc_13_io_pipe_phv_out_data_100; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_101 = proc_13_io_pipe_phv_out_data_101; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_102 = proc_13_io_pipe_phv_out_data_102; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_103 = proc_13_io_pipe_phv_out_data_103; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_104 = proc_13_io_pipe_phv_out_data_104; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_105 = proc_13_io_pipe_phv_out_data_105; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_106 = proc_13_io_pipe_phv_out_data_106; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_107 = proc_13_io_pipe_phv_out_data_107; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_108 = proc_13_io_pipe_phv_out_data_108; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_109 = proc_13_io_pipe_phv_out_data_109; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_110 = proc_13_io_pipe_phv_out_data_110; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_111 = proc_13_io_pipe_phv_out_data_111; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_112 = proc_13_io_pipe_phv_out_data_112; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_113 = proc_13_io_pipe_phv_out_data_113; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_114 = proc_13_io_pipe_phv_out_data_114; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_115 = proc_13_io_pipe_phv_out_data_115; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_116 = proc_13_io_pipe_phv_out_data_116; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_117 = proc_13_io_pipe_phv_out_data_117; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_118 = proc_13_io_pipe_phv_out_data_118; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_119 = proc_13_io_pipe_phv_out_data_119; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_120 = proc_13_io_pipe_phv_out_data_120; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_121 = proc_13_io_pipe_phv_out_data_121; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_122 = proc_13_io_pipe_phv_out_data_122; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_123 = proc_13_io_pipe_phv_out_data_123; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_124 = proc_13_io_pipe_phv_out_data_124; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_125 = proc_13_io_pipe_phv_out_data_125; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_126 = proc_13_io_pipe_phv_out_data_126; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_127 = proc_13_io_pipe_phv_out_data_127; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_128 = proc_13_io_pipe_phv_out_data_128; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_129 = proc_13_io_pipe_phv_out_data_129; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_130 = proc_13_io_pipe_phv_out_data_130; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_131 = proc_13_io_pipe_phv_out_data_131; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_132 = proc_13_io_pipe_phv_out_data_132; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_133 = proc_13_io_pipe_phv_out_data_133; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_134 = proc_13_io_pipe_phv_out_data_134; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_135 = proc_13_io_pipe_phv_out_data_135; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_136 = proc_13_io_pipe_phv_out_data_136; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_137 = proc_13_io_pipe_phv_out_data_137; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_138 = proc_13_io_pipe_phv_out_data_138; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_139 = proc_13_io_pipe_phv_out_data_139; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_140 = proc_13_io_pipe_phv_out_data_140; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_141 = proc_13_io_pipe_phv_out_data_141; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_142 = proc_13_io_pipe_phv_out_data_142; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_143 = proc_13_io_pipe_phv_out_data_143; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_144 = proc_13_io_pipe_phv_out_data_144; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_145 = proc_13_io_pipe_phv_out_data_145; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_146 = proc_13_io_pipe_phv_out_data_146; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_147 = proc_13_io_pipe_phv_out_data_147; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_148 = proc_13_io_pipe_phv_out_data_148; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_149 = proc_13_io_pipe_phv_out_data_149; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_150 = proc_13_io_pipe_phv_out_data_150; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_151 = proc_13_io_pipe_phv_out_data_151; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_152 = proc_13_io_pipe_phv_out_data_152; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_153 = proc_13_io_pipe_phv_out_data_153; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_154 = proc_13_io_pipe_phv_out_data_154; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_155 = proc_13_io_pipe_phv_out_data_155; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_156 = proc_13_io_pipe_phv_out_data_156; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_157 = proc_13_io_pipe_phv_out_data_157; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_158 = proc_13_io_pipe_phv_out_data_158; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_data_159 = proc_13_io_pipe_phv_out_data_159; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_header_0 = proc_13_io_pipe_phv_out_header_0; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_header_1 = proc_13_io_pipe_phv_out_header_1; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_header_2 = proc_13_io_pipe_phv_out_header_2; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_header_3 = proc_13_io_pipe_phv_out_header_3; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_header_4 = proc_13_io_pipe_phv_out_header_4; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_header_5 = proc_13_io_pipe_phv_out_header_5; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_header_6 = proc_13_io_pipe_phv_out_header_6; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_header_7 = proc_13_io_pipe_phv_out_header_7; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_header_8 = proc_13_io_pipe_phv_out_header_8; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_header_9 = proc_13_io_pipe_phv_out_header_9; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_header_10 = proc_13_io_pipe_phv_out_header_10; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_header_11 = proc_13_io_pipe_phv_out_header_11; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_header_12 = proc_13_io_pipe_phv_out_header_12; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_header_13 = proc_13_io_pipe_phv_out_header_13; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_header_14 = proc_13_io_pipe_phv_out_header_14; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_header_15 = proc_13_io_pipe_phv_out_header_15; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_parse_current_state = proc_13_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_parse_current_offset = proc_13_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_parse_transition_field = proc_13_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_next_processor_id = proc_13_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_next_config_id = proc_13_io_pipe_phv_out_next_config_id; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_valid = proc_13_io_pipe_phv_out_valid; // @[ipsa.scala 82:32]
  assign trans_13_io_pipe_phv_in_last = proc_13_io_pipe_phv_out_last; // @[ipsa.scala 82:32]
  assign trans_13_io_next_proc_exist = 1'h1; // @[ipsa.scala 80:48]
  assign trans_14_clock = clock;
  assign trans_14_io_pipe_phv_in_data_0 = proc_14_io_pipe_phv_out_data_0; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_1 = proc_14_io_pipe_phv_out_data_1; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_2 = proc_14_io_pipe_phv_out_data_2; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_3 = proc_14_io_pipe_phv_out_data_3; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_4 = proc_14_io_pipe_phv_out_data_4; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_5 = proc_14_io_pipe_phv_out_data_5; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_6 = proc_14_io_pipe_phv_out_data_6; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_7 = proc_14_io_pipe_phv_out_data_7; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_8 = proc_14_io_pipe_phv_out_data_8; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_9 = proc_14_io_pipe_phv_out_data_9; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_10 = proc_14_io_pipe_phv_out_data_10; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_11 = proc_14_io_pipe_phv_out_data_11; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_12 = proc_14_io_pipe_phv_out_data_12; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_13 = proc_14_io_pipe_phv_out_data_13; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_14 = proc_14_io_pipe_phv_out_data_14; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_15 = proc_14_io_pipe_phv_out_data_15; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_16 = proc_14_io_pipe_phv_out_data_16; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_17 = proc_14_io_pipe_phv_out_data_17; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_18 = proc_14_io_pipe_phv_out_data_18; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_19 = proc_14_io_pipe_phv_out_data_19; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_20 = proc_14_io_pipe_phv_out_data_20; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_21 = proc_14_io_pipe_phv_out_data_21; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_22 = proc_14_io_pipe_phv_out_data_22; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_23 = proc_14_io_pipe_phv_out_data_23; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_24 = proc_14_io_pipe_phv_out_data_24; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_25 = proc_14_io_pipe_phv_out_data_25; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_26 = proc_14_io_pipe_phv_out_data_26; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_27 = proc_14_io_pipe_phv_out_data_27; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_28 = proc_14_io_pipe_phv_out_data_28; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_29 = proc_14_io_pipe_phv_out_data_29; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_30 = proc_14_io_pipe_phv_out_data_30; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_31 = proc_14_io_pipe_phv_out_data_31; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_32 = proc_14_io_pipe_phv_out_data_32; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_33 = proc_14_io_pipe_phv_out_data_33; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_34 = proc_14_io_pipe_phv_out_data_34; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_35 = proc_14_io_pipe_phv_out_data_35; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_36 = proc_14_io_pipe_phv_out_data_36; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_37 = proc_14_io_pipe_phv_out_data_37; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_38 = proc_14_io_pipe_phv_out_data_38; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_39 = proc_14_io_pipe_phv_out_data_39; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_40 = proc_14_io_pipe_phv_out_data_40; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_41 = proc_14_io_pipe_phv_out_data_41; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_42 = proc_14_io_pipe_phv_out_data_42; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_43 = proc_14_io_pipe_phv_out_data_43; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_44 = proc_14_io_pipe_phv_out_data_44; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_45 = proc_14_io_pipe_phv_out_data_45; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_46 = proc_14_io_pipe_phv_out_data_46; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_47 = proc_14_io_pipe_phv_out_data_47; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_48 = proc_14_io_pipe_phv_out_data_48; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_49 = proc_14_io_pipe_phv_out_data_49; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_50 = proc_14_io_pipe_phv_out_data_50; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_51 = proc_14_io_pipe_phv_out_data_51; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_52 = proc_14_io_pipe_phv_out_data_52; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_53 = proc_14_io_pipe_phv_out_data_53; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_54 = proc_14_io_pipe_phv_out_data_54; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_55 = proc_14_io_pipe_phv_out_data_55; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_56 = proc_14_io_pipe_phv_out_data_56; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_57 = proc_14_io_pipe_phv_out_data_57; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_58 = proc_14_io_pipe_phv_out_data_58; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_59 = proc_14_io_pipe_phv_out_data_59; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_60 = proc_14_io_pipe_phv_out_data_60; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_61 = proc_14_io_pipe_phv_out_data_61; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_62 = proc_14_io_pipe_phv_out_data_62; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_63 = proc_14_io_pipe_phv_out_data_63; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_64 = proc_14_io_pipe_phv_out_data_64; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_65 = proc_14_io_pipe_phv_out_data_65; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_66 = proc_14_io_pipe_phv_out_data_66; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_67 = proc_14_io_pipe_phv_out_data_67; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_68 = proc_14_io_pipe_phv_out_data_68; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_69 = proc_14_io_pipe_phv_out_data_69; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_70 = proc_14_io_pipe_phv_out_data_70; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_71 = proc_14_io_pipe_phv_out_data_71; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_72 = proc_14_io_pipe_phv_out_data_72; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_73 = proc_14_io_pipe_phv_out_data_73; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_74 = proc_14_io_pipe_phv_out_data_74; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_75 = proc_14_io_pipe_phv_out_data_75; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_76 = proc_14_io_pipe_phv_out_data_76; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_77 = proc_14_io_pipe_phv_out_data_77; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_78 = proc_14_io_pipe_phv_out_data_78; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_79 = proc_14_io_pipe_phv_out_data_79; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_80 = proc_14_io_pipe_phv_out_data_80; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_81 = proc_14_io_pipe_phv_out_data_81; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_82 = proc_14_io_pipe_phv_out_data_82; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_83 = proc_14_io_pipe_phv_out_data_83; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_84 = proc_14_io_pipe_phv_out_data_84; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_85 = proc_14_io_pipe_phv_out_data_85; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_86 = proc_14_io_pipe_phv_out_data_86; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_87 = proc_14_io_pipe_phv_out_data_87; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_88 = proc_14_io_pipe_phv_out_data_88; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_89 = proc_14_io_pipe_phv_out_data_89; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_90 = proc_14_io_pipe_phv_out_data_90; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_91 = proc_14_io_pipe_phv_out_data_91; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_92 = proc_14_io_pipe_phv_out_data_92; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_93 = proc_14_io_pipe_phv_out_data_93; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_94 = proc_14_io_pipe_phv_out_data_94; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_95 = proc_14_io_pipe_phv_out_data_95; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_96 = proc_14_io_pipe_phv_out_data_96; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_97 = proc_14_io_pipe_phv_out_data_97; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_98 = proc_14_io_pipe_phv_out_data_98; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_99 = proc_14_io_pipe_phv_out_data_99; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_100 = proc_14_io_pipe_phv_out_data_100; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_101 = proc_14_io_pipe_phv_out_data_101; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_102 = proc_14_io_pipe_phv_out_data_102; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_103 = proc_14_io_pipe_phv_out_data_103; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_104 = proc_14_io_pipe_phv_out_data_104; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_105 = proc_14_io_pipe_phv_out_data_105; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_106 = proc_14_io_pipe_phv_out_data_106; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_107 = proc_14_io_pipe_phv_out_data_107; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_108 = proc_14_io_pipe_phv_out_data_108; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_109 = proc_14_io_pipe_phv_out_data_109; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_110 = proc_14_io_pipe_phv_out_data_110; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_111 = proc_14_io_pipe_phv_out_data_111; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_112 = proc_14_io_pipe_phv_out_data_112; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_113 = proc_14_io_pipe_phv_out_data_113; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_114 = proc_14_io_pipe_phv_out_data_114; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_115 = proc_14_io_pipe_phv_out_data_115; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_116 = proc_14_io_pipe_phv_out_data_116; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_117 = proc_14_io_pipe_phv_out_data_117; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_118 = proc_14_io_pipe_phv_out_data_118; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_119 = proc_14_io_pipe_phv_out_data_119; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_120 = proc_14_io_pipe_phv_out_data_120; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_121 = proc_14_io_pipe_phv_out_data_121; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_122 = proc_14_io_pipe_phv_out_data_122; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_123 = proc_14_io_pipe_phv_out_data_123; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_124 = proc_14_io_pipe_phv_out_data_124; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_125 = proc_14_io_pipe_phv_out_data_125; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_126 = proc_14_io_pipe_phv_out_data_126; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_127 = proc_14_io_pipe_phv_out_data_127; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_128 = proc_14_io_pipe_phv_out_data_128; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_129 = proc_14_io_pipe_phv_out_data_129; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_130 = proc_14_io_pipe_phv_out_data_130; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_131 = proc_14_io_pipe_phv_out_data_131; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_132 = proc_14_io_pipe_phv_out_data_132; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_133 = proc_14_io_pipe_phv_out_data_133; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_134 = proc_14_io_pipe_phv_out_data_134; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_135 = proc_14_io_pipe_phv_out_data_135; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_136 = proc_14_io_pipe_phv_out_data_136; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_137 = proc_14_io_pipe_phv_out_data_137; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_138 = proc_14_io_pipe_phv_out_data_138; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_139 = proc_14_io_pipe_phv_out_data_139; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_140 = proc_14_io_pipe_phv_out_data_140; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_141 = proc_14_io_pipe_phv_out_data_141; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_142 = proc_14_io_pipe_phv_out_data_142; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_143 = proc_14_io_pipe_phv_out_data_143; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_144 = proc_14_io_pipe_phv_out_data_144; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_145 = proc_14_io_pipe_phv_out_data_145; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_146 = proc_14_io_pipe_phv_out_data_146; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_147 = proc_14_io_pipe_phv_out_data_147; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_148 = proc_14_io_pipe_phv_out_data_148; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_149 = proc_14_io_pipe_phv_out_data_149; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_150 = proc_14_io_pipe_phv_out_data_150; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_151 = proc_14_io_pipe_phv_out_data_151; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_152 = proc_14_io_pipe_phv_out_data_152; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_153 = proc_14_io_pipe_phv_out_data_153; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_154 = proc_14_io_pipe_phv_out_data_154; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_155 = proc_14_io_pipe_phv_out_data_155; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_156 = proc_14_io_pipe_phv_out_data_156; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_157 = proc_14_io_pipe_phv_out_data_157; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_158 = proc_14_io_pipe_phv_out_data_158; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_data_159 = proc_14_io_pipe_phv_out_data_159; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_header_0 = proc_14_io_pipe_phv_out_header_0; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_header_1 = proc_14_io_pipe_phv_out_header_1; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_header_2 = proc_14_io_pipe_phv_out_header_2; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_header_3 = proc_14_io_pipe_phv_out_header_3; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_header_4 = proc_14_io_pipe_phv_out_header_4; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_header_5 = proc_14_io_pipe_phv_out_header_5; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_header_6 = proc_14_io_pipe_phv_out_header_6; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_header_7 = proc_14_io_pipe_phv_out_header_7; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_header_8 = proc_14_io_pipe_phv_out_header_8; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_header_9 = proc_14_io_pipe_phv_out_header_9; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_header_10 = proc_14_io_pipe_phv_out_header_10; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_header_11 = proc_14_io_pipe_phv_out_header_11; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_header_12 = proc_14_io_pipe_phv_out_header_12; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_header_13 = proc_14_io_pipe_phv_out_header_13; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_header_14 = proc_14_io_pipe_phv_out_header_14; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_header_15 = proc_14_io_pipe_phv_out_header_15; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_parse_current_state = proc_14_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_parse_current_offset = proc_14_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_parse_transition_field = proc_14_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_next_processor_id = proc_14_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_next_config_id = proc_14_io_pipe_phv_out_next_config_id; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_valid = proc_14_io_pipe_phv_out_valid; // @[ipsa.scala 82:32]
  assign trans_14_io_pipe_phv_in_last = proc_14_io_pipe_phv_out_last; // @[ipsa.scala 82:32]
  assign trans_14_io_next_proc_exist = 1'h1; // @[ipsa.scala 80:48]
  assign trans_15_clock = clock;
  assign trans_15_io_pipe_phv_in_data_0 = proc_15_io_pipe_phv_out_data_0; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_1 = proc_15_io_pipe_phv_out_data_1; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_2 = proc_15_io_pipe_phv_out_data_2; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_3 = proc_15_io_pipe_phv_out_data_3; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_4 = proc_15_io_pipe_phv_out_data_4; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_5 = proc_15_io_pipe_phv_out_data_5; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_6 = proc_15_io_pipe_phv_out_data_6; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_7 = proc_15_io_pipe_phv_out_data_7; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_8 = proc_15_io_pipe_phv_out_data_8; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_9 = proc_15_io_pipe_phv_out_data_9; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_10 = proc_15_io_pipe_phv_out_data_10; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_11 = proc_15_io_pipe_phv_out_data_11; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_12 = proc_15_io_pipe_phv_out_data_12; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_13 = proc_15_io_pipe_phv_out_data_13; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_14 = proc_15_io_pipe_phv_out_data_14; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_15 = proc_15_io_pipe_phv_out_data_15; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_16 = proc_15_io_pipe_phv_out_data_16; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_17 = proc_15_io_pipe_phv_out_data_17; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_18 = proc_15_io_pipe_phv_out_data_18; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_19 = proc_15_io_pipe_phv_out_data_19; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_20 = proc_15_io_pipe_phv_out_data_20; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_21 = proc_15_io_pipe_phv_out_data_21; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_22 = proc_15_io_pipe_phv_out_data_22; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_23 = proc_15_io_pipe_phv_out_data_23; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_24 = proc_15_io_pipe_phv_out_data_24; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_25 = proc_15_io_pipe_phv_out_data_25; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_26 = proc_15_io_pipe_phv_out_data_26; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_27 = proc_15_io_pipe_phv_out_data_27; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_28 = proc_15_io_pipe_phv_out_data_28; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_29 = proc_15_io_pipe_phv_out_data_29; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_30 = proc_15_io_pipe_phv_out_data_30; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_31 = proc_15_io_pipe_phv_out_data_31; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_32 = proc_15_io_pipe_phv_out_data_32; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_33 = proc_15_io_pipe_phv_out_data_33; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_34 = proc_15_io_pipe_phv_out_data_34; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_35 = proc_15_io_pipe_phv_out_data_35; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_36 = proc_15_io_pipe_phv_out_data_36; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_37 = proc_15_io_pipe_phv_out_data_37; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_38 = proc_15_io_pipe_phv_out_data_38; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_39 = proc_15_io_pipe_phv_out_data_39; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_40 = proc_15_io_pipe_phv_out_data_40; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_41 = proc_15_io_pipe_phv_out_data_41; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_42 = proc_15_io_pipe_phv_out_data_42; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_43 = proc_15_io_pipe_phv_out_data_43; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_44 = proc_15_io_pipe_phv_out_data_44; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_45 = proc_15_io_pipe_phv_out_data_45; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_46 = proc_15_io_pipe_phv_out_data_46; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_47 = proc_15_io_pipe_phv_out_data_47; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_48 = proc_15_io_pipe_phv_out_data_48; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_49 = proc_15_io_pipe_phv_out_data_49; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_50 = proc_15_io_pipe_phv_out_data_50; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_51 = proc_15_io_pipe_phv_out_data_51; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_52 = proc_15_io_pipe_phv_out_data_52; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_53 = proc_15_io_pipe_phv_out_data_53; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_54 = proc_15_io_pipe_phv_out_data_54; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_55 = proc_15_io_pipe_phv_out_data_55; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_56 = proc_15_io_pipe_phv_out_data_56; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_57 = proc_15_io_pipe_phv_out_data_57; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_58 = proc_15_io_pipe_phv_out_data_58; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_59 = proc_15_io_pipe_phv_out_data_59; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_60 = proc_15_io_pipe_phv_out_data_60; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_61 = proc_15_io_pipe_phv_out_data_61; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_62 = proc_15_io_pipe_phv_out_data_62; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_63 = proc_15_io_pipe_phv_out_data_63; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_64 = proc_15_io_pipe_phv_out_data_64; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_65 = proc_15_io_pipe_phv_out_data_65; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_66 = proc_15_io_pipe_phv_out_data_66; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_67 = proc_15_io_pipe_phv_out_data_67; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_68 = proc_15_io_pipe_phv_out_data_68; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_69 = proc_15_io_pipe_phv_out_data_69; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_70 = proc_15_io_pipe_phv_out_data_70; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_71 = proc_15_io_pipe_phv_out_data_71; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_72 = proc_15_io_pipe_phv_out_data_72; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_73 = proc_15_io_pipe_phv_out_data_73; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_74 = proc_15_io_pipe_phv_out_data_74; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_75 = proc_15_io_pipe_phv_out_data_75; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_76 = proc_15_io_pipe_phv_out_data_76; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_77 = proc_15_io_pipe_phv_out_data_77; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_78 = proc_15_io_pipe_phv_out_data_78; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_79 = proc_15_io_pipe_phv_out_data_79; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_80 = proc_15_io_pipe_phv_out_data_80; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_81 = proc_15_io_pipe_phv_out_data_81; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_82 = proc_15_io_pipe_phv_out_data_82; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_83 = proc_15_io_pipe_phv_out_data_83; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_84 = proc_15_io_pipe_phv_out_data_84; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_85 = proc_15_io_pipe_phv_out_data_85; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_86 = proc_15_io_pipe_phv_out_data_86; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_87 = proc_15_io_pipe_phv_out_data_87; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_88 = proc_15_io_pipe_phv_out_data_88; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_89 = proc_15_io_pipe_phv_out_data_89; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_90 = proc_15_io_pipe_phv_out_data_90; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_91 = proc_15_io_pipe_phv_out_data_91; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_92 = proc_15_io_pipe_phv_out_data_92; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_93 = proc_15_io_pipe_phv_out_data_93; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_94 = proc_15_io_pipe_phv_out_data_94; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_95 = proc_15_io_pipe_phv_out_data_95; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_96 = proc_15_io_pipe_phv_out_data_96; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_97 = proc_15_io_pipe_phv_out_data_97; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_98 = proc_15_io_pipe_phv_out_data_98; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_99 = proc_15_io_pipe_phv_out_data_99; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_100 = proc_15_io_pipe_phv_out_data_100; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_101 = proc_15_io_pipe_phv_out_data_101; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_102 = proc_15_io_pipe_phv_out_data_102; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_103 = proc_15_io_pipe_phv_out_data_103; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_104 = proc_15_io_pipe_phv_out_data_104; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_105 = proc_15_io_pipe_phv_out_data_105; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_106 = proc_15_io_pipe_phv_out_data_106; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_107 = proc_15_io_pipe_phv_out_data_107; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_108 = proc_15_io_pipe_phv_out_data_108; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_109 = proc_15_io_pipe_phv_out_data_109; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_110 = proc_15_io_pipe_phv_out_data_110; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_111 = proc_15_io_pipe_phv_out_data_111; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_112 = proc_15_io_pipe_phv_out_data_112; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_113 = proc_15_io_pipe_phv_out_data_113; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_114 = proc_15_io_pipe_phv_out_data_114; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_115 = proc_15_io_pipe_phv_out_data_115; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_116 = proc_15_io_pipe_phv_out_data_116; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_117 = proc_15_io_pipe_phv_out_data_117; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_118 = proc_15_io_pipe_phv_out_data_118; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_119 = proc_15_io_pipe_phv_out_data_119; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_120 = proc_15_io_pipe_phv_out_data_120; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_121 = proc_15_io_pipe_phv_out_data_121; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_122 = proc_15_io_pipe_phv_out_data_122; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_123 = proc_15_io_pipe_phv_out_data_123; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_124 = proc_15_io_pipe_phv_out_data_124; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_125 = proc_15_io_pipe_phv_out_data_125; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_126 = proc_15_io_pipe_phv_out_data_126; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_127 = proc_15_io_pipe_phv_out_data_127; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_128 = proc_15_io_pipe_phv_out_data_128; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_129 = proc_15_io_pipe_phv_out_data_129; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_130 = proc_15_io_pipe_phv_out_data_130; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_131 = proc_15_io_pipe_phv_out_data_131; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_132 = proc_15_io_pipe_phv_out_data_132; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_133 = proc_15_io_pipe_phv_out_data_133; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_134 = proc_15_io_pipe_phv_out_data_134; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_135 = proc_15_io_pipe_phv_out_data_135; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_136 = proc_15_io_pipe_phv_out_data_136; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_137 = proc_15_io_pipe_phv_out_data_137; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_138 = proc_15_io_pipe_phv_out_data_138; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_139 = proc_15_io_pipe_phv_out_data_139; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_140 = proc_15_io_pipe_phv_out_data_140; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_141 = proc_15_io_pipe_phv_out_data_141; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_142 = proc_15_io_pipe_phv_out_data_142; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_143 = proc_15_io_pipe_phv_out_data_143; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_144 = proc_15_io_pipe_phv_out_data_144; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_145 = proc_15_io_pipe_phv_out_data_145; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_146 = proc_15_io_pipe_phv_out_data_146; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_147 = proc_15_io_pipe_phv_out_data_147; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_148 = proc_15_io_pipe_phv_out_data_148; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_149 = proc_15_io_pipe_phv_out_data_149; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_150 = proc_15_io_pipe_phv_out_data_150; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_151 = proc_15_io_pipe_phv_out_data_151; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_152 = proc_15_io_pipe_phv_out_data_152; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_153 = proc_15_io_pipe_phv_out_data_153; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_154 = proc_15_io_pipe_phv_out_data_154; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_155 = proc_15_io_pipe_phv_out_data_155; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_156 = proc_15_io_pipe_phv_out_data_156; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_157 = proc_15_io_pipe_phv_out_data_157; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_158 = proc_15_io_pipe_phv_out_data_158; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_data_159 = proc_15_io_pipe_phv_out_data_159; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_header_0 = proc_15_io_pipe_phv_out_header_0; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_header_1 = proc_15_io_pipe_phv_out_header_1; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_header_2 = proc_15_io_pipe_phv_out_header_2; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_header_3 = proc_15_io_pipe_phv_out_header_3; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_header_4 = proc_15_io_pipe_phv_out_header_4; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_header_5 = proc_15_io_pipe_phv_out_header_5; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_header_6 = proc_15_io_pipe_phv_out_header_6; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_header_7 = proc_15_io_pipe_phv_out_header_7; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_header_8 = proc_15_io_pipe_phv_out_header_8; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_header_9 = proc_15_io_pipe_phv_out_header_9; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_header_10 = proc_15_io_pipe_phv_out_header_10; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_header_11 = proc_15_io_pipe_phv_out_header_11; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_header_12 = proc_15_io_pipe_phv_out_header_12; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_header_13 = proc_15_io_pipe_phv_out_header_13; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_header_14 = proc_15_io_pipe_phv_out_header_14; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_header_15 = proc_15_io_pipe_phv_out_header_15; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_parse_current_state = proc_15_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_parse_current_offset = proc_15_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_parse_transition_field = proc_15_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_next_processor_id = proc_15_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_next_config_id = proc_15_io_pipe_phv_out_next_config_id; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_valid = proc_15_io_pipe_phv_out_valid; // @[ipsa.scala 82:32]
  assign trans_15_io_pipe_phv_in_last = proc_15_io_pipe_phv_out_last; // @[ipsa.scala 82:32]
  assign trans_15_io_next_proc_exist = 1'h1; // @[ipsa.scala 80:48]
endmodule
