module PrimitiveWriteBack(
  input         clock,
  input  [7:0]  io_pipe_phv_in_data_0,
  input  [7:0]  io_pipe_phv_in_data_1,
  input  [7:0]  io_pipe_phv_in_data_2,
  input  [7:0]  io_pipe_phv_in_data_3,
  input  [7:0]  io_pipe_phv_in_data_4,
  input  [7:0]  io_pipe_phv_in_data_5,
  input  [7:0]  io_pipe_phv_in_data_6,
  input  [7:0]  io_pipe_phv_in_data_7,
  input  [7:0]  io_pipe_phv_in_data_8,
  input  [7:0]  io_pipe_phv_in_data_9,
  input  [7:0]  io_pipe_phv_in_data_10,
  input  [7:0]  io_pipe_phv_in_data_11,
  input  [7:0]  io_pipe_phv_in_data_12,
  input  [7:0]  io_pipe_phv_in_data_13,
  input  [7:0]  io_pipe_phv_in_data_14,
  input  [7:0]  io_pipe_phv_in_data_15,
  input  [7:0]  io_pipe_phv_in_data_16,
  input  [7:0]  io_pipe_phv_in_data_17,
  input  [7:0]  io_pipe_phv_in_data_18,
  input  [7:0]  io_pipe_phv_in_data_19,
  input  [7:0]  io_pipe_phv_in_data_20,
  input  [7:0]  io_pipe_phv_in_data_21,
  input  [7:0]  io_pipe_phv_in_data_22,
  input  [7:0]  io_pipe_phv_in_data_23,
  input  [7:0]  io_pipe_phv_in_data_24,
  input  [7:0]  io_pipe_phv_in_data_25,
  input  [7:0]  io_pipe_phv_in_data_26,
  input  [7:0]  io_pipe_phv_in_data_27,
  input  [7:0]  io_pipe_phv_in_data_28,
  input  [7:0]  io_pipe_phv_in_data_29,
  input  [7:0]  io_pipe_phv_in_data_30,
  input  [7:0]  io_pipe_phv_in_data_31,
  input  [7:0]  io_pipe_phv_in_data_32,
  input  [7:0]  io_pipe_phv_in_data_33,
  input  [7:0]  io_pipe_phv_in_data_34,
  input  [7:0]  io_pipe_phv_in_data_35,
  input  [7:0]  io_pipe_phv_in_data_36,
  input  [7:0]  io_pipe_phv_in_data_37,
  input  [7:0]  io_pipe_phv_in_data_38,
  input  [7:0]  io_pipe_phv_in_data_39,
  input  [7:0]  io_pipe_phv_in_data_40,
  input  [7:0]  io_pipe_phv_in_data_41,
  input  [7:0]  io_pipe_phv_in_data_42,
  input  [7:0]  io_pipe_phv_in_data_43,
  input  [7:0]  io_pipe_phv_in_data_44,
  input  [7:0]  io_pipe_phv_in_data_45,
  input  [7:0]  io_pipe_phv_in_data_46,
  input  [7:0]  io_pipe_phv_in_data_47,
  input  [7:0]  io_pipe_phv_in_data_48,
  input  [7:0]  io_pipe_phv_in_data_49,
  input  [7:0]  io_pipe_phv_in_data_50,
  input  [7:0]  io_pipe_phv_in_data_51,
  input  [7:0]  io_pipe_phv_in_data_52,
  input  [7:0]  io_pipe_phv_in_data_53,
  input  [7:0]  io_pipe_phv_in_data_54,
  input  [7:0]  io_pipe_phv_in_data_55,
  input  [7:0]  io_pipe_phv_in_data_56,
  input  [7:0]  io_pipe_phv_in_data_57,
  input  [7:0]  io_pipe_phv_in_data_58,
  input  [7:0]  io_pipe_phv_in_data_59,
  input  [7:0]  io_pipe_phv_in_data_60,
  input  [7:0]  io_pipe_phv_in_data_61,
  input  [7:0]  io_pipe_phv_in_data_62,
  input  [7:0]  io_pipe_phv_in_data_63,
  input  [7:0]  io_pipe_phv_in_data_64,
  input  [7:0]  io_pipe_phv_in_data_65,
  input  [7:0]  io_pipe_phv_in_data_66,
  input  [7:0]  io_pipe_phv_in_data_67,
  input  [7:0]  io_pipe_phv_in_data_68,
  input  [7:0]  io_pipe_phv_in_data_69,
  input  [7:0]  io_pipe_phv_in_data_70,
  input  [7:0]  io_pipe_phv_in_data_71,
  input  [7:0]  io_pipe_phv_in_data_72,
  input  [7:0]  io_pipe_phv_in_data_73,
  input  [7:0]  io_pipe_phv_in_data_74,
  input  [7:0]  io_pipe_phv_in_data_75,
  input  [7:0]  io_pipe_phv_in_data_76,
  input  [7:0]  io_pipe_phv_in_data_77,
  input  [7:0]  io_pipe_phv_in_data_78,
  input  [7:0]  io_pipe_phv_in_data_79,
  input  [7:0]  io_pipe_phv_in_data_80,
  input  [7:0]  io_pipe_phv_in_data_81,
  input  [7:0]  io_pipe_phv_in_data_82,
  input  [7:0]  io_pipe_phv_in_data_83,
  input  [7:0]  io_pipe_phv_in_data_84,
  input  [7:0]  io_pipe_phv_in_data_85,
  input  [7:0]  io_pipe_phv_in_data_86,
  input  [7:0]  io_pipe_phv_in_data_87,
  input  [7:0]  io_pipe_phv_in_data_88,
  input  [7:0]  io_pipe_phv_in_data_89,
  input  [7:0]  io_pipe_phv_in_data_90,
  input  [7:0]  io_pipe_phv_in_data_91,
  input  [7:0]  io_pipe_phv_in_data_92,
  input  [7:0]  io_pipe_phv_in_data_93,
  input  [7:0]  io_pipe_phv_in_data_94,
  input  [7:0]  io_pipe_phv_in_data_95,
  input  [7:0]  io_pipe_phv_in_data_96,
  input  [7:0]  io_pipe_phv_in_data_97,
  input  [7:0]  io_pipe_phv_in_data_98,
  input  [7:0]  io_pipe_phv_in_data_99,
  input  [7:0]  io_pipe_phv_in_data_100,
  input  [7:0]  io_pipe_phv_in_data_101,
  input  [7:0]  io_pipe_phv_in_data_102,
  input  [7:0]  io_pipe_phv_in_data_103,
  input  [7:0]  io_pipe_phv_in_data_104,
  input  [7:0]  io_pipe_phv_in_data_105,
  input  [7:0]  io_pipe_phv_in_data_106,
  input  [7:0]  io_pipe_phv_in_data_107,
  input  [7:0]  io_pipe_phv_in_data_108,
  input  [7:0]  io_pipe_phv_in_data_109,
  input  [7:0]  io_pipe_phv_in_data_110,
  input  [7:0]  io_pipe_phv_in_data_111,
  input  [7:0]  io_pipe_phv_in_data_112,
  input  [7:0]  io_pipe_phv_in_data_113,
  input  [7:0]  io_pipe_phv_in_data_114,
  input  [7:0]  io_pipe_phv_in_data_115,
  input  [7:0]  io_pipe_phv_in_data_116,
  input  [7:0]  io_pipe_phv_in_data_117,
  input  [7:0]  io_pipe_phv_in_data_118,
  input  [7:0]  io_pipe_phv_in_data_119,
  input  [7:0]  io_pipe_phv_in_data_120,
  input  [7:0]  io_pipe_phv_in_data_121,
  input  [7:0]  io_pipe_phv_in_data_122,
  input  [7:0]  io_pipe_phv_in_data_123,
  input  [7:0]  io_pipe_phv_in_data_124,
  input  [7:0]  io_pipe_phv_in_data_125,
  input  [7:0]  io_pipe_phv_in_data_126,
  input  [7:0]  io_pipe_phv_in_data_127,
  input  [7:0]  io_pipe_phv_in_data_128,
  input  [7:0]  io_pipe_phv_in_data_129,
  input  [7:0]  io_pipe_phv_in_data_130,
  input  [7:0]  io_pipe_phv_in_data_131,
  input  [7:0]  io_pipe_phv_in_data_132,
  input  [7:0]  io_pipe_phv_in_data_133,
  input  [7:0]  io_pipe_phv_in_data_134,
  input  [7:0]  io_pipe_phv_in_data_135,
  input  [7:0]  io_pipe_phv_in_data_136,
  input  [7:0]  io_pipe_phv_in_data_137,
  input  [7:0]  io_pipe_phv_in_data_138,
  input  [7:0]  io_pipe_phv_in_data_139,
  input  [7:0]  io_pipe_phv_in_data_140,
  input  [7:0]  io_pipe_phv_in_data_141,
  input  [7:0]  io_pipe_phv_in_data_142,
  input  [7:0]  io_pipe_phv_in_data_143,
  input  [7:0]  io_pipe_phv_in_data_144,
  input  [7:0]  io_pipe_phv_in_data_145,
  input  [7:0]  io_pipe_phv_in_data_146,
  input  [7:0]  io_pipe_phv_in_data_147,
  input  [7:0]  io_pipe_phv_in_data_148,
  input  [7:0]  io_pipe_phv_in_data_149,
  input  [7:0]  io_pipe_phv_in_data_150,
  input  [7:0]  io_pipe_phv_in_data_151,
  input  [7:0]  io_pipe_phv_in_data_152,
  input  [7:0]  io_pipe_phv_in_data_153,
  input  [7:0]  io_pipe_phv_in_data_154,
  input  [7:0]  io_pipe_phv_in_data_155,
  input  [7:0]  io_pipe_phv_in_data_156,
  input  [7:0]  io_pipe_phv_in_data_157,
  input  [7:0]  io_pipe_phv_in_data_158,
  input  [7:0]  io_pipe_phv_in_data_159,
  input  [15:0] io_pipe_phv_in_header_0,
  input  [15:0] io_pipe_phv_in_header_1,
  input  [15:0] io_pipe_phv_in_header_2,
  input  [15:0] io_pipe_phv_in_header_3,
  input  [15:0] io_pipe_phv_in_header_4,
  input  [15:0] io_pipe_phv_in_header_5,
  input  [15:0] io_pipe_phv_in_header_6,
  input  [15:0] io_pipe_phv_in_header_7,
  input  [15:0] io_pipe_phv_in_header_8,
  input  [15:0] io_pipe_phv_in_header_9,
  input  [15:0] io_pipe_phv_in_header_10,
  input  [15:0] io_pipe_phv_in_header_11,
  input  [15:0] io_pipe_phv_in_header_12,
  input  [15:0] io_pipe_phv_in_header_13,
  input  [15:0] io_pipe_phv_in_header_14,
  input  [15:0] io_pipe_phv_in_header_15,
  input  [7:0]  io_pipe_phv_in_parse_current_state,
  input  [7:0]  io_pipe_phv_in_parse_current_offset,
  input  [15:0] io_pipe_phv_in_parse_transition_field,
  input  [3:0]  io_pipe_phv_in_next_processor_id,
  input         io_pipe_phv_in_next_config_id,
  input         io_pipe_phv_in_is_valid_processor,
  input         io_pipe_phv_in_valid,
  output [7:0]  io_pipe_phv_out_data_0,
  output [7:0]  io_pipe_phv_out_data_1,
  output [7:0]  io_pipe_phv_out_data_2,
  output [7:0]  io_pipe_phv_out_data_3,
  output [7:0]  io_pipe_phv_out_data_4,
  output [7:0]  io_pipe_phv_out_data_5,
  output [7:0]  io_pipe_phv_out_data_6,
  output [7:0]  io_pipe_phv_out_data_7,
  output [7:0]  io_pipe_phv_out_data_8,
  output [7:0]  io_pipe_phv_out_data_9,
  output [7:0]  io_pipe_phv_out_data_10,
  output [7:0]  io_pipe_phv_out_data_11,
  output [7:0]  io_pipe_phv_out_data_12,
  output [7:0]  io_pipe_phv_out_data_13,
  output [7:0]  io_pipe_phv_out_data_14,
  output [7:0]  io_pipe_phv_out_data_15,
  output [7:0]  io_pipe_phv_out_data_16,
  output [7:0]  io_pipe_phv_out_data_17,
  output [7:0]  io_pipe_phv_out_data_18,
  output [7:0]  io_pipe_phv_out_data_19,
  output [7:0]  io_pipe_phv_out_data_20,
  output [7:0]  io_pipe_phv_out_data_21,
  output [7:0]  io_pipe_phv_out_data_22,
  output [7:0]  io_pipe_phv_out_data_23,
  output [7:0]  io_pipe_phv_out_data_24,
  output [7:0]  io_pipe_phv_out_data_25,
  output [7:0]  io_pipe_phv_out_data_26,
  output [7:0]  io_pipe_phv_out_data_27,
  output [7:0]  io_pipe_phv_out_data_28,
  output [7:0]  io_pipe_phv_out_data_29,
  output [7:0]  io_pipe_phv_out_data_30,
  output [7:0]  io_pipe_phv_out_data_31,
  output [7:0]  io_pipe_phv_out_data_32,
  output [7:0]  io_pipe_phv_out_data_33,
  output [7:0]  io_pipe_phv_out_data_34,
  output [7:0]  io_pipe_phv_out_data_35,
  output [7:0]  io_pipe_phv_out_data_36,
  output [7:0]  io_pipe_phv_out_data_37,
  output [7:0]  io_pipe_phv_out_data_38,
  output [7:0]  io_pipe_phv_out_data_39,
  output [7:0]  io_pipe_phv_out_data_40,
  output [7:0]  io_pipe_phv_out_data_41,
  output [7:0]  io_pipe_phv_out_data_42,
  output [7:0]  io_pipe_phv_out_data_43,
  output [7:0]  io_pipe_phv_out_data_44,
  output [7:0]  io_pipe_phv_out_data_45,
  output [7:0]  io_pipe_phv_out_data_46,
  output [7:0]  io_pipe_phv_out_data_47,
  output [7:0]  io_pipe_phv_out_data_48,
  output [7:0]  io_pipe_phv_out_data_49,
  output [7:0]  io_pipe_phv_out_data_50,
  output [7:0]  io_pipe_phv_out_data_51,
  output [7:0]  io_pipe_phv_out_data_52,
  output [7:0]  io_pipe_phv_out_data_53,
  output [7:0]  io_pipe_phv_out_data_54,
  output [7:0]  io_pipe_phv_out_data_55,
  output [7:0]  io_pipe_phv_out_data_56,
  output [7:0]  io_pipe_phv_out_data_57,
  output [7:0]  io_pipe_phv_out_data_58,
  output [7:0]  io_pipe_phv_out_data_59,
  output [7:0]  io_pipe_phv_out_data_60,
  output [7:0]  io_pipe_phv_out_data_61,
  output [7:0]  io_pipe_phv_out_data_62,
  output [7:0]  io_pipe_phv_out_data_63,
  output [7:0]  io_pipe_phv_out_data_64,
  output [7:0]  io_pipe_phv_out_data_65,
  output [7:0]  io_pipe_phv_out_data_66,
  output [7:0]  io_pipe_phv_out_data_67,
  output [7:0]  io_pipe_phv_out_data_68,
  output [7:0]  io_pipe_phv_out_data_69,
  output [7:0]  io_pipe_phv_out_data_70,
  output [7:0]  io_pipe_phv_out_data_71,
  output [7:0]  io_pipe_phv_out_data_72,
  output [7:0]  io_pipe_phv_out_data_73,
  output [7:0]  io_pipe_phv_out_data_74,
  output [7:0]  io_pipe_phv_out_data_75,
  output [7:0]  io_pipe_phv_out_data_76,
  output [7:0]  io_pipe_phv_out_data_77,
  output [7:0]  io_pipe_phv_out_data_78,
  output [7:0]  io_pipe_phv_out_data_79,
  output [7:0]  io_pipe_phv_out_data_80,
  output [7:0]  io_pipe_phv_out_data_81,
  output [7:0]  io_pipe_phv_out_data_82,
  output [7:0]  io_pipe_phv_out_data_83,
  output [7:0]  io_pipe_phv_out_data_84,
  output [7:0]  io_pipe_phv_out_data_85,
  output [7:0]  io_pipe_phv_out_data_86,
  output [7:0]  io_pipe_phv_out_data_87,
  output [7:0]  io_pipe_phv_out_data_88,
  output [7:0]  io_pipe_phv_out_data_89,
  output [7:0]  io_pipe_phv_out_data_90,
  output [7:0]  io_pipe_phv_out_data_91,
  output [7:0]  io_pipe_phv_out_data_92,
  output [7:0]  io_pipe_phv_out_data_93,
  output [7:0]  io_pipe_phv_out_data_94,
  output [7:0]  io_pipe_phv_out_data_95,
  output [7:0]  io_pipe_phv_out_data_96,
  output [7:0]  io_pipe_phv_out_data_97,
  output [7:0]  io_pipe_phv_out_data_98,
  output [7:0]  io_pipe_phv_out_data_99,
  output [7:0]  io_pipe_phv_out_data_100,
  output [7:0]  io_pipe_phv_out_data_101,
  output [7:0]  io_pipe_phv_out_data_102,
  output [7:0]  io_pipe_phv_out_data_103,
  output [7:0]  io_pipe_phv_out_data_104,
  output [7:0]  io_pipe_phv_out_data_105,
  output [7:0]  io_pipe_phv_out_data_106,
  output [7:0]  io_pipe_phv_out_data_107,
  output [7:0]  io_pipe_phv_out_data_108,
  output [7:0]  io_pipe_phv_out_data_109,
  output [7:0]  io_pipe_phv_out_data_110,
  output [7:0]  io_pipe_phv_out_data_111,
  output [7:0]  io_pipe_phv_out_data_112,
  output [7:0]  io_pipe_phv_out_data_113,
  output [7:0]  io_pipe_phv_out_data_114,
  output [7:0]  io_pipe_phv_out_data_115,
  output [7:0]  io_pipe_phv_out_data_116,
  output [7:0]  io_pipe_phv_out_data_117,
  output [7:0]  io_pipe_phv_out_data_118,
  output [7:0]  io_pipe_phv_out_data_119,
  output [7:0]  io_pipe_phv_out_data_120,
  output [7:0]  io_pipe_phv_out_data_121,
  output [7:0]  io_pipe_phv_out_data_122,
  output [7:0]  io_pipe_phv_out_data_123,
  output [7:0]  io_pipe_phv_out_data_124,
  output [7:0]  io_pipe_phv_out_data_125,
  output [7:0]  io_pipe_phv_out_data_126,
  output [7:0]  io_pipe_phv_out_data_127,
  output [7:0]  io_pipe_phv_out_data_128,
  output [7:0]  io_pipe_phv_out_data_129,
  output [7:0]  io_pipe_phv_out_data_130,
  output [7:0]  io_pipe_phv_out_data_131,
  output [7:0]  io_pipe_phv_out_data_132,
  output [7:0]  io_pipe_phv_out_data_133,
  output [7:0]  io_pipe_phv_out_data_134,
  output [7:0]  io_pipe_phv_out_data_135,
  output [7:0]  io_pipe_phv_out_data_136,
  output [7:0]  io_pipe_phv_out_data_137,
  output [7:0]  io_pipe_phv_out_data_138,
  output [7:0]  io_pipe_phv_out_data_139,
  output [7:0]  io_pipe_phv_out_data_140,
  output [7:0]  io_pipe_phv_out_data_141,
  output [7:0]  io_pipe_phv_out_data_142,
  output [7:0]  io_pipe_phv_out_data_143,
  output [7:0]  io_pipe_phv_out_data_144,
  output [7:0]  io_pipe_phv_out_data_145,
  output [7:0]  io_pipe_phv_out_data_146,
  output [7:0]  io_pipe_phv_out_data_147,
  output [7:0]  io_pipe_phv_out_data_148,
  output [7:0]  io_pipe_phv_out_data_149,
  output [7:0]  io_pipe_phv_out_data_150,
  output [7:0]  io_pipe_phv_out_data_151,
  output [7:0]  io_pipe_phv_out_data_152,
  output [7:0]  io_pipe_phv_out_data_153,
  output [7:0]  io_pipe_phv_out_data_154,
  output [7:0]  io_pipe_phv_out_data_155,
  output [7:0]  io_pipe_phv_out_data_156,
  output [7:0]  io_pipe_phv_out_data_157,
  output [7:0]  io_pipe_phv_out_data_158,
  output [7:0]  io_pipe_phv_out_data_159,
  output [15:0] io_pipe_phv_out_header_0,
  output [15:0] io_pipe_phv_out_header_1,
  output [15:0] io_pipe_phv_out_header_2,
  output [15:0] io_pipe_phv_out_header_3,
  output [15:0] io_pipe_phv_out_header_4,
  output [15:0] io_pipe_phv_out_header_5,
  output [15:0] io_pipe_phv_out_header_6,
  output [15:0] io_pipe_phv_out_header_7,
  output [15:0] io_pipe_phv_out_header_8,
  output [15:0] io_pipe_phv_out_header_9,
  output [15:0] io_pipe_phv_out_header_10,
  output [15:0] io_pipe_phv_out_header_11,
  output [15:0] io_pipe_phv_out_header_12,
  output [15:0] io_pipe_phv_out_header_13,
  output [15:0] io_pipe_phv_out_header_14,
  output [15:0] io_pipe_phv_out_header_15,
  output [7:0]  io_pipe_phv_out_parse_current_state,
  output [7:0]  io_pipe_phv_out_parse_current_offset,
  output [15:0] io_pipe_phv_out_parse_transition_field,
  output [3:0]  io_pipe_phv_out_next_processor_id,
  output        io_pipe_phv_out_next_config_id,
  output        io_pipe_phv_out_valid,
  input  [31:0] io_vliw_in_0,
  input  [31:0] io_vliw_in_1,
  input  [31:0] io_vliw_in_2,
  input  [31:0] io_vliw_in_3,
  input  [31:0] io_field_in_0,
  input  [31:0] io_field_in_1,
  input  [31:0] io_field_in_2,
  input  [31:0] io_field_in_3,
  input  [3:0]  io_mask_in_0,
  input  [3:0]  io_mask_in_1,
  input  [3:0]  io_mask_in_2,
  input  [3:0]  io_mask_in_3,
  input  [5:0]  io_dst_offset_in_0,
  input  [5:0]  io_dst_offset_in_1,
  input  [5:0]  io_dst_offset_in_2,
  input  [5:0]  io_dst_offset_in_3
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] phv_data_0; // @[executor.scala 448:22]
  reg [7:0] phv_data_1; // @[executor.scala 448:22]
  reg [7:0] phv_data_2; // @[executor.scala 448:22]
  reg [7:0] phv_data_3; // @[executor.scala 448:22]
  reg [7:0] phv_data_4; // @[executor.scala 448:22]
  reg [7:0] phv_data_5; // @[executor.scala 448:22]
  reg [7:0] phv_data_6; // @[executor.scala 448:22]
  reg [7:0] phv_data_7; // @[executor.scala 448:22]
  reg [7:0] phv_data_8; // @[executor.scala 448:22]
  reg [7:0] phv_data_9; // @[executor.scala 448:22]
  reg [7:0] phv_data_10; // @[executor.scala 448:22]
  reg [7:0] phv_data_11; // @[executor.scala 448:22]
  reg [7:0] phv_data_12; // @[executor.scala 448:22]
  reg [7:0] phv_data_13; // @[executor.scala 448:22]
  reg [7:0] phv_data_14; // @[executor.scala 448:22]
  reg [7:0] phv_data_15; // @[executor.scala 448:22]
  reg [7:0] phv_data_16; // @[executor.scala 448:22]
  reg [7:0] phv_data_17; // @[executor.scala 448:22]
  reg [7:0] phv_data_18; // @[executor.scala 448:22]
  reg [7:0] phv_data_19; // @[executor.scala 448:22]
  reg [7:0] phv_data_20; // @[executor.scala 448:22]
  reg [7:0] phv_data_21; // @[executor.scala 448:22]
  reg [7:0] phv_data_22; // @[executor.scala 448:22]
  reg [7:0] phv_data_23; // @[executor.scala 448:22]
  reg [7:0] phv_data_24; // @[executor.scala 448:22]
  reg [7:0] phv_data_25; // @[executor.scala 448:22]
  reg [7:0] phv_data_26; // @[executor.scala 448:22]
  reg [7:0] phv_data_27; // @[executor.scala 448:22]
  reg [7:0] phv_data_28; // @[executor.scala 448:22]
  reg [7:0] phv_data_29; // @[executor.scala 448:22]
  reg [7:0] phv_data_30; // @[executor.scala 448:22]
  reg [7:0] phv_data_31; // @[executor.scala 448:22]
  reg [7:0] phv_data_32; // @[executor.scala 448:22]
  reg [7:0] phv_data_33; // @[executor.scala 448:22]
  reg [7:0] phv_data_34; // @[executor.scala 448:22]
  reg [7:0] phv_data_35; // @[executor.scala 448:22]
  reg [7:0] phv_data_36; // @[executor.scala 448:22]
  reg [7:0] phv_data_37; // @[executor.scala 448:22]
  reg [7:0] phv_data_38; // @[executor.scala 448:22]
  reg [7:0] phv_data_39; // @[executor.scala 448:22]
  reg [7:0] phv_data_40; // @[executor.scala 448:22]
  reg [7:0] phv_data_41; // @[executor.scala 448:22]
  reg [7:0] phv_data_42; // @[executor.scala 448:22]
  reg [7:0] phv_data_43; // @[executor.scala 448:22]
  reg [7:0] phv_data_44; // @[executor.scala 448:22]
  reg [7:0] phv_data_45; // @[executor.scala 448:22]
  reg [7:0] phv_data_46; // @[executor.scala 448:22]
  reg [7:0] phv_data_47; // @[executor.scala 448:22]
  reg [7:0] phv_data_48; // @[executor.scala 448:22]
  reg [7:0] phv_data_49; // @[executor.scala 448:22]
  reg [7:0] phv_data_50; // @[executor.scala 448:22]
  reg [7:0] phv_data_51; // @[executor.scala 448:22]
  reg [7:0] phv_data_52; // @[executor.scala 448:22]
  reg [7:0] phv_data_53; // @[executor.scala 448:22]
  reg [7:0] phv_data_54; // @[executor.scala 448:22]
  reg [7:0] phv_data_55; // @[executor.scala 448:22]
  reg [7:0] phv_data_56; // @[executor.scala 448:22]
  reg [7:0] phv_data_57; // @[executor.scala 448:22]
  reg [7:0] phv_data_58; // @[executor.scala 448:22]
  reg [7:0] phv_data_59; // @[executor.scala 448:22]
  reg [7:0] phv_data_60; // @[executor.scala 448:22]
  reg [7:0] phv_data_61; // @[executor.scala 448:22]
  reg [7:0] phv_data_62; // @[executor.scala 448:22]
  reg [7:0] phv_data_63; // @[executor.scala 448:22]
  reg [7:0] phv_data_64; // @[executor.scala 448:22]
  reg [7:0] phv_data_65; // @[executor.scala 448:22]
  reg [7:0] phv_data_66; // @[executor.scala 448:22]
  reg [7:0] phv_data_67; // @[executor.scala 448:22]
  reg [7:0] phv_data_68; // @[executor.scala 448:22]
  reg [7:0] phv_data_69; // @[executor.scala 448:22]
  reg [7:0] phv_data_70; // @[executor.scala 448:22]
  reg [7:0] phv_data_71; // @[executor.scala 448:22]
  reg [7:0] phv_data_72; // @[executor.scala 448:22]
  reg [7:0] phv_data_73; // @[executor.scala 448:22]
  reg [7:0] phv_data_74; // @[executor.scala 448:22]
  reg [7:0] phv_data_75; // @[executor.scala 448:22]
  reg [7:0] phv_data_76; // @[executor.scala 448:22]
  reg [7:0] phv_data_77; // @[executor.scala 448:22]
  reg [7:0] phv_data_78; // @[executor.scala 448:22]
  reg [7:0] phv_data_79; // @[executor.scala 448:22]
  reg [7:0] phv_data_80; // @[executor.scala 448:22]
  reg [7:0] phv_data_81; // @[executor.scala 448:22]
  reg [7:0] phv_data_82; // @[executor.scala 448:22]
  reg [7:0] phv_data_83; // @[executor.scala 448:22]
  reg [7:0] phv_data_84; // @[executor.scala 448:22]
  reg [7:0] phv_data_85; // @[executor.scala 448:22]
  reg [7:0] phv_data_86; // @[executor.scala 448:22]
  reg [7:0] phv_data_87; // @[executor.scala 448:22]
  reg [7:0] phv_data_88; // @[executor.scala 448:22]
  reg [7:0] phv_data_89; // @[executor.scala 448:22]
  reg [7:0] phv_data_90; // @[executor.scala 448:22]
  reg [7:0] phv_data_91; // @[executor.scala 448:22]
  reg [7:0] phv_data_92; // @[executor.scala 448:22]
  reg [7:0] phv_data_93; // @[executor.scala 448:22]
  reg [7:0] phv_data_94; // @[executor.scala 448:22]
  reg [7:0] phv_data_95; // @[executor.scala 448:22]
  reg [7:0] phv_data_96; // @[executor.scala 448:22]
  reg [7:0] phv_data_97; // @[executor.scala 448:22]
  reg [7:0] phv_data_98; // @[executor.scala 448:22]
  reg [7:0] phv_data_99; // @[executor.scala 448:22]
  reg [7:0] phv_data_100; // @[executor.scala 448:22]
  reg [7:0] phv_data_101; // @[executor.scala 448:22]
  reg [7:0] phv_data_102; // @[executor.scala 448:22]
  reg [7:0] phv_data_103; // @[executor.scala 448:22]
  reg [7:0] phv_data_104; // @[executor.scala 448:22]
  reg [7:0] phv_data_105; // @[executor.scala 448:22]
  reg [7:0] phv_data_106; // @[executor.scala 448:22]
  reg [7:0] phv_data_107; // @[executor.scala 448:22]
  reg [7:0] phv_data_108; // @[executor.scala 448:22]
  reg [7:0] phv_data_109; // @[executor.scala 448:22]
  reg [7:0] phv_data_110; // @[executor.scala 448:22]
  reg [7:0] phv_data_111; // @[executor.scala 448:22]
  reg [7:0] phv_data_112; // @[executor.scala 448:22]
  reg [7:0] phv_data_113; // @[executor.scala 448:22]
  reg [7:0] phv_data_114; // @[executor.scala 448:22]
  reg [7:0] phv_data_115; // @[executor.scala 448:22]
  reg [7:0] phv_data_116; // @[executor.scala 448:22]
  reg [7:0] phv_data_117; // @[executor.scala 448:22]
  reg [7:0] phv_data_118; // @[executor.scala 448:22]
  reg [7:0] phv_data_119; // @[executor.scala 448:22]
  reg [7:0] phv_data_120; // @[executor.scala 448:22]
  reg [7:0] phv_data_121; // @[executor.scala 448:22]
  reg [7:0] phv_data_122; // @[executor.scala 448:22]
  reg [7:0] phv_data_123; // @[executor.scala 448:22]
  reg [7:0] phv_data_124; // @[executor.scala 448:22]
  reg [7:0] phv_data_125; // @[executor.scala 448:22]
  reg [7:0] phv_data_126; // @[executor.scala 448:22]
  reg [7:0] phv_data_127; // @[executor.scala 448:22]
  reg [7:0] phv_data_128; // @[executor.scala 448:22]
  reg [7:0] phv_data_129; // @[executor.scala 448:22]
  reg [7:0] phv_data_130; // @[executor.scala 448:22]
  reg [7:0] phv_data_131; // @[executor.scala 448:22]
  reg [7:0] phv_data_132; // @[executor.scala 448:22]
  reg [7:0] phv_data_133; // @[executor.scala 448:22]
  reg [7:0] phv_data_134; // @[executor.scala 448:22]
  reg [7:0] phv_data_135; // @[executor.scala 448:22]
  reg [7:0] phv_data_136; // @[executor.scala 448:22]
  reg [7:0] phv_data_137; // @[executor.scala 448:22]
  reg [7:0] phv_data_138; // @[executor.scala 448:22]
  reg [7:0] phv_data_139; // @[executor.scala 448:22]
  reg [7:0] phv_data_140; // @[executor.scala 448:22]
  reg [7:0] phv_data_141; // @[executor.scala 448:22]
  reg [7:0] phv_data_142; // @[executor.scala 448:22]
  reg [7:0] phv_data_143; // @[executor.scala 448:22]
  reg [7:0] phv_data_144; // @[executor.scala 448:22]
  reg [7:0] phv_data_145; // @[executor.scala 448:22]
  reg [7:0] phv_data_146; // @[executor.scala 448:22]
  reg [7:0] phv_data_147; // @[executor.scala 448:22]
  reg [7:0] phv_data_148; // @[executor.scala 448:22]
  reg [7:0] phv_data_149; // @[executor.scala 448:22]
  reg [7:0] phv_data_150; // @[executor.scala 448:22]
  reg [7:0] phv_data_151; // @[executor.scala 448:22]
  reg [7:0] phv_data_152; // @[executor.scala 448:22]
  reg [7:0] phv_data_153; // @[executor.scala 448:22]
  reg [7:0] phv_data_154; // @[executor.scala 448:22]
  reg [7:0] phv_data_155; // @[executor.scala 448:22]
  reg [7:0] phv_data_156; // @[executor.scala 448:22]
  reg [7:0] phv_data_157; // @[executor.scala 448:22]
  reg [7:0] phv_data_158; // @[executor.scala 448:22]
  reg [7:0] phv_data_159; // @[executor.scala 448:22]
  reg [15:0] phv_header_0; // @[executor.scala 448:22]
  reg [15:0] phv_header_1; // @[executor.scala 448:22]
  reg [15:0] phv_header_2; // @[executor.scala 448:22]
  reg [15:0] phv_header_3; // @[executor.scala 448:22]
  reg [15:0] phv_header_4; // @[executor.scala 448:22]
  reg [15:0] phv_header_5; // @[executor.scala 448:22]
  reg [15:0] phv_header_6; // @[executor.scala 448:22]
  reg [15:0] phv_header_7; // @[executor.scala 448:22]
  reg [15:0] phv_header_8; // @[executor.scala 448:22]
  reg [15:0] phv_header_9; // @[executor.scala 448:22]
  reg [15:0] phv_header_10; // @[executor.scala 448:22]
  reg [15:0] phv_header_11; // @[executor.scala 448:22]
  reg [15:0] phv_header_12; // @[executor.scala 448:22]
  reg [15:0] phv_header_13; // @[executor.scala 448:22]
  reg [15:0] phv_header_14; // @[executor.scala 448:22]
  reg [15:0] phv_header_15; // @[executor.scala 448:22]
  reg [7:0] phv_parse_current_state; // @[executor.scala 448:22]
  reg [7:0] phv_parse_current_offset; // @[executor.scala 448:22]
  reg [15:0] phv_parse_transition_field; // @[executor.scala 448:22]
  reg [3:0] phv_next_processor_id; // @[executor.scala 448:22]
  reg  phv_next_config_id; // @[executor.scala 448:22]
  reg  phv_is_valid_processor; // @[executor.scala 448:22]
  reg  phv_valid; // @[executor.scala 448:22]
  reg [31:0] vliw_0; // @[executor.scala 452:23]
  reg [31:0] vliw_1; // @[executor.scala 452:23]
  reg [31:0] vliw_2; // @[executor.scala 452:23]
  reg [31:0] vliw_3; // @[executor.scala 452:23]
  reg [31:0] field_0; // @[executor.scala 454:24]
  reg [31:0] field_1; // @[executor.scala 454:24]
  reg [31:0] field_2; // @[executor.scala 454:24]
  reg [31:0] field_3; // @[executor.scala 454:24]
  reg [3:0] mask_0; // @[executor.scala 456:23]
  reg [3:0] mask_1; // @[executor.scala 456:23]
  reg [3:0] mask_2; // @[executor.scala 456:23]
  reg [3:0] mask_3; // @[executor.scala 456:23]
  reg [5:0] dst_offset_0; // @[executor.scala 458:29]
  reg [5:0] dst_offset_1; // @[executor.scala 458:29]
  reg [5:0] dst_offset_2; // @[executor.scala 458:29]
  reg [5:0] dst_offset_3; // @[executor.scala 458:29]
  wire [3:0] opcode = vliw_0[31:28]; // @[primitive.scala 9:44]
  wire [13:0] parameter_2 = vliw_0[13:0]; // @[primitive.scala 11:44]
  wire [7:0] _GEN_2730 = {{2'd0}, dst_offset_0}; // @[executor.scala 473:49]
  wire [7:0] byte_ = field_0[7:0]; // @[executor.scala 475:56]
  wire [7:0] _GEN_0 = mask_0[0] ? byte_ : phv_data_3; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] byte_1 = field_0[15:8]; // @[executor.scala 475:56]
  wire [7:0] _GEN_1 = mask_0[1] ? byte_1 : phv_data_2; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] byte_2 = field_0[23:16]; // @[executor.scala 475:56]
  wire [7:0] _GEN_2 = mask_0[2] ? byte_2 : phv_data_1; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] byte_3 = field_0[31:24]; // @[executor.scala 475:56]
  wire [7:0] _GEN_3 = mask_0[3] ? byte_3 : phv_data_0; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_4 = _GEN_2730 == 8'h0 ? _GEN_0 : phv_data_3; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_5 = _GEN_2730 == 8'h0 ? _GEN_1 : phv_data_2; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_6 = _GEN_2730 == 8'h0 ? _GEN_2 : phv_data_1; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_7 = _GEN_2730 == 8'h0 ? _GEN_3 : phv_data_0; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_8 = mask_0[0] ? byte_ : phv_data_7; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_9 = mask_0[1] ? byte_1 : phv_data_6; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_10 = mask_0[2] ? byte_2 : phv_data_5; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_11 = mask_0[3] ? byte_3 : phv_data_4; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_12 = _GEN_2730 == 8'h1 ? _GEN_8 : phv_data_7; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_13 = _GEN_2730 == 8'h1 ? _GEN_9 : phv_data_6; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_14 = _GEN_2730 == 8'h1 ? _GEN_10 : phv_data_5; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_15 = _GEN_2730 == 8'h1 ? _GEN_11 : phv_data_4; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_16 = mask_0[0] ? byte_ : phv_data_11; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_17 = mask_0[1] ? byte_1 : phv_data_10; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_18 = mask_0[2] ? byte_2 : phv_data_9; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_19 = mask_0[3] ? byte_3 : phv_data_8; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_20 = _GEN_2730 == 8'h2 ? _GEN_16 : phv_data_11; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_21 = _GEN_2730 == 8'h2 ? _GEN_17 : phv_data_10; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_22 = _GEN_2730 == 8'h2 ? _GEN_18 : phv_data_9; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_23 = _GEN_2730 == 8'h2 ? _GEN_19 : phv_data_8; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_24 = mask_0[0] ? byte_ : phv_data_15; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_25 = mask_0[1] ? byte_1 : phv_data_14; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_26 = mask_0[2] ? byte_2 : phv_data_13; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_27 = mask_0[3] ? byte_3 : phv_data_12; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_28 = _GEN_2730 == 8'h3 ? _GEN_24 : phv_data_15; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_29 = _GEN_2730 == 8'h3 ? _GEN_25 : phv_data_14; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_30 = _GEN_2730 == 8'h3 ? _GEN_26 : phv_data_13; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_31 = _GEN_2730 == 8'h3 ? _GEN_27 : phv_data_12; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_32 = mask_0[0] ? byte_ : phv_data_19; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_33 = mask_0[1] ? byte_1 : phv_data_18; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_34 = mask_0[2] ? byte_2 : phv_data_17; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_35 = mask_0[3] ? byte_3 : phv_data_16; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_36 = _GEN_2730 == 8'h4 ? _GEN_32 : phv_data_19; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_37 = _GEN_2730 == 8'h4 ? _GEN_33 : phv_data_18; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_38 = _GEN_2730 == 8'h4 ? _GEN_34 : phv_data_17; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_39 = _GEN_2730 == 8'h4 ? _GEN_35 : phv_data_16; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_40 = mask_0[0] ? byte_ : phv_data_23; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_41 = mask_0[1] ? byte_1 : phv_data_22; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_42 = mask_0[2] ? byte_2 : phv_data_21; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_43 = mask_0[3] ? byte_3 : phv_data_20; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_44 = _GEN_2730 == 8'h5 ? _GEN_40 : phv_data_23; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_45 = _GEN_2730 == 8'h5 ? _GEN_41 : phv_data_22; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_46 = _GEN_2730 == 8'h5 ? _GEN_42 : phv_data_21; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_47 = _GEN_2730 == 8'h5 ? _GEN_43 : phv_data_20; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_48 = mask_0[0] ? byte_ : phv_data_27; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_49 = mask_0[1] ? byte_1 : phv_data_26; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_50 = mask_0[2] ? byte_2 : phv_data_25; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_51 = mask_0[3] ? byte_3 : phv_data_24; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_52 = _GEN_2730 == 8'h6 ? _GEN_48 : phv_data_27; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_53 = _GEN_2730 == 8'h6 ? _GEN_49 : phv_data_26; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_54 = _GEN_2730 == 8'h6 ? _GEN_50 : phv_data_25; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_55 = _GEN_2730 == 8'h6 ? _GEN_51 : phv_data_24; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_56 = mask_0[0] ? byte_ : phv_data_31; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_57 = mask_0[1] ? byte_1 : phv_data_30; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_58 = mask_0[2] ? byte_2 : phv_data_29; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_59 = mask_0[3] ? byte_3 : phv_data_28; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_60 = _GEN_2730 == 8'h7 ? _GEN_56 : phv_data_31; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_61 = _GEN_2730 == 8'h7 ? _GEN_57 : phv_data_30; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_62 = _GEN_2730 == 8'h7 ? _GEN_58 : phv_data_29; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_63 = _GEN_2730 == 8'h7 ? _GEN_59 : phv_data_28; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_64 = mask_0[0] ? byte_ : phv_data_35; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_65 = mask_0[1] ? byte_1 : phv_data_34; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_66 = mask_0[2] ? byte_2 : phv_data_33; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_67 = mask_0[3] ? byte_3 : phv_data_32; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_68 = _GEN_2730 == 8'h8 ? _GEN_64 : phv_data_35; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_69 = _GEN_2730 == 8'h8 ? _GEN_65 : phv_data_34; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_70 = _GEN_2730 == 8'h8 ? _GEN_66 : phv_data_33; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_71 = _GEN_2730 == 8'h8 ? _GEN_67 : phv_data_32; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_72 = mask_0[0] ? byte_ : phv_data_39; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_73 = mask_0[1] ? byte_1 : phv_data_38; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_74 = mask_0[2] ? byte_2 : phv_data_37; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_75 = mask_0[3] ? byte_3 : phv_data_36; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_76 = _GEN_2730 == 8'h9 ? _GEN_72 : phv_data_39; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_77 = _GEN_2730 == 8'h9 ? _GEN_73 : phv_data_38; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_78 = _GEN_2730 == 8'h9 ? _GEN_74 : phv_data_37; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_79 = _GEN_2730 == 8'h9 ? _GEN_75 : phv_data_36; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_80 = mask_0[0] ? byte_ : phv_data_43; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_81 = mask_0[1] ? byte_1 : phv_data_42; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_82 = mask_0[2] ? byte_2 : phv_data_41; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_83 = mask_0[3] ? byte_3 : phv_data_40; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_84 = _GEN_2730 == 8'ha ? _GEN_80 : phv_data_43; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_85 = _GEN_2730 == 8'ha ? _GEN_81 : phv_data_42; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_86 = _GEN_2730 == 8'ha ? _GEN_82 : phv_data_41; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_87 = _GEN_2730 == 8'ha ? _GEN_83 : phv_data_40; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_88 = mask_0[0] ? byte_ : phv_data_47; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_89 = mask_0[1] ? byte_1 : phv_data_46; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_90 = mask_0[2] ? byte_2 : phv_data_45; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_91 = mask_0[3] ? byte_3 : phv_data_44; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_92 = _GEN_2730 == 8'hb ? _GEN_88 : phv_data_47; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_93 = _GEN_2730 == 8'hb ? _GEN_89 : phv_data_46; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_94 = _GEN_2730 == 8'hb ? _GEN_90 : phv_data_45; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_95 = _GEN_2730 == 8'hb ? _GEN_91 : phv_data_44; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_96 = mask_0[0] ? byte_ : phv_data_51; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_97 = mask_0[1] ? byte_1 : phv_data_50; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_98 = mask_0[2] ? byte_2 : phv_data_49; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_99 = mask_0[3] ? byte_3 : phv_data_48; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_100 = _GEN_2730 == 8'hc ? _GEN_96 : phv_data_51; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_101 = _GEN_2730 == 8'hc ? _GEN_97 : phv_data_50; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_102 = _GEN_2730 == 8'hc ? _GEN_98 : phv_data_49; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_103 = _GEN_2730 == 8'hc ? _GEN_99 : phv_data_48; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_104 = mask_0[0] ? byte_ : phv_data_55; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_105 = mask_0[1] ? byte_1 : phv_data_54; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_106 = mask_0[2] ? byte_2 : phv_data_53; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_107 = mask_0[3] ? byte_3 : phv_data_52; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_108 = _GEN_2730 == 8'hd ? _GEN_104 : phv_data_55; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_109 = _GEN_2730 == 8'hd ? _GEN_105 : phv_data_54; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_110 = _GEN_2730 == 8'hd ? _GEN_106 : phv_data_53; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_111 = _GEN_2730 == 8'hd ? _GEN_107 : phv_data_52; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_112 = mask_0[0] ? byte_ : phv_data_59; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_113 = mask_0[1] ? byte_1 : phv_data_58; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_114 = mask_0[2] ? byte_2 : phv_data_57; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_115 = mask_0[3] ? byte_3 : phv_data_56; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_116 = _GEN_2730 == 8'he ? _GEN_112 : phv_data_59; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_117 = _GEN_2730 == 8'he ? _GEN_113 : phv_data_58; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_118 = _GEN_2730 == 8'he ? _GEN_114 : phv_data_57; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_119 = _GEN_2730 == 8'he ? _GEN_115 : phv_data_56; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_120 = mask_0[0] ? byte_ : phv_data_63; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_121 = mask_0[1] ? byte_1 : phv_data_62; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_122 = mask_0[2] ? byte_2 : phv_data_61; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_123 = mask_0[3] ? byte_3 : phv_data_60; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_124 = _GEN_2730 == 8'hf ? _GEN_120 : phv_data_63; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_125 = _GEN_2730 == 8'hf ? _GEN_121 : phv_data_62; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_126 = _GEN_2730 == 8'hf ? _GEN_122 : phv_data_61; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_127 = _GEN_2730 == 8'hf ? _GEN_123 : phv_data_60; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_128 = mask_0[0] ? byte_ : phv_data_67; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_129 = mask_0[1] ? byte_1 : phv_data_66; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_130 = mask_0[2] ? byte_2 : phv_data_65; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_131 = mask_0[3] ? byte_3 : phv_data_64; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_132 = _GEN_2730 == 8'h10 ? _GEN_128 : phv_data_67; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_133 = _GEN_2730 == 8'h10 ? _GEN_129 : phv_data_66; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_134 = _GEN_2730 == 8'h10 ? _GEN_130 : phv_data_65; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_135 = _GEN_2730 == 8'h10 ? _GEN_131 : phv_data_64; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_136 = mask_0[0] ? byte_ : phv_data_71; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_137 = mask_0[1] ? byte_1 : phv_data_70; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_138 = mask_0[2] ? byte_2 : phv_data_69; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_139 = mask_0[3] ? byte_3 : phv_data_68; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_140 = _GEN_2730 == 8'h11 ? _GEN_136 : phv_data_71; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_141 = _GEN_2730 == 8'h11 ? _GEN_137 : phv_data_70; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_142 = _GEN_2730 == 8'h11 ? _GEN_138 : phv_data_69; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_143 = _GEN_2730 == 8'h11 ? _GEN_139 : phv_data_68; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_144 = mask_0[0] ? byte_ : phv_data_75; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_145 = mask_0[1] ? byte_1 : phv_data_74; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_146 = mask_0[2] ? byte_2 : phv_data_73; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_147 = mask_0[3] ? byte_3 : phv_data_72; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_148 = _GEN_2730 == 8'h12 ? _GEN_144 : phv_data_75; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_149 = _GEN_2730 == 8'h12 ? _GEN_145 : phv_data_74; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_150 = _GEN_2730 == 8'h12 ? _GEN_146 : phv_data_73; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_151 = _GEN_2730 == 8'h12 ? _GEN_147 : phv_data_72; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_152 = mask_0[0] ? byte_ : phv_data_79; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_153 = mask_0[1] ? byte_1 : phv_data_78; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_154 = mask_0[2] ? byte_2 : phv_data_77; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_155 = mask_0[3] ? byte_3 : phv_data_76; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_156 = _GEN_2730 == 8'h13 ? _GEN_152 : phv_data_79; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_157 = _GEN_2730 == 8'h13 ? _GEN_153 : phv_data_78; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_158 = _GEN_2730 == 8'h13 ? _GEN_154 : phv_data_77; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_159 = _GEN_2730 == 8'h13 ? _GEN_155 : phv_data_76; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_160 = mask_0[0] ? byte_ : phv_data_83; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_161 = mask_0[1] ? byte_1 : phv_data_82; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_162 = mask_0[2] ? byte_2 : phv_data_81; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_163 = mask_0[3] ? byte_3 : phv_data_80; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_164 = _GEN_2730 == 8'h14 ? _GEN_160 : phv_data_83; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_165 = _GEN_2730 == 8'h14 ? _GEN_161 : phv_data_82; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_166 = _GEN_2730 == 8'h14 ? _GEN_162 : phv_data_81; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_167 = _GEN_2730 == 8'h14 ? _GEN_163 : phv_data_80; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_168 = mask_0[0] ? byte_ : phv_data_87; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_169 = mask_0[1] ? byte_1 : phv_data_86; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_170 = mask_0[2] ? byte_2 : phv_data_85; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_171 = mask_0[3] ? byte_3 : phv_data_84; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_172 = _GEN_2730 == 8'h15 ? _GEN_168 : phv_data_87; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_173 = _GEN_2730 == 8'h15 ? _GEN_169 : phv_data_86; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_174 = _GEN_2730 == 8'h15 ? _GEN_170 : phv_data_85; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_175 = _GEN_2730 == 8'h15 ? _GEN_171 : phv_data_84; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_176 = mask_0[0] ? byte_ : phv_data_91; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_177 = mask_0[1] ? byte_1 : phv_data_90; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_178 = mask_0[2] ? byte_2 : phv_data_89; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_179 = mask_0[3] ? byte_3 : phv_data_88; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_180 = _GEN_2730 == 8'h16 ? _GEN_176 : phv_data_91; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_181 = _GEN_2730 == 8'h16 ? _GEN_177 : phv_data_90; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_182 = _GEN_2730 == 8'h16 ? _GEN_178 : phv_data_89; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_183 = _GEN_2730 == 8'h16 ? _GEN_179 : phv_data_88; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_184 = mask_0[0] ? byte_ : phv_data_95; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_185 = mask_0[1] ? byte_1 : phv_data_94; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_186 = mask_0[2] ? byte_2 : phv_data_93; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_187 = mask_0[3] ? byte_3 : phv_data_92; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_188 = _GEN_2730 == 8'h17 ? _GEN_184 : phv_data_95; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_189 = _GEN_2730 == 8'h17 ? _GEN_185 : phv_data_94; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_190 = _GEN_2730 == 8'h17 ? _GEN_186 : phv_data_93; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_191 = _GEN_2730 == 8'h17 ? _GEN_187 : phv_data_92; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_192 = mask_0[0] ? byte_ : phv_data_99; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_193 = mask_0[1] ? byte_1 : phv_data_98; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_194 = mask_0[2] ? byte_2 : phv_data_97; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_195 = mask_0[3] ? byte_3 : phv_data_96; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_196 = _GEN_2730 == 8'h18 ? _GEN_192 : phv_data_99; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_197 = _GEN_2730 == 8'h18 ? _GEN_193 : phv_data_98; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_198 = _GEN_2730 == 8'h18 ? _GEN_194 : phv_data_97; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_199 = _GEN_2730 == 8'h18 ? _GEN_195 : phv_data_96; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_200 = mask_0[0] ? byte_ : phv_data_103; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_201 = mask_0[1] ? byte_1 : phv_data_102; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_202 = mask_0[2] ? byte_2 : phv_data_101; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_203 = mask_0[3] ? byte_3 : phv_data_100; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_204 = _GEN_2730 == 8'h19 ? _GEN_200 : phv_data_103; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_205 = _GEN_2730 == 8'h19 ? _GEN_201 : phv_data_102; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_206 = _GEN_2730 == 8'h19 ? _GEN_202 : phv_data_101; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_207 = _GEN_2730 == 8'h19 ? _GEN_203 : phv_data_100; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_208 = mask_0[0] ? byte_ : phv_data_107; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_209 = mask_0[1] ? byte_1 : phv_data_106; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_210 = mask_0[2] ? byte_2 : phv_data_105; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_211 = mask_0[3] ? byte_3 : phv_data_104; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_212 = _GEN_2730 == 8'h1a ? _GEN_208 : phv_data_107; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_213 = _GEN_2730 == 8'h1a ? _GEN_209 : phv_data_106; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_214 = _GEN_2730 == 8'h1a ? _GEN_210 : phv_data_105; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_215 = _GEN_2730 == 8'h1a ? _GEN_211 : phv_data_104; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_216 = mask_0[0] ? byte_ : phv_data_111; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_217 = mask_0[1] ? byte_1 : phv_data_110; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_218 = mask_0[2] ? byte_2 : phv_data_109; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_219 = mask_0[3] ? byte_3 : phv_data_108; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_220 = _GEN_2730 == 8'h1b ? _GEN_216 : phv_data_111; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_221 = _GEN_2730 == 8'h1b ? _GEN_217 : phv_data_110; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_222 = _GEN_2730 == 8'h1b ? _GEN_218 : phv_data_109; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_223 = _GEN_2730 == 8'h1b ? _GEN_219 : phv_data_108; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_224 = mask_0[0] ? byte_ : phv_data_115; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_225 = mask_0[1] ? byte_1 : phv_data_114; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_226 = mask_0[2] ? byte_2 : phv_data_113; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_227 = mask_0[3] ? byte_3 : phv_data_112; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_228 = _GEN_2730 == 8'h1c ? _GEN_224 : phv_data_115; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_229 = _GEN_2730 == 8'h1c ? _GEN_225 : phv_data_114; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_230 = _GEN_2730 == 8'h1c ? _GEN_226 : phv_data_113; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_231 = _GEN_2730 == 8'h1c ? _GEN_227 : phv_data_112; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_232 = mask_0[0] ? byte_ : phv_data_119; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_233 = mask_0[1] ? byte_1 : phv_data_118; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_234 = mask_0[2] ? byte_2 : phv_data_117; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_235 = mask_0[3] ? byte_3 : phv_data_116; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_236 = _GEN_2730 == 8'h1d ? _GEN_232 : phv_data_119; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_237 = _GEN_2730 == 8'h1d ? _GEN_233 : phv_data_118; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_238 = _GEN_2730 == 8'h1d ? _GEN_234 : phv_data_117; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_239 = _GEN_2730 == 8'h1d ? _GEN_235 : phv_data_116; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_240 = mask_0[0] ? byte_ : phv_data_123; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_241 = mask_0[1] ? byte_1 : phv_data_122; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_242 = mask_0[2] ? byte_2 : phv_data_121; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_243 = mask_0[3] ? byte_3 : phv_data_120; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_244 = _GEN_2730 == 8'h1e ? _GEN_240 : phv_data_123; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_245 = _GEN_2730 == 8'h1e ? _GEN_241 : phv_data_122; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_246 = _GEN_2730 == 8'h1e ? _GEN_242 : phv_data_121; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_247 = _GEN_2730 == 8'h1e ? _GEN_243 : phv_data_120; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_248 = mask_0[0] ? byte_ : phv_data_127; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_249 = mask_0[1] ? byte_1 : phv_data_126; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_250 = mask_0[2] ? byte_2 : phv_data_125; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_251 = mask_0[3] ? byte_3 : phv_data_124; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_252 = _GEN_2730 == 8'h1f ? _GEN_248 : phv_data_127; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_253 = _GEN_2730 == 8'h1f ? _GEN_249 : phv_data_126; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_254 = _GEN_2730 == 8'h1f ? _GEN_250 : phv_data_125; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_255 = _GEN_2730 == 8'h1f ? _GEN_251 : phv_data_124; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_256 = mask_0[0] ? byte_ : phv_data_131; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_257 = mask_0[1] ? byte_1 : phv_data_130; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_258 = mask_0[2] ? byte_2 : phv_data_129; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_259 = mask_0[3] ? byte_3 : phv_data_128; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_260 = _GEN_2730 == 8'h20 ? _GEN_256 : phv_data_131; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_261 = _GEN_2730 == 8'h20 ? _GEN_257 : phv_data_130; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_262 = _GEN_2730 == 8'h20 ? _GEN_258 : phv_data_129; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_263 = _GEN_2730 == 8'h20 ? _GEN_259 : phv_data_128; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_264 = mask_0[0] ? byte_ : phv_data_135; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_265 = mask_0[1] ? byte_1 : phv_data_134; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_266 = mask_0[2] ? byte_2 : phv_data_133; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_267 = mask_0[3] ? byte_3 : phv_data_132; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_268 = _GEN_2730 == 8'h21 ? _GEN_264 : phv_data_135; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_269 = _GEN_2730 == 8'h21 ? _GEN_265 : phv_data_134; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_270 = _GEN_2730 == 8'h21 ? _GEN_266 : phv_data_133; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_271 = _GEN_2730 == 8'h21 ? _GEN_267 : phv_data_132; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_272 = mask_0[0] ? byte_ : phv_data_139; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_273 = mask_0[1] ? byte_1 : phv_data_138; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_274 = mask_0[2] ? byte_2 : phv_data_137; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_275 = mask_0[3] ? byte_3 : phv_data_136; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_276 = _GEN_2730 == 8'h22 ? _GEN_272 : phv_data_139; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_277 = _GEN_2730 == 8'h22 ? _GEN_273 : phv_data_138; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_278 = _GEN_2730 == 8'h22 ? _GEN_274 : phv_data_137; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_279 = _GEN_2730 == 8'h22 ? _GEN_275 : phv_data_136; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_280 = mask_0[0] ? byte_ : phv_data_143; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_281 = mask_0[1] ? byte_1 : phv_data_142; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_282 = mask_0[2] ? byte_2 : phv_data_141; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_283 = mask_0[3] ? byte_3 : phv_data_140; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_284 = _GEN_2730 == 8'h23 ? _GEN_280 : phv_data_143; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_285 = _GEN_2730 == 8'h23 ? _GEN_281 : phv_data_142; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_286 = _GEN_2730 == 8'h23 ? _GEN_282 : phv_data_141; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_287 = _GEN_2730 == 8'h23 ? _GEN_283 : phv_data_140; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_288 = mask_0[0] ? byte_ : phv_data_147; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_289 = mask_0[1] ? byte_1 : phv_data_146; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_290 = mask_0[2] ? byte_2 : phv_data_145; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_291 = mask_0[3] ? byte_3 : phv_data_144; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_292 = _GEN_2730 == 8'h24 ? _GEN_288 : phv_data_147; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_293 = _GEN_2730 == 8'h24 ? _GEN_289 : phv_data_146; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_294 = _GEN_2730 == 8'h24 ? _GEN_290 : phv_data_145; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_295 = _GEN_2730 == 8'h24 ? _GEN_291 : phv_data_144; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_296 = mask_0[0] ? byte_ : phv_data_151; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_297 = mask_0[1] ? byte_1 : phv_data_150; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_298 = mask_0[2] ? byte_2 : phv_data_149; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_299 = mask_0[3] ? byte_3 : phv_data_148; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_300 = _GEN_2730 == 8'h25 ? _GEN_296 : phv_data_151; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_301 = _GEN_2730 == 8'h25 ? _GEN_297 : phv_data_150; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_302 = _GEN_2730 == 8'h25 ? _GEN_298 : phv_data_149; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_303 = _GEN_2730 == 8'h25 ? _GEN_299 : phv_data_148; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_304 = mask_0[0] ? byte_ : phv_data_155; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_305 = mask_0[1] ? byte_1 : phv_data_154; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_306 = mask_0[2] ? byte_2 : phv_data_153; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_307 = mask_0[3] ? byte_3 : phv_data_152; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_308 = _GEN_2730 == 8'h26 ? _GEN_304 : phv_data_155; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_309 = _GEN_2730 == 8'h26 ? _GEN_305 : phv_data_154; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_310 = _GEN_2730 == 8'h26 ? _GEN_306 : phv_data_153; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_311 = _GEN_2730 == 8'h26 ? _GEN_307 : phv_data_152; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_312 = mask_0[0] ? byte_ : phv_data_159; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_313 = mask_0[1] ? byte_1 : phv_data_158; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_314 = mask_0[2] ? byte_2 : phv_data_157; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_315 = mask_0[3] ? byte_3 : phv_data_156; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_316 = _GEN_2730 == 8'h27 ? _GEN_312 : phv_data_159; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_317 = _GEN_2730 == 8'h27 ? _GEN_313 : phv_data_158; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_318 = _GEN_2730 == 8'h27 ? _GEN_314 : phv_data_157; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_319 = _GEN_2730 == 8'h27 ? _GEN_315 : phv_data_156; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_320 = opcode != 4'h0 ? _GEN_4 : phv_data_3; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_321 = opcode != 4'h0 ? _GEN_5 : phv_data_2; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_322 = opcode != 4'h0 ? _GEN_6 : phv_data_1; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_323 = opcode != 4'h0 ? _GEN_7 : phv_data_0; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_324 = opcode != 4'h0 ? _GEN_12 : phv_data_7; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_325 = opcode != 4'h0 ? _GEN_13 : phv_data_6; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_326 = opcode != 4'h0 ? _GEN_14 : phv_data_5; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_327 = opcode != 4'h0 ? _GEN_15 : phv_data_4; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_328 = opcode != 4'h0 ? _GEN_20 : phv_data_11; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_329 = opcode != 4'h0 ? _GEN_21 : phv_data_10; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_330 = opcode != 4'h0 ? _GEN_22 : phv_data_9; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_331 = opcode != 4'h0 ? _GEN_23 : phv_data_8; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_332 = opcode != 4'h0 ? _GEN_28 : phv_data_15; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_333 = opcode != 4'h0 ? _GEN_29 : phv_data_14; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_334 = opcode != 4'h0 ? _GEN_30 : phv_data_13; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_335 = opcode != 4'h0 ? _GEN_31 : phv_data_12; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_336 = opcode != 4'h0 ? _GEN_36 : phv_data_19; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_337 = opcode != 4'h0 ? _GEN_37 : phv_data_18; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_338 = opcode != 4'h0 ? _GEN_38 : phv_data_17; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_339 = opcode != 4'h0 ? _GEN_39 : phv_data_16; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_340 = opcode != 4'h0 ? _GEN_44 : phv_data_23; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_341 = opcode != 4'h0 ? _GEN_45 : phv_data_22; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_342 = opcode != 4'h0 ? _GEN_46 : phv_data_21; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_343 = opcode != 4'h0 ? _GEN_47 : phv_data_20; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_344 = opcode != 4'h0 ? _GEN_52 : phv_data_27; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_345 = opcode != 4'h0 ? _GEN_53 : phv_data_26; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_346 = opcode != 4'h0 ? _GEN_54 : phv_data_25; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_347 = opcode != 4'h0 ? _GEN_55 : phv_data_24; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_348 = opcode != 4'h0 ? _GEN_60 : phv_data_31; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_349 = opcode != 4'h0 ? _GEN_61 : phv_data_30; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_350 = opcode != 4'h0 ? _GEN_62 : phv_data_29; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_351 = opcode != 4'h0 ? _GEN_63 : phv_data_28; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_352 = opcode != 4'h0 ? _GEN_68 : phv_data_35; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_353 = opcode != 4'h0 ? _GEN_69 : phv_data_34; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_354 = opcode != 4'h0 ? _GEN_70 : phv_data_33; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_355 = opcode != 4'h0 ? _GEN_71 : phv_data_32; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_356 = opcode != 4'h0 ? _GEN_76 : phv_data_39; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_357 = opcode != 4'h0 ? _GEN_77 : phv_data_38; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_358 = opcode != 4'h0 ? _GEN_78 : phv_data_37; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_359 = opcode != 4'h0 ? _GEN_79 : phv_data_36; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_360 = opcode != 4'h0 ? _GEN_84 : phv_data_43; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_361 = opcode != 4'h0 ? _GEN_85 : phv_data_42; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_362 = opcode != 4'h0 ? _GEN_86 : phv_data_41; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_363 = opcode != 4'h0 ? _GEN_87 : phv_data_40; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_364 = opcode != 4'h0 ? _GEN_92 : phv_data_47; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_365 = opcode != 4'h0 ? _GEN_93 : phv_data_46; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_366 = opcode != 4'h0 ? _GEN_94 : phv_data_45; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_367 = opcode != 4'h0 ? _GEN_95 : phv_data_44; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_368 = opcode != 4'h0 ? _GEN_100 : phv_data_51; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_369 = opcode != 4'h0 ? _GEN_101 : phv_data_50; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_370 = opcode != 4'h0 ? _GEN_102 : phv_data_49; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_371 = opcode != 4'h0 ? _GEN_103 : phv_data_48; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_372 = opcode != 4'h0 ? _GEN_108 : phv_data_55; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_373 = opcode != 4'h0 ? _GEN_109 : phv_data_54; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_374 = opcode != 4'h0 ? _GEN_110 : phv_data_53; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_375 = opcode != 4'h0 ? _GEN_111 : phv_data_52; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_376 = opcode != 4'h0 ? _GEN_116 : phv_data_59; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_377 = opcode != 4'h0 ? _GEN_117 : phv_data_58; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_378 = opcode != 4'h0 ? _GEN_118 : phv_data_57; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_379 = opcode != 4'h0 ? _GEN_119 : phv_data_56; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_380 = opcode != 4'h0 ? _GEN_124 : phv_data_63; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_381 = opcode != 4'h0 ? _GEN_125 : phv_data_62; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_382 = opcode != 4'h0 ? _GEN_126 : phv_data_61; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_383 = opcode != 4'h0 ? _GEN_127 : phv_data_60; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_384 = opcode != 4'h0 ? _GEN_132 : phv_data_67; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_385 = opcode != 4'h0 ? _GEN_133 : phv_data_66; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_386 = opcode != 4'h0 ? _GEN_134 : phv_data_65; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_387 = opcode != 4'h0 ? _GEN_135 : phv_data_64; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_388 = opcode != 4'h0 ? _GEN_140 : phv_data_71; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_389 = opcode != 4'h0 ? _GEN_141 : phv_data_70; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_390 = opcode != 4'h0 ? _GEN_142 : phv_data_69; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_391 = opcode != 4'h0 ? _GEN_143 : phv_data_68; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_392 = opcode != 4'h0 ? _GEN_148 : phv_data_75; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_393 = opcode != 4'h0 ? _GEN_149 : phv_data_74; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_394 = opcode != 4'h0 ? _GEN_150 : phv_data_73; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_395 = opcode != 4'h0 ? _GEN_151 : phv_data_72; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_396 = opcode != 4'h0 ? _GEN_156 : phv_data_79; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_397 = opcode != 4'h0 ? _GEN_157 : phv_data_78; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_398 = opcode != 4'h0 ? _GEN_158 : phv_data_77; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_399 = opcode != 4'h0 ? _GEN_159 : phv_data_76; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_400 = opcode != 4'h0 ? _GEN_164 : phv_data_83; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_401 = opcode != 4'h0 ? _GEN_165 : phv_data_82; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_402 = opcode != 4'h0 ? _GEN_166 : phv_data_81; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_403 = opcode != 4'h0 ? _GEN_167 : phv_data_80; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_404 = opcode != 4'h0 ? _GEN_172 : phv_data_87; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_405 = opcode != 4'h0 ? _GEN_173 : phv_data_86; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_406 = opcode != 4'h0 ? _GEN_174 : phv_data_85; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_407 = opcode != 4'h0 ? _GEN_175 : phv_data_84; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_408 = opcode != 4'h0 ? _GEN_180 : phv_data_91; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_409 = opcode != 4'h0 ? _GEN_181 : phv_data_90; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_410 = opcode != 4'h0 ? _GEN_182 : phv_data_89; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_411 = opcode != 4'h0 ? _GEN_183 : phv_data_88; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_412 = opcode != 4'h0 ? _GEN_188 : phv_data_95; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_413 = opcode != 4'h0 ? _GEN_189 : phv_data_94; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_414 = opcode != 4'h0 ? _GEN_190 : phv_data_93; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_415 = opcode != 4'h0 ? _GEN_191 : phv_data_92; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_416 = opcode != 4'h0 ? _GEN_196 : phv_data_99; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_417 = opcode != 4'h0 ? _GEN_197 : phv_data_98; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_418 = opcode != 4'h0 ? _GEN_198 : phv_data_97; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_419 = opcode != 4'h0 ? _GEN_199 : phv_data_96; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_420 = opcode != 4'h0 ? _GEN_204 : phv_data_103; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_421 = opcode != 4'h0 ? _GEN_205 : phv_data_102; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_422 = opcode != 4'h0 ? _GEN_206 : phv_data_101; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_423 = opcode != 4'h0 ? _GEN_207 : phv_data_100; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_424 = opcode != 4'h0 ? _GEN_212 : phv_data_107; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_425 = opcode != 4'h0 ? _GEN_213 : phv_data_106; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_426 = opcode != 4'h0 ? _GEN_214 : phv_data_105; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_427 = opcode != 4'h0 ? _GEN_215 : phv_data_104; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_428 = opcode != 4'h0 ? _GEN_220 : phv_data_111; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_429 = opcode != 4'h0 ? _GEN_221 : phv_data_110; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_430 = opcode != 4'h0 ? _GEN_222 : phv_data_109; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_431 = opcode != 4'h0 ? _GEN_223 : phv_data_108; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_432 = opcode != 4'h0 ? _GEN_228 : phv_data_115; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_433 = opcode != 4'h0 ? _GEN_229 : phv_data_114; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_434 = opcode != 4'h0 ? _GEN_230 : phv_data_113; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_435 = opcode != 4'h0 ? _GEN_231 : phv_data_112; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_436 = opcode != 4'h0 ? _GEN_236 : phv_data_119; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_437 = opcode != 4'h0 ? _GEN_237 : phv_data_118; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_438 = opcode != 4'h0 ? _GEN_238 : phv_data_117; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_439 = opcode != 4'h0 ? _GEN_239 : phv_data_116; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_440 = opcode != 4'h0 ? _GEN_244 : phv_data_123; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_441 = opcode != 4'h0 ? _GEN_245 : phv_data_122; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_442 = opcode != 4'h0 ? _GEN_246 : phv_data_121; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_443 = opcode != 4'h0 ? _GEN_247 : phv_data_120; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_444 = opcode != 4'h0 ? _GEN_252 : phv_data_127; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_445 = opcode != 4'h0 ? _GEN_253 : phv_data_126; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_446 = opcode != 4'h0 ? _GEN_254 : phv_data_125; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_447 = opcode != 4'h0 ? _GEN_255 : phv_data_124; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_448 = opcode != 4'h0 ? _GEN_260 : phv_data_131; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_449 = opcode != 4'h0 ? _GEN_261 : phv_data_130; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_450 = opcode != 4'h0 ? _GEN_262 : phv_data_129; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_451 = opcode != 4'h0 ? _GEN_263 : phv_data_128; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_452 = opcode != 4'h0 ? _GEN_268 : phv_data_135; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_453 = opcode != 4'h0 ? _GEN_269 : phv_data_134; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_454 = opcode != 4'h0 ? _GEN_270 : phv_data_133; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_455 = opcode != 4'h0 ? _GEN_271 : phv_data_132; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_456 = opcode != 4'h0 ? _GEN_276 : phv_data_139; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_457 = opcode != 4'h0 ? _GEN_277 : phv_data_138; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_458 = opcode != 4'h0 ? _GEN_278 : phv_data_137; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_459 = opcode != 4'h0 ? _GEN_279 : phv_data_136; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_460 = opcode != 4'h0 ? _GEN_284 : phv_data_143; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_461 = opcode != 4'h0 ? _GEN_285 : phv_data_142; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_462 = opcode != 4'h0 ? _GEN_286 : phv_data_141; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_463 = opcode != 4'h0 ? _GEN_287 : phv_data_140; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_464 = opcode != 4'h0 ? _GEN_292 : phv_data_147; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_465 = opcode != 4'h0 ? _GEN_293 : phv_data_146; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_466 = opcode != 4'h0 ? _GEN_294 : phv_data_145; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_467 = opcode != 4'h0 ? _GEN_295 : phv_data_144; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_468 = opcode != 4'h0 ? _GEN_300 : phv_data_151; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_469 = opcode != 4'h0 ? _GEN_301 : phv_data_150; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_470 = opcode != 4'h0 ? _GEN_302 : phv_data_149; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_471 = opcode != 4'h0 ? _GEN_303 : phv_data_148; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_472 = opcode != 4'h0 ? _GEN_308 : phv_data_155; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_473 = opcode != 4'h0 ? _GEN_309 : phv_data_154; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_474 = opcode != 4'h0 ? _GEN_310 : phv_data_153; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_475 = opcode != 4'h0 ? _GEN_311 : phv_data_152; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_476 = opcode != 4'h0 ? _GEN_316 : phv_data_159; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_477 = opcode != 4'h0 ? _GEN_317 : phv_data_158; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_478 = opcode != 4'h0 ? _GEN_318 : phv_data_157; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_479 = opcode != 4'h0 ? _GEN_319 : phv_data_156; // @[executor.scala 470:55 executor.scala 450:25]
  wire [3:0] _GEN_480 = opcode == 4'hf ? parameter_2[13:10] : phv_next_processor_id; // @[executor.scala 466:52 executor.scala 467:55 executor.scala 450:25]
  wire  _GEN_481 = opcode == 4'hf ? parameter_2[0] : phv_next_config_id; // @[executor.scala 466:52 executor.scala 468:55 executor.scala 450:25]
  wire [7:0] _GEN_482 = opcode == 4'hf ? phv_data_3 : _GEN_320; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_483 = opcode == 4'hf ? phv_data_2 : _GEN_321; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_484 = opcode == 4'hf ? phv_data_1 : _GEN_322; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_485 = opcode == 4'hf ? phv_data_0 : _GEN_323; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_486 = opcode == 4'hf ? phv_data_7 : _GEN_324; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_487 = opcode == 4'hf ? phv_data_6 : _GEN_325; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_488 = opcode == 4'hf ? phv_data_5 : _GEN_326; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_489 = opcode == 4'hf ? phv_data_4 : _GEN_327; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_490 = opcode == 4'hf ? phv_data_11 : _GEN_328; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_491 = opcode == 4'hf ? phv_data_10 : _GEN_329; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_492 = opcode == 4'hf ? phv_data_9 : _GEN_330; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_493 = opcode == 4'hf ? phv_data_8 : _GEN_331; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_494 = opcode == 4'hf ? phv_data_15 : _GEN_332; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_495 = opcode == 4'hf ? phv_data_14 : _GEN_333; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_496 = opcode == 4'hf ? phv_data_13 : _GEN_334; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_497 = opcode == 4'hf ? phv_data_12 : _GEN_335; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_498 = opcode == 4'hf ? phv_data_19 : _GEN_336; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_499 = opcode == 4'hf ? phv_data_18 : _GEN_337; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_500 = opcode == 4'hf ? phv_data_17 : _GEN_338; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_501 = opcode == 4'hf ? phv_data_16 : _GEN_339; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_502 = opcode == 4'hf ? phv_data_23 : _GEN_340; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_503 = opcode == 4'hf ? phv_data_22 : _GEN_341; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_504 = opcode == 4'hf ? phv_data_21 : _GEN_342; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_505 = opcode == 4'hf ? phv_data_20 : _GEN_343; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_506 = opcode == 4'hf ? phv_data_27 : _GEN_344; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_507 = opcode == 4'hf ? phv_data_26 : _GEN_345; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_508 = opcode == 4'hf ? phv_data_25 : _GEN_346; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_509 = opcode == 4'hf ? phv_data_24 : _GEN_347; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_510 = opcode == 4'hf ? phv_data_31 : _GEN_348; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_511 = opcode == 4'hf ? phv_data_30 : _GEN_349; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_512 = opcode == 4'hf ? phv_data_29 : _GEN_350; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_513 = opcode == 4'hf ? phv_data_28 : _GEN_351; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_514 = opcode == 4'hf ? phv_data_35 : _GEN_352; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_515 = opcode == 4'hf ? phv_data_34 : _GEN_353; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_516 = opcode == 4'hf ? phv_data_33 : _GEN_354; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_517 = opcode == 4'hf ? phv_data_32 : _GEN_355; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_518 = opcode == 4'hf ? phv_data_39 : _GEN_356; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_519 = opcode == 4'hf ? phv_data_38 : _GEN_357; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_520 = opcode == 4'hf ? phv_data_37 : _GEN_358; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_521 = opcode == 4'hf ? phv_data_36 : _GEN_359; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_522 = opcode == 4'hf ? phv_data_43 : _GEN_360; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_523 = opcode == 4'hf ? phv_data_42 : _GEN_361; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_524 = opcode == 4'hf ? phv_data_41 : _GEN_362; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_525 = opcode == 4'hf ? phv_data_40 : _GEN_363; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_526 = opcode == 4'hf ? phv_data_47 : _GEN_364; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_527 = opcode == 4'hf ? phv_data_46 : _GEN_365; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_528 = opcode == 4'hf ? phv_data_45 : _GEN_366; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_529 = opcode == 4'hf ? phv_data_44 : _GEN_367; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_530 = opcode == 4'hf ? phv_data_51 : _GEN_368; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_531 = opcode == 4'hf ? phv_data_50 : _GEN_369; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_532 = opcode == 4'hf ? phv_data_49 : _GEN_370; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_533 = opcode == 4'hf ? phv_data_48 : _GEN_371; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_534 = opcode == 4'hf ? phv_data_55 : _GEN_372; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_535 = opcode == 4'hf ? phv_data_54 : _GEN_373; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_536 = opcode == 4'hf ? phv_data_53 : _GEN_374; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_537 = opcode == 4'hf ? phv_data_52 : _GEN_375; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_538 = opcode == 4'hf ? phv_data_59 : _GEN_376; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_539 = opcode == 4'hf ? phv_data_58 : _GEN_377; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_540 = opcode == 4'hf ? phv_data_57 : _GEN_378; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_541 = opcode == 4'hf ? phv_data_56 : _GEN_379; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_542 = opcode == 4'hf ? phv_data_63 : _GEN_380; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_543 = opcode == 4'hf ? phv_data_62 : _GEN_381; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_544 = opcode == 4'hf ? phv_data_61 : _GEN_382; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_545 = opcode == 4'hf ? phv_data_60 : _GEN_383; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_546 = opcode == 4'hf ? phv_data_67 : _GEN_384; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_547 = opcode == 4'hf ? phv_data_66 : _GEN_385; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_548 = opcode == 4'hf ? phv_data_65 : _GEN_386; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_549 = opcode == 4'hf ? phv_data_64 : _GEN_387; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_550 = opcode == 4'hf ? phv_data_71 : _GEN_388; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_551 = opcode == 4'hf ? phv_data_70 : _GEN_389; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_552 = opcode == 4'hf ? phv_data_69 : _GEN_390; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_553 = opcode == 4'hf ? phv_data_68 : _GEN_391; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_554 = opcode == 4'hf ? phv_data_75 : _GEN_392; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_555 = opcode == 4'hf ? phv_data_74 : _GEN_393; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_556 = opcode == 4'hf ? phv_data_73 : _GEN_394; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_557 = opcode == 4'hf ? phv_data_72 : _GEN_395; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_558 = opcode == 4'hf ? phv_data_79 : _GEN_396; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_559 = opcode == 4'hf ? phv_data_78 : _GEN_397; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_560 = opcode == 4'hf ? phv_data_77 : _GEN_398; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_561 = opcode == 4'hf ? phv_data_76 : _GEN_399; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_562 = opcode == 4'hf ? phv_data_83 : _GEN_400; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_563 = opcode == 4'hf ? phv_data_82 : _GEN_401; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_564 = opcode == 4'hf ? phv_data_81 : _GEN_402; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_565 = opcode == 4'hf ? phv_data_80 : _GEN_403; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_566 = opcode == 4'hf ? phv_data_87 : _GEN_404; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_567 = opcode == 4'hf ? phv_data_86 : _GEN_405; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_568 = opcode == 4'hf ? phv_data_85 : _GEN_406; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_569 = opcode == 4'hf ? phv_data_84 : _GEN_407; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_570 = opcode == 4'hf ? phv_data_91 : _GEN_408; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_571 = opcode == 4'hf ? phv_data_90 : _GEN_409; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_572 = opcode == 4'hf ? phv_data_89 : _GEN_410; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_573 = opcode == 4'hf ? phv_data_88 : _GEN_411; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_574 = opcode == 4'hf ? phv_data_95 : _GEN_412; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_575 = opcode == 4'hf ? phv_data_94 : _GEN_413; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_576 = opcode == 4'hf ? phv_data_93 : _GEN_414; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_577 = opcode == 4'hf ? phv_data_92 : _GEN_415; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_578 = opcode == 4'hf ? phv_data_99 : _GEN_416; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_579 = opcode == 4'hf ? phv_data_98 : _GEN_417; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_580 = opcode == 4'hf ? phv_data_97 : _GEN_418; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_581 = opcode == 4'hf ? phv_data_96 : _GEN_419; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_582 = opcode == 4'hf ? phv_data_103 : _GEN_420; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_583 = opcode == 4'hf ? phv_data_102 : _GEN_421; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_584 = opcode == 4'hf ? phv_data_101 : _GEN_422; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_585 = opcode == 4'hf ? phv_data_100 : _GEN_423; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_586 = opcode == 4'hf ? phv_data_107 : _GEN_424; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_587 = opcode == 4'hf ? phv_data_106 : _GEN_425; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_588 = opcode == 4'hf ? phv_data_105 : _GEN_426; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_589 = opcode == 4'hf ? phv_data_104 : _GEN_427; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_590 = opcode == 4'hf ? phv_data_111 : _GEN_428; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_591 = opcode == 4'hf ? phv_data_110 : _GEN_429; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_592 = opcode == 4'hf ? phv_data_109 : _GEN_430; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_593 = opcode == 4'hf ? phv_data_108 : _GEN_431; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_594 = opcode == 4'hf ? phv_data_115 : _GEN_432; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_595 = opcode == 4'hf ? phv_data_114 : _GEN_433; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_596 = opcode == 4'hf ? phv_data_113 : _GEN_434; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_597 = opcode == 4'hf ? phv_data_112 : _GEN_435; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_598 = opcode == 4'hf ? phv_data_119 : _GEN_436; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_599 = opcode == 4'hf ? phv_data_118 : _GEN_437; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_600 = opcode == 4'hf ? phv_data_117 : _GEN_438; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_601 = opcode == 4'hf ? phv_data_116 : _GEN_439; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_602 = opcode == 4'hf ? phv_data_123 : _GEN_440; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_603 = opcode == 4'hf ? phv_data_122 : _GEN_441; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_604 = opcode == 4'hf ? phv_data_121 : _GEN_442; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_605 = opcode == 4'hf ? phv_data_120 : _GEN_443; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_606 = opcode == 4'hf ? phv_data_127 : _GEN_444; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_607 = opcode == 4'hf ? phv_data_126 : _GEN_445; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_608 = opcode == 4'hf ? phv_data_125 : _GEN_446; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_609 = opcode == 4'hf ? phv_data_124 : _GEN_447; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_610 = opcode == 4'hf ? phv_data_131 : _GEN_448; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_611 = opcode == 4'hf ? phv_data_130 : _GEN_449; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_612 = opcode == 4'hf ? phv_data_129 : _GEN_450; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_613 = opcode == 4'hf ? phv_data_128 : _GEN_451; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_614 = opcode == 4'hf ? phv_data_135 : _GEN_452; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_615 = opcode == 4'hf ? phv_data_134 : _GEN_453; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_616 = opcode == 4'hf ? phv_data_133 : _GEN_454; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_617 = opcode == 4'hf ? phv_data_132 : _GEN_455; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_618 = opcode == 4'hf ? phv_data_139 : _GEN_456; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_619 = opcode == 4'hf ? phv_data_138 : _GEN_457; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_620 = opcode == 4'hf ? phv_data_137 : _GEN_458; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_621 = opcode == 4'hf ? phv_data_136 : _GEN_459; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_622 = opcode == 4'hf ? phv_data_143 : _GEN_460; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_623 = opcode == 4'hf ? phv_data_142 : _GEN_461; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_624 = opcode == 4'hf ? phv_data_141 : _GEN_462; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_625 = opcode == 4'hf ? phv_data_140 : _GEN_463; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_626 = opcode == 4'hf ? phv_data_147 : _GEN_464; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_627 = opcode == 4'hf ? phv_data_146 : _GEN_465; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_628 = opcode == 4'hf ? phv_data_145 : _GEN_466; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_629 = opcode == 4'hf ? phv_data_144 : _GEN_467; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_630 = opcode == 4'hf ? phv_data_151 : _GEN_468; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_631 = opcode == 4'hf ? phv_data_150 : _GEN_469; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_632 = opcode == 4'hf ? phv_data_149 : _GEN_470; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_633 = opcode == 4'hf ? phv_data_148 : _GEN_471; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_634 = opcode == 4'hf ? phv_data_155 : _GEN_472; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_635 = opcode == 4'hf ? phv_data_154 : _GEN_473; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_636 = opcode == 4'hf ? phv_data_153 : _GEN_474; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_637 = opcode == 4'hf ? phv_data_152 : _GEN_475; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_638 = opcode == 4'hf ? phv_data_159 : _GEN_476; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_639 = opcode == 4'hf ? phv_data_158 : _GEN_477; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_640 = opcode == 4'hf ? phv_data_157 : _GEN_478; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_641 = opcode == 4'hf ? phv_data_156 : _GEN_479; // @[executor.scala 466:52 executor.scala 450:25]
  wire [3:0] opcode_1 = vliw_1[31:28]; // @[primitive.scala 9:44]
  wire [13:0] parameter_2_1 = vliw_1[13:0]; // @[primitive.scala 11:44]
  wire [7:0] _GEN_2770 = {{2'd0}, dst_offset_1}; // @[executor.scala 473:49]
  wire [7:0] byte_160 = field_1[7:0]; // @[executor.scala 475:56]
  wire [7:0] _GEN_642 = mask_1[0] ? byte_160 : _GEN_482; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] byte_161 = field_1[15:8]; // @[executor.scala 475:56]
  wire [7:0] _GEN_643 = mask_1[1] ? byte_161 : _GEN_483; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] byte_162 = field_1[23:16]; // @[executor.scala 475:56]
  wire [7:0] _GEN_644 = mask_1[2] ? byte_162 : _GEN_484; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] byte_163 = field_1[31:24]; // @[executor.scala 475:56]
  wire [7:0] _GEN_645 = mask_1[3] ? byte_163 : _GEN_485; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_646 = _GEN_2770 == 8'h0 ? _GEN_642 : _GEN_482; // @[executor.scala 473:84]
  wire [7:0] _GEN_647 = _GEN_2770 == 8'h0 ? _GEN_643 : _GEN_483; // @[executor.scala 473:84]
  wire [7:0] _GEN_648 = _GEN_2770 == 8'h0 ? _GEN_644 : _GEN_484; // @[executor.scala 473:84]
  wire [7:0] _GEN_649 = _GEN_2770 == 8'h0 ? _GEN_645 : _GEN_485; // @[executor.scala 473:84]
  wire [7:0] _GEN_650 = mask_1[0] ? byte_160 : _GEN_486; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_651 = mask_1[1] ? byte_161 : _GEN_487; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_652 = mask_1[2] ? byte_162 : _GEN_488; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_653 = mask_1[3] ? byte_163 : _GEN_489; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_654 = _GEN_2770 == 8'h1 ? _GEN_650 : _GEN_486; // @[executor.scala 473:84]
  wire [7:0] _GEN_655 = _GEN_2770 == 8'h1 ? _GEN_651 : _GEN_487; // @[executor.scala 473:84]
  wire [7:0] _GEN_656 = _GEN_2770 == 8'h1 ? _GEN_652 : _GEN_488; // @[executor.scala 473:84]
  wire [7:0] _GEN_657 = _GEN_2770 == 8'h1 ? _GEN_653 : _GEN_489; // @[executor.scala 473:84]
  wire [7:0] _GEN_658 = mask_1[0] ? byte_160 : _GEN_490; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_659 = mask_1[1] ? byte_161 : _GEN_491; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_660 = mask_1[2] ? byte_162 : _GEN_492; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_661 = mask_1[3] ? byte_163 : _GEN_493; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_662 = _GEN_2770 == 8'h2 ? _GEN_658 : _GEN_490; // @[executor.scala 473:84]
  wire [7:0] _GEN_663 = _GEN_2770 == 8'h2 ? _GEN_659 : _GEN_491; // @[executor.scala 473:84]
  wire [7:0] _GEN_664 = _GEN_2770 == 8'h2 ? _GEN_660 : _GEN_492; // @[executor.scala 473:84]
  wire [7:0] _GEN_665 = _GEN_2770 == 8'h2 ? _GEN_661 : _GEN_493; // @[executor.scala 473:84]
  wire [7:0] _GEN_666 = mask_1[0] ? byte_160 : _GEN_494; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_667 = mask_1[1] ? byte_161 : _GEN_495; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_668 = mask_1[2] ? byte_162 : _GEN_496; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_669 = mask_1[3] ? byte_163 : _GEN_497; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_670 = _GEN_2770 == 8'h3 ? _GEN_666 : _GEN_494; // @[executor.scala 473:84]
  wire [7:0] _GEN_671 = _GEN_2770 == 8'h3 ? _GEN_667 : _GEN_495; // @[executor.scala 473:84]
  wire [7:0] _GEN_672 = _GEN_2770 == 8'h3 ? _GEN_668 : _GEN_496; // @[executor.scala 473:84]
  wire [7:0] _GEN_673 = _GEN_2770 == 8'h3 ? _GEN_669 : _GEN_497; // @[executor.scala 473:84]
  wire [7:0] _GEN_674 = mask_1[0] ? byte_160 : _GEN_498; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_675 = mask_1[1] ? byte_161 : _GEN_499; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_676 = mask_1[2] ? byte_162 : _GEN_500; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_677 = mask_1[3] ? byte_163 : _GEN_501; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_678 = _GEN_2770 == 8'h4 ? _GEN_674 : _GEN_498; // @[executor.scala 473:84]
  wire [7:0] _GEN_679 = _GEN_2770 == 8'h4 ? _GEN_675 : _GEN_499; // @[executor.scala 473:84]
  wire [7:0] _GEN_680 = _GEN_2770 == 8'h4 ? _GEN_676 : _GEN_500; // @[executor.scala 473:84]
  wire [7:0] _GEN_681 = _GEN_2770 == 8'h4 ? _GEN_677 : _GEN_501; // @[executor.scala 473:84]
  wire [7:0] _GEN_682 = mask_1[0] ? byte_160 : _GEN_502; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_683 = mask_1[1] ? byte_161 : _GEN_503; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_684 = mask_1[2] ? byte_162 : _GEN_504; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_685 = mask_1[3] ? byte_163 : _GEN_505; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_686 = _GEN_2770 == 8'h5 ? _GEN_682 : _GEN_502; // @[executor.scala 473:84]
  wire [7:0] _GEN_687 = _GEN_2770 == 8'h5 ? _GEN_683 : _GEN_503; // @[executor.scala 473:84]
  wire [7:0] _GEN_688 = _GEN_2770 == 8'h5 ? _GEN_684 : _GEN_504; // @[executor.scala 473:84]
  wire [7:0] _GEN_689 = _GEN_2770 == 8'h5 ? _GEN_685 : _GEN_505; // @[executor.scala 473:84]
  wire [7:0] _GEN_690 = mask_1[0] ? byte_160 : _GEN_506; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_691 = mask_1[1] ? byte_161 : _GEN_507; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_692 = mask_1[2] ? byte_162 : _GEN_508; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_693 = mask_1[3] ? byte_163 : _GEN_509; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_694 = _GEN_2770 == 8'h6 ? _GEN_690 : _GEN_506; // @[executor.scala 473:84]
  wire [7:0] _GEN_695 = _GEN_2770 == 8'h6 ? _GEN_691 : _GEN_507; // @[executor.scala 473:84]
  wire [7:0] _GEN_696 = _GEN_2770 == 8'h6 ? _GEN_692 : _GEN_508; // @[executor.scala 473:84]
  wire [7:0] _GEN_697 = _GEN_2770 == 8'h6 ? _GEN_693 : _GEN_509; // @[executor.scala 473:84]
  wire [7:0] _GEN_698 = mask_1[0] ? byte_160 : _GEN_510; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_699 = mask_1[1] ? byte_161 : _GEN_511; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_700 = mask_1[2] ? byte_162 : _GEN_512; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_701 = mask_1[3] ? byte_163 : _GEN_513; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_702 = _GEN_2770 == 8'h7 ? _GEN_698 : _GEN_510; // @[executor.scala 473:84]
  wire [7:0] _GEN_703 = _GEN_2770 == 8'h7 ? _GEN_699 : _GEN_511; // @[executor.scala 473:84]
  wire [7:0] _GEN_704 = _GEN_2770 == 8'h7 ? _GEN_700 : _GEN_512; // @[executor.scala 473:84]
  wire [7:0] _GEN_705 = _GEN_2770 == 8'h7 ? _GEN_701 : _GEN_513; // @[executor.scala 473:84]
  wire [7:0] _GEN_706 = mask_1[0] ? byte_160 : _GEN_514; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_707 = mask_1[1] ? byte_161 : _GEN_515; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_708 = mask_1[2] ? byte_162 : _GEN_516; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_709 = mask_1[3] ? byte_163 : _GEN_517; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_710 = _GEN_2770 == 8'h8 ? _GEN_706 : _GEN_514; // @[executor.scala 473:84]
  wire [7:0] _GEN_711 = _GEN_2770 == 8'h8 ? _GEN_707 : _GEN_515; // @[executor.scala 473:84]
  wire [7:0] _GEN_712 = _GEN_2770 == 8'h8 ? _GEN_708 : _GEN_516; // @[executor.scala 473:84]
  wire [7:0] _GEN_713 = _GEN_2770 == 8'h8 ? _GEN_709 : _GEN_517; // @[executor.scala 473:84]
  wire [7:0] _GEN_714 = mask_1[0] ? byte_160 : _GEN_518; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_715 = mask_1[1] ? byte_161 : _GEN_519; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_716 = mask_1[2] ? byte_162 : _GEN_520; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_717 = mask_1[3] ? byte_163 : _GEN_521; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_718 = _GEN_2770 == 8'h9 ? _GEN_714 : _GEN_518; // @[executor.scala 473:84]
  wire [7:0] _GEN_719 = _GEN_2770 == 8'h9 ? _GEN_715 : _GEN_519; // @[executor.scala 473:84]
  wire [7:0] _GEN_720 = _GEN_2770 == 8'h9 ? _GEN_716 : _GEN_520; // @[executor.scala 473:84]
  wire [7:0] _GEN_721 = _GEN_2770 == 8'h9 ? _GEN_717 : _GEN_521; // @[executor.scala 473:84]
  wire [7:0] _GEN_722 = mask_1[0] ? byte_160 : _GEN_522; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_723 = mask_1[1] ? byte_161 : _GEN_523; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_724 = mask_1[2] ? byte_162 : _GEN_524; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_725 = mask_1[3] ? byte_163 : _GEN_525; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_726 = _GEN_2770 == 8'ha ? _GEN_722 : _GEN_522; // @[executor.scala 473:84]
  wire [7:0] _GEN_727 = _GEN_2770 == 8'ha ? _GEN_723 : _GEN_523; // @[executor.scala 473:84]
  wire [7:0] _GEN_728 = _GEN_2770 == 8'ha ? _GEN_724 : _GEN_524; // @[executor.scala 473:84]
  wire [7:0] _GEN_729 = _GEN_2770 == 8'ha ? _GEN_725 : _GEN_525; // @[executor.scala 473:84]
  wire [7:0] _GEN_730 = mask_1[0] ? byte_160 : _GEN_526; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_731 = mask_1[1] ? byte_161 : _GEN_527; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_732 = mask_1[2] ? byte_162 : _GEN_528; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_733 = mask_1[3] ? byte_163 : _GEN_529; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_734 = _GEN_2770 == 8'hb ? _GEN_730 : _GEN_526; // @[executor.scala 473:84]
  wire [7:0] _GEN_735 = _GEN_2770 == 8'hb ? _GEN_731 : _GEN_527; // @[executor.scala 473:84]
  wire [7:0] _GEN_736 = _GEN_2770 == 8'hb ? _GEN_732 : _GEN_528; // @[executor.scala 473:84]
  wire [7:0] _GEN_737 = _GEN_2770 == 8'hb ? _GEN_733 : _GEN_529; // @[executor.scala 473:84]
  wire [7:0] _GEN_738 = mask_1[0] ? byte_160 : _GEN_530; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_739 = mask_1[1] ? byte_161 : _GEN_531; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_740 = mask_1[2] ? byte_162 : _GEN_532; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_741 = mask_1[3] ? byte_163 : _GEN_533; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_742 = _GEN_2770 == 8'hc ? _GEN_738 : _GEN_530; // @[executor.scala 473:84]
  wire [7:0] _GEN_743 = _GEN_2770 == 8'hc ? _GEN_739 : _GEN_531; // @[executor.scala 473:84]
  wire [7:0] _GEN_744 = _GEN_2770 == 8'hc ? _GEN_740 : _GEN_532; // @[executor.scala 473:84]
  wire [7:0] _GEN_745 = _GEN_2770 == 8'hc ? _GEN_741 : _GEN_533; // @[executor.scala 473:84]
  wire [7:0] _GEN_746 = mask_1[0] ? byte_160 : _GEN_534; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_747 = mask_1[1] ? byte_161 : _GEN_535; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_748 = mask_1[2] ? byte_162 : _GEN_536; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_749 = mask_1[3] ? byte_163 : _GEN_537; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_750 = _GEN_2770 == 8'hd ? _GEN_746 : _GEN_534; // @[executor.scala 473:84]
  wire [7:0] _GEN_751 = _GEN_2770 == 8'hd ? _GEN_747 : _GEN_535; // @[executor.scala 473:84]
  wire [7:0] _GEN_752 = _GEN_2770 == 8'hd ? _GEN_748 : _GEN_536; // @[executor.scala 473:84]
  wire [7:0] _GEN_753 = _GEN_2770 == 8'hd ? _GEN_749 : _GEN_537; // @[executor.scala 473:84]
  wire [7:0] _GEN_754 = mask_1[0] ? byte_160 : _GEN_538; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_755 = mask_1[1] ? byte_161 : _GEN_539; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_756 = mask_1[2] ? byte_162 : _GEN_540; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_757 = mask_1[3] ? byte_163 : _GEN_541; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_758 = _GEN_2770 == 8'he ? _GEN_754 : _GEN_538; // @[executor.scala 473:84]
  wire [7:0] _GEN_759 = _GEN_2770 == 8'he ? _GEN_755 : _GEN_539; // @[executor.scala 473:84]
  wire [7:0] _GEN_760 = _GEN_2770 == 8'he ? _GEN_756 : _GEN_540; // @[executor.scala 473:84]
  wire [7:0] _GEN_761 = _GEN_2770 == 8'he ? _GEN_757 : _GEN_541; // @[executor.scala 473:84]
  wire [7:0] _GEN_762 = mask_1[0] ? byte_160 : _GEN_542; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_763 = mask_1[1] ? byte_161 : _GEN_543; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_764 = mask_1[2] ? byte_162 : _GEN_544; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_765 = mask_1[3] ? byte_163 : _GEN_545; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_766 = _GEN_2770 == 8'hf ? _GEN_762 : _GEN_542; // @[executor.scala 473:84]
  wire [7:0] _GEN_767 = _GEN_2770 == 8'hf ? _GEN_763 : _GEN_543; // @[executor.scala 473:84]
  wire [7:0] _GEN_768 = _GEN_2770 == 8'hf ? _GEN_764 : _GEN_544; // @[executor.scala 473:84]
  wire [7:0] _GEN_769 = _GEN_2770 == 8'hf ? _GEN_765 : _GEN_545; // @[executor.scala 473:84]
  wire [7:0] _GEN_770 = mask_1[0] ? byte_160 : _GEN_546; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_771 = mask_1[1] ? byte_161 : _GEN_547; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_772 = mask_1[2] ? byte_162 : _GEN_548; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_773 = mask_1[3] ? byte_163 : _GEN_549; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_774 = _GEN_2770 == 8'h10 ? _GEN_770 : _GEN_546; // @[executor.scala 473:84]
  wire [7:0] _GEN_775 = _GEN_2770 == 8'h10 ? _GEN_771 : _GEN_547; // @[executor.scala 473:84]
  wire [7:0] _GEN_776 = _GEN_2770 == 8'h10 ? _GEN_772 : _GEN_548; // @[executor.scala 473:84]
  wire [7:0] _GEN_777 = _GEN_2770 == 8'h10 ? _GEN_773 : _GEN_549; // @[executor.scala 473:84]
  wire [7:0] _GEN_778 = mask_1[0] ? byte_160 : _GEN_550; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_779 = mask_1[1] ? byte_161 : _GEN_551; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_780 = mask_1[2] ? byte_162 : _GEN_552; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_781 = mask_1[3] ? byte_163 : _GEN_553; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_782 = _GEN_2770 == 8'h11 ? _GEN_778 : _GEN_550; // @[executor.scala 473:84]
  wire [7:0] _GEN_783 = _GEN_2770 == 8'h11 ? _GEN_779 : _GEN_551; // @[executor.scala 473:84]
  wire [7:0] _GEN_784 = _GEN_2770 == 8'h11 ? _GEN_780 : _GEN_552; // @[executor.scala 473:84]
  wire [7:0] _GEN_785 = _GEN_2770 == 8'h11 ? _GEN_781 : _GEN_553; // @[executor.scala 473:84]
  wire [7:0] _GEN_786 = mask_1[0] ? byte_160 : _GEN_554; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_787 = mask_1[1] ? byte_161 : _GEN_555; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_788 = mask_1[2] ? byte_162 : _GEN_556; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_789 = mask_1[3] ? byte_163 : _GEN_557; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_790 = _GEN_2770 == 8'h12 ? _GEN_786 : _GEN_554; // @[executor.scala 473:84]
  wire [7:0] _GEN_791 = _GEN_2770 == 8'h12 ? _GEN_787 : _GEN_555; // @[executor.scala 473:84]
  wire [7:0] _GEN_792 = _GEN_2770 == 8'h12 ? _GEN_788 : _GEN_556; // @[executor.scala 473:84]
  wire [7:0] _GEN_793 = _GEN_2770 == 8'h12 ? _GEN_789 : _GEN_557; // @[executor.scala 473:84]
  wire [7:0] _GEN_794 = mask_1[0] ? byte_160 : _GEN_558; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_795 = mask_1[1] ? byte_161 : _GEN_559; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_796 = mask_1[2] ? byte_162 : _GEN_560; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_797 = mask_1[3] ? byte_163 : _GEN_561; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_798 = _GEN_2770 == 8'h13 ? _GEN_794 : _GEN_558; // @[executor.scala 473:84]
  wire [7:0] _GEN_799 = _GEN_2770 == 8'h13 ? _GEN_795 : _GEN_559; // @[executor.scala 473:84]
  wire [7:0] _GEN_800 = _GEN_2770 == 8'h13 ? _GEN_796 : _GEN_560; // @[executor.scala 473:84]
  wire [7:0] _GEN_801 = _GEN_2770 == 8'h13 ? _GEN_797 : _GEN_561; // @[executor.scala 473:84]
  wire [7:0] _GEN_802 = mask_1[0] ? byte_160 : _GEN_562; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_803 = mask_1[1] ? byte_161 : _GEN_563; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_804 = mask_1[2] ? byte_162 : _GEN_564; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_805 = mask_1[3] ? byte_163 : _GEN_565; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_806 = _GEN_2770 == 8'h14 ? _GEN_802 : _GEN_562; // @[executor.scala 473:84]
  wire [7:0] _GEN_807 = _GEN_2770 == 8'h14 ? _GEN_803 : _GEN_563; // @[executor.scala 473:84]
  wire [7:0] _GEN_808 = _GEN_2770 == 8'h14 ? _GEN_804 : _GEN_564; // @[executor.scala 473:84]
  wire [7:0] _GEN_809 = _GEN_2770 == 8'h14 ? _GEN_805 : _GEN_565; // @[executor.scala 473:84]
  wire [7:0] _GEN_810 = mask_1[0] ? byte_160 : _GEN_566; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_811 = mask_1[1] ? byte_161 : _GEN_567; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_812 = mask_1[2] ? byte_162 : _GEN_568; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_813 = mask_1[3] ? byte_163 : _GEN_569; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_814 = _GEN_2770 == 8'h15 ? _GEN_810 : _GEN_566; // @[executor.scala 473:84]
  wire [7:0] _GEN_815 = _GEN_2770 == 8'h15 ? _GEN_811 : _GEN_567; // @[executor.scala 473:84]
  wire [7:0] _GEN_816 = _GEN_2770 == 8'h15 ? _GEN_812 : _GEN_568; // @[executor.scala 473:84]
  wire [7:0] _GEN_817 = _GEN_2770 == 8'h15 ? _GEN_813 : _GEN_569; // @[executor.scala 473:84]
  wire [7:0] _GEN_818 = mask_1[0] ? byte_160 : _GEN_570; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_819 = mask_1[1] ? byte_161 : _GEN_571; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_820 = mask_1[2] ? byte_162 : _GEN_572; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_821 = mask_1[3] ? byte_163 : _GEN_573; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_822 = _GEN_2770 == 8'h16 ? _GEN_818 : _GEN_570; // @[executor.scala 473:84]
  wire [7:0] _GEN_823 = _GEN_2770 == 8'h16 ? _GEN_819 : _GEN_571; // @[executor.scala 473:84]
  wire [7:0] _GEN_824 = _GEN_2770 == 8'h16 ? _GEN_820 : _GEN_572; // @[executor.scala 473:84]
  wire [7:0] _GEN_825 = _GEN_2770 == 8'h16 ? _GEN_821 : _GEN_573; // @[executor.scala 473:84]
  wire [7:0] _GEN_826 = mask_1[0] ? byte_160 : _GEN_574; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_827 = mask_1[1] ? byte_161 : _GEN_575; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_828 = mask_1[2] ? byte_162 : _GEN_576; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_829 = mask_1[3] ? byte_163 : _GEN_577; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_830 = _GEN_2770 == 8'h17 ? _GEN_826 : _GEN_574; // @[executor.scala 473:84]
  wire [7:0] _GEN_831 = _GEN_2770 == 8'h17 ? _GEN_827 : _GEN_575; // @[executor.scala 473:84]
  wire [7:0] _GEN_832 = _GEN_2770 == 8'h17 ? _GEN_828 : _GEN_576; // @[executor.scala 473:84]
  wire [7:0] _GEN_833 = _GEN_2770 == 8'h17 ? _GEN_829 : _GEN_577; // @[executor.scala 473:84]
  wire [7:0] _GEN_834 = mask_1[0] ? byte_160 : _GEN_578; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_835 = mask_1[1] ? byte_161 : _GEN_579; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_836 = mask_1[2] ? byte_162 : _GEN_580; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_837 = mask_1[3] ? byte_163 : _GEN_581; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_838 = _GEN_2770 == 8'h18 ? _GEN_834 : _GEN_578; // @[executor.scala 473:84]
  wire [7:0] _GEN_839 = _GEN_2770 == 8'h18 ? _GEN_835 : _GEN_579; // @[executor.scala 473:84]
  wire [7:0] _GEN_840 = _GEN_2770 == 8'h18 ? _GEN_836 : _GEN_580; // @[executor.scala 473:84]
  wire [7:0] _GEN_841 = _GEN_2770 == 8'h18 ? _GEN_837 : _GEN_581; // @[executor.scala 473:84]
  wire [7:0] _GEN_842 = mask_1[0] ? byte_160 : _GEN_582; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_843 = mask_1[1] ? byte_161 : _GEN_583; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_844 = mask_1[2] ? byte_162 : _GEN_584; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_845 = mask_1[3] ? byte_163 : _GEN_585; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_846 = _GEN_2770 == 8'h19 ? _GEN_842 : _GEN_582; // @[executor.scala 473:84]
  wire [7:0] _GEN_847 = _GEN_2770 == 8'h19 ? _GEN_843 : _GEN_583; // @[executor.scala 473:84]
  wire [7:0] _GEN_848 = _GEN_2770 == 8'h19 ? _GEN_844 : _GEN_584; // @[executor.scala 473:84]
  wire [7:0] _GEN_849 = _GEN_2770 == 8'h19 ? _GEN_845 : _GEN_585; // @[executor.scala 473:84]
  wire [7:0] _GEN_850 = mask_1[0] ? byte_160 : _GEN_586; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_851 = mask_1[1] ? byte_161 : _GEN_587; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_852 = mask_1[2] ? byte_162 : _GEN_588; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_853 = mask_1[3] ? byte_163 : _GEN_589; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_854 = _GEN_2770 == 8'h1a ? _GEN_850 : _GEN_586; // @[executor.scala 473:84]
  wire [7:0] _GEN_855 = _GEN_2770 == 8'h1a ? _GEN_851 : _GEN_587; // @[executor.scala 473:84]
  wire [7:0] _GEN_856 = _GEN_2770 == 8'h1a ? _GEN_852 : _GEN_588; // @[executor.scala 473:84]
  wire [7:0] _GEN_857 = _GEN_2770 == 8'h1a ? _GEN_853 : _GEN_589; // @[executor.scala 473:84]
  wire [7:0] _GEN_858 = mask_1[0] ? byte_160 : _GEN_590; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_859 = mask_1[1] ? byte_161 : _GEN_591; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_860 = mask_1[2] ? byte_162 : _GEN_592; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_861 = mask_1[3] ? byte_163 : _GEN_593; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_862 = _GEN_2770 == 8'h1b ? _GEN_858 : _GEN_590; // @[executor.scala 473:84]
  wire [7:0] _GEN_863 = _GEN_2770 == 8'h1b ? _GEN_859 : _GEN_591; // @[executor.scala 473:84]
  wire [7:0] _GEN_864 = _GEN_2770 == 8'h1b ? _GEN_860 : _GEN_592; // @[executor.scala 473:84]
  wire [7:0] _GEN_865 = _GEN_2770 == 8'h1b ? _GEN_861 : _GEN_593; // @[executor.scala 473:84]
  wire [7:0] _GEN_866 = mask_1[0] ? byte_160 : _GEN_594; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_867 = mask_1[1] ? byte_161 : _GEN_595; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_868 = mask_1[2] ? byte_162 : _GEN_596; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_869 = mask_1[3] ? byte_163 : _GEN_597; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_870 = _GEN_2770 == 8'h1c ? _GEN_866 : _GEN_594; // @[executor.scala 473:84]
  wire [7:0] _GEN_871 = _GEN_2770 == 8'h1c ? _GEN_867 : _GEN_595; // @[executor.scala 473:84]
  wire [7:0] _GEN_872 = _GEN_2770 == 8'h1c ? _GEN_868 : _GEN_596; // @[executor.scala 473:84]
  wire [7:0] _GEN_873 = _GEN_2770 == 8'h1c ? _GEN_869 : _GEN_597; // @[executor.scala 473:84]
  wire [7:0] _GEN_874 = mask_1[0] ? byte_160 : _GEN_598; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_875 = mask_1[1] ? byte_161 : _GEN_599; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_876 = mask_1[2] ? byte_162 : _GEN_600; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_877 = mask_1[3] ? byte_163 : _GEN_601; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_878 = _GEN_2770 == 8'h1d ? _GEN_874 : _GEN_598; // @[executor.scala 473:84]
  wire [7:0] _GEN_879 = _GEN_2770 == 8'h1d ? _GEN_875 : _GEN_599; // @[executor.scala 473:84]
  wire [7:0] _GEN_880 = _GEN_2770 == 8'h1d ? _GEN_876 : _GEN_600; // @[executor.scala 473:84]
  wire [7:0] _GEN_881 = _GEN_2770 == 8'h1d ? _GEN_877 : _GEN_601; // @[executor.scala 473:84]
  wire [7:0] _GEN_882 = mask_1[0] ? byte_160 : _GEN_602; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_883 = mask_1[1] ? byte_161 : _GEN_603; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_884 = mask_1[2] ? byte_162 : _GEN_604; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_885 = mask_1[3] ? byte_163 : _GEN_605; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_886 = _GEN_2770 == 8'h1e ? _GEN_882 : _GEN_602; // @[executor.scala 473:84]
  wire [7:0] _GEN_887 = _GEN_2770 == 8'h1e ? _GEN_883 : _GEN_603; // @[executor.scala 473:84]
  wire [7:0] _GEN_888 = _GEN_2770 == 8'h1e ? _GEN_884 : _GEN_604; // @[executor.scala 473:84]
  wire [7:0] _GEN_889 = _GEN_2770 == 8'h1e ? _GEN_885 : _GEN_605; // @[executor.scala 473:84]
  wire [7:0] _GEN_890 = mask_1[0] ? byte_160 : _GEN_606; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_891 = mask_1[1] ? byte_161 : _GEN_607; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_892 = mask_1[2] ? byte_162 : _GEN_608; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_893 = mask_1[3] ? byte_163 : _GEN_609; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_894 = _GEN_2770 == 8'h1f ? _GEN_890 : _GEN_606; // @[executor.scala 473:84]
  wire [7:0] _GEN_895 = _GEN_2770 == 8'h1f ? _GEN_891 : _GEN_607; // @[executor.scala 473:84]
  wire [7:0] _GEN_896 = _GEN_2770 == 8'h1f ? _GEN_892 : _GEN_608; // @[executor.scala 473:84]
  wire [7:0] _GEN_897 = _GEN_2770 == 8'h1f ? _GEN_893 : _GEN_609; // @[executor.scala 473:84]
  wire [7:0] _GEN_898 = mask_1[0] ? byte_160 : _GEN_610; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_899 = mask_1[1] ? byte_161 : _GEN_611; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_900 = mask_1[2] ? byte_162 : _GEN_612; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_901 = mask_1[3] ? byte_163 : _GEN_613; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_902 = _GEN_2770 == 8'h20 ? _GEN_898 : _GEN_610; // @[executor.scala 473:84]
  wire [7:0] _GEN_903 = _GEN_2770 == 8'h20 ? _GEN_899 : _GEN_611; // @[executor.scala 473:84]
  wire [7:0] _GEN_904 = _GEN_2770 == 8'h20 ? _GEN_900 : _GEN_612; // @[executor.scala 473:84]
  wire [7:0] _GEN_905 = _GEN_2770 == 8'h20 ? _GEN_901 : _GEN_613; // @[executor.scala 473:84]
  wire [7:0] _GEN_906 = mask_1[0] ? byte_160 : _GEN_614; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_907 = mask_1[1] ? byte_161 : _GEN_615; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_908 = mask_1[2] ? byte_162 : _GEN_616; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_909 = mask_1[3] ? byte_163 : _GEN_617; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_910 = _GEN_2770 == 8'h21 ? _GEN_906 : _GEN_614; // @[executor.scala 473:84]
  wire [7:0] _GEN_911 = _GEN_2770 == 8'h21 ? _GEN_907 : _GEN_615; // @[executor.scala 473:84]
  wire [7:0] _GEN_912 = _GEN_2770 == 8'h21 ? _GEN_908 : _GEN_616; // @[executor.scala 473:84]
  wire [7:0] _GEN_913 = _GEN_2770 == 8'h21 ? _GEN_909 : _GEN_617; // @[executor.scala 473:84]
  wire [7:0] _GEN_914 = mask_1[0] ? byte_160 : _GEN_618; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_915 = mask_1[1] ? byte_161 : _GEN_619; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_916 = mask_1[2] ? byte_162 : _GEN_620; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_917 = mask_1[3] ? byte_163 : _GEN_621; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_918 = _GEN_2770 == 8'h22 ? _GEN_914 : _GEN_618; // @[executor.scala 473:84]
  wire [7:0] _GEN_919 = _GEN_2770 == 8'h22 ? _GEN_915 : _GEN_619; // @[executor.scala 473:84]
  wire [7:0] _GEN_920 = _GEN_2770 == 8'h22 ? _GEN_916 : _GEN_620; // @[executor.scala 473:84]
  wire [7:0] _GEN_921 = _GEN_2770 == 8'h22 ? _GEN_917 : _GEN_621; // @[executor.scala 473:84]
  wire [7:0] _GEN_922 = mask_1[0] ? byte_160 : _GEN_622; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_923 = mask_1[1] ? byte_161 : _GEN_623; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_924 = mask_1[2] ? byte_162 : _GEN_624; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_925 = mask_1[3] ? byte_163 : _GEN_625; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_926 = _GEN_2770 == 8'h23 ? _GEN_922 : _GEN_622; // @[executor.scala 473:84]
  wire [7:0] _GEN_927 = _GEN_2770 == 8'h23 ? _GEN_923 : _GEN_623; // @[executor.scala 473:84]
  wire [7:0] _GEN_928 = _GEN_2770 == 8'h23 ? _GEN_924 : _GEN_624; // @[executor.scala 473:84]
  wire [7:0] _GEN_929 = _GEN_2770 == 8'h23 ? _GEN_925 : _GEN_625; // @[executor.scala 473:84]
  wire [7:0] _GEN_930 = mask_1[0] ? byte_160 : _GEN_626; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_931 = mask_1[1] ? byte_161 : _GEN_627; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_932 = mask_1[2] ? byte_162 : _GEN_628; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_933 = mask_1[3] ? byte_163 : _GEN_629; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_934 = _GEN_2770 == 8'h24 ? _GEN_930 : _GEN_626; // @[executor.scala 473:84]
  wire [7:0] _GEN_935 = _GEN_2770 == 8'h24 ? _GEN_931 : _GEN_627; // @[executor.scala 473:84]
  wire [7:0] _GEN_936 = _GEN_2770 == 8'h24 ? _GEN_932 : _GEN_628; // @[executor.scala 473:84]
  wire [7:0] _GEN_937 = _GEN_2770 == 8'h24 ? _GEN_933 : _GEN_629; // @[executor.scala 473:84]
  wire [7:0] _GEN_938 = mask_1[0] ? byte_160 : _GEN_630; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_939 = mask_1[1] ? byte_161 : _GEN_631; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_940 = mask_1[2] ? byte_162 : _GEN_632; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_941 = mask_1[3] ? byte_163 : _GEN_633; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_942 = _GEN_2770 == 8'h25 ? _GEN_938 : _GEN_630; // @[executor.scala 473:84]
  wire [7:0] _GEN_943 = _GEN_2770 == 8'h25 ? _GEN_939 : _GEN_631; // @[executor.scala 473:84]
  wire [7:0] _GEN_944 = _GEN_2770 == 8'h25 ? _GEN_940 : _GEN_632; // @[executor.scala 473:84]
  wire [7:0] _GEN_945 = _GEN_2770 == 8'h25 ? _GEN_941 : _GEN_633; // @[executor.scala 473:84]
  wire [7:0] _GEN_946 = mask_1[0] ? byte_160 : _GEN_634; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_947 = mask_1[1] ? byte_161 : _GEN_635; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_948 = mask_1[2] ? byte_162 : _GEN_636; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_949 = mask_1[3] ? byte_163 : _GEN_637; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_950 = _GEN_2770 == 8'h26 ? _GEN_946 : _GEN_634; // @[executor.scala 473:84]
  wire [7:0] _GEN_951 = _GEN_2770 == 8'h26 ? _GEN_947 : _GEN_635; // @[executor.scala 473:84]
  wire [7:0] _GEN_952 = _GEN_2770 == 8'h26 ? _GEN_948 : _GEN_636; // @[executor.scala 473:84]
  wire [7:0] _GEN_953 = _GEN_2770 == 8'h26 ? _GEN_949 : _GEN_637; // @[executor.scala 473:84]
  wire [7:0] _GEN_954 = mask_1[0] ? byte_160 : _GEN_638; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_955 = mask_1[1] ? byte_161 : _GEN_639; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_956 = mask_1[2] ? byte_162 : _GEN_640; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_957 = mask_1[3] ? byte_163 : _GEN_641; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_958 = _GEN_2770 == 8'h27 ? _GEN_954 : _GEN_638; // @[executor.scala 473:84]
  wire [7:0] _GEN_959 = _GEN_2770 == 8'h27 ? _GEN_955 : _GEN_639; // @[executor.scala 473:84]
  wire [7:0] _GEN_960 = _GEN_2770 == 8'h27 ? _GEN_956 : _GEN_640; // @[executor.scala 473:84]
  wire [7:0] _GEN_961 = _GEN_2770 == 8'h27 ? _GEN_957 : _GEN_641; // @[executor.scala 473:84]
  wire [7:0] _GEN_962 = opcode_1 != 4'h0 ? _GEN_646 : _GEN_482; // @[executor.scala 470:55]
  wire [7:0] _GEN_963 = opcode_1 != 4'h0 ? _GEN_647 : _GEN_483; // @[executor.scala 470:55]
  wire [7:0] _GEN_964 = opcode_1 != 4'h0 ? _GEN_648 : _GEN_484; // @[executor.scala 470:55]
  wire [7:0] _GEN_965 = opcode_1 != 4'h0 ? _GEN_649 : _GEN_485; // @[executor.scala 470:55]
  wire [7:0] _GEN_966 = opcode_1 != 4'h0 ? _GEN_654 : _GEN_486; // @[executor.scala 470:55]
  wire [7:0] _GEN_967 = opcode_1 != 4'h0 ? _GEN_655 : _GEN_487; // @[executor.scala 470:55]
  wire [7:0] _GEN_968 = opcode_1 != 4'h0 ? _GEN_656 : _GEN_488; // @[executor.scala 470:55]
  wire [7:0] _GEN_969 = opcode_1 != 4'h0 ? _GEN_657 : _GEN_489; // @[executor.scala 470:55]
  wire [7:0] _GEN_970 = opcode_1 != 4'h0 ? _GEN_662 : _GEN_490; // @[executor.scala 470:55]
  wire [7:0] _GEN_971 = opcode_1 != 4'h0 ? _GEN_663 : _GEN_491; // @[executor.scala 470:55]
  wire [7:0] _GEN_972 = opcode_1 != 4'h0 ? _GEN_664 : _GEN_492; // @[executor.scala 470:55]
  wire [7:0] _GEN_973 = opcode_1 != 4'h0 ? _GEN_665 : _GEN_493; // @[executor.scala 470:55]
  wire [7:0] _GEN_974 = opcode_1 != 4'h0 ? _GEN_670 : _GEN_494; // @[executor.scala 470:55]
  wire [7:0] _GEN_975 = opcode_1 != 4'h0 ? _GEN_671 : _GEN_495; // @[executor.scala 470:55]
  wire [7:0] _GEN_976 = opcode_1 != 4'h0 ? _GEN_672 : _GEN_496; // @[executor.scala 470:55]
  wire [7:0] _GEN_977 = opcode_1 != 4'h0 ? _GEN_673 : _GEN_497; // @[executor.scala 470:55]
  wire [7:0] _GEN_978 = opcode_1 != 4'h0 ? _GEN_678 : _GEN_498; // @[executor.scala 470:55]
  wire [7:0] _GEN_979 = opcode_1 != 4'h0 ? _GEN_679 : _GEN_499; // @[executor.scala 470:55]
  wire [7:0] _GEN_980 = opcode_1 != 4'h0 ? _GEN_680 : _GEN_500; // @[executor.scala 470:55]
  wire [7:0] _GEN_981 = opcode_1 != 4'h0 ? _GEN_681 : _GEN_501; // @[executor.scala 470:55]
  wire [7:0] _GEN_982 = opcode_1 != 4'h0 ? _GEN_686 : _GEN_502; // @[executor.scala 470:55]
  wire [7:0] _GEN_983 = opcode_1 != 4'h0 ? _GEN_687 : _GEN_503; // @[executor.scala 470:55]
  wire [7:0] _GEN_984 = opcode_1 != 4'h0 ? _GEN_688 : _GEN_504; // @[executor.scala 470:55]
  wire [7:0] _GEN_985 = opcode_1 != 4'h0 ? _GEN_689 : _GEN_505; // @[executor.scala 470:55]
  wire [7:0] _GEN_986 = opcode_1 != 4'h0 ? _GEN_694 : _GEN_506; // @[executor.scala 470:55]
  wire [7:0] _GEN_987 = opcode_1 != 4'h0 ? _GEN_695 : _GEN_507; // @[executor.scala 470:55]
  wire [7:0] _GEN_988 = opcode_1 != 4'h0 ? _GEN_696 : _GEN_508; // @[executor.scala 470:55]
  wire [7:0] _GEN_989 = opcode_1 != 4'h0 ? _GEN_697 : _GEN_509; // @[executor.scala 470:55]
  wire [7:0] _GEN_990 = opcode_1 != 4'h0 ? _GEN_702 : _GEN_510; // @[executor.scala 470:55]
  wire [7:0] _GEN_991 = opcode_1 != 4'h0 ? _GEN_703 : _GEN_511; // @[executor.scala 470:55]
  wire [7:0] _GEN_992 = opcode_1 != 4'h0 ? _GEN_704 : _GEN_512; // @[executor.scala 470:55]
  wire [7:0] _GEN_993 = opcode_1 != 4'h0 ? _GEN_705 : _GEN_513; // @[executor.scala 470:55]
  wire [7:0] _GEN_994 = opcode_1 != 4'h0 ? _GEN_710 : _GEN_514; // @[executor.scala 470:55]
  wire [7:0] _GEN_995 = opcode_1 != 4'h0 ? _GEN_711 : _GEN_515; // @[executor.scala 470:55]
  wire [7:0] _GEN_996 = opcode_1 != 4'h0 ? _GEN_712 : _GEN_516; // @[executor.scala 470:55]
  wire [7:0] _GEN_997 = opcode_1 != 4'h0 ? _GEN_713 : _GEN_517; // @[executor.scala 470:55]
  wire [7:0] _GEN_998 = opcode_1 != 4'h0 ? _GEN_718 : _GEN_518; // @[executor.scala 470:55]
  wire [7:0] _GEN_999 = opcode_1 != 4'h0 ? _GEN_719 : _GEN_519; // @[executor.scala 470:55]
  wire [7:0] _GEN_1000 = opcode_1 != 4'h0 ? _GEN_720 : _GEN_520; // @[executor.scala 470:55]
  wire [7:0] _GEN_1001 = opcode_1 != 4'h0 ? _GEN_721 : _GEN_521; // @[executor.scala 470:55]
  wire [7:0] _GEN_1002 = opcode_1 != 4'h0 ? _GEN_726 : _GEN_522; // @[executor.scala 470:55]
  wire [7:0] _GEN_1003 = opcode_1 != 4'h0 ? _GEN_727 : _GEN_523; // @[executor.scala 470:55]
  wire [7:0] _GEN_1004 = opcode_1 != 4'h0 ? _GEN_728 : _GEN_524; // @[executor.scala 470:55]
  wire [7:0] _GEN_1005 = opcode_1 != 4'h0 ? _GEN_729 : _GEN_525; // @[executor.scala 470:55]
  wire [7:0] _GEN_1006 = opcode_1 != 4'h0 ? _GEN_734 : _GEN_526; // @[executor.scala 470:55]
  wire [7:0] _GEN_1007 = opcode_1 != 4'h0 ? _GEN_735 : _GEN_527; // @[executor.scala 470:55]
  wire [7:0] _GEN_1008 = opcode_1 != 4'h0 ? _GEN_736 : _GEN_528; // @[executor.scala 470:55]
  wire [7:0] _GEN_1009 = opcode_1 != 4'h0 ? _GEN_737 : _GEN_529; // @[executor.scala 470:55]
  wire [7:0] _GEN_1010 = opcode_1 != 4'h0 ? _GEN_742 : _GEN_530; // @[executor.scala 470:55]
  wire [7:0] _GEN_1011 = opcode_1 != 4'h0 ? _GEN_743 : _GEN_531; // @[executor.scala 470:55]
  wire [7:0] _GEN_1012 = opcode_1 != 4'h0 ? _GEN_744 : _GEN_532; // @[executor.scala 470:55]
  wire [7:0] _GEN_1013 = opcode_1 != 4'h0 ? _GEN_745 : _GEN_533; // @[executor.scala 470:55]
  wire [7:0] _GEN_1014 = opcode_1 != 4'h0 ? _GEN_750 : _GEN_534; // @[executor.scala 470:55]
  wire [7:0] _GEN_1015 = opcode_1 != 4'h0 ? _GEN_751 : _GEN_535; // @[executor.scala 470:55]
  wire [7:0] _GEN_1016 = opcode_1 != 4'h0 ? _GEN_752 : _GEN_536; // @[executor.scala 470:55]
  wire [7:0] _GEN_1017 = opcode_1 != 4'h0 ? _GEN_753 : _GEN_537; // @[executor.scala 470:55]
  wire [7:0] _GEN_1018 = opcode_1 != 4'h0 ? _GEN_758 : _GEN_538; // @[executor.scala 470:55]
  wire [7:0] _GEN_1019 = opcode_1 != 4'h0 ? _GEN_759 : _GEN_539; // @[executor.scala 470:55]
  wire [7:0] _GEN_1020 = opcode_1 != 4'h0 ? _GEN_760 : _GEN_540; // @[executor.scala 470:55]
  wire [7:0] _GEN_1021 = opcode_1 != 4'h0 ? _GEN_761 : _GEN_541; // @[executor.scala 470:55]
  wire [7:0] _GEN_1022 = opcode_1 != 4'h0 ? _GEN_766 : _GEN_542; // @[executor.scala 470:55]
  wire [7:0] _GEN_1023 = opcode_1 != 4'h0 ? _GEN_767 : _GEN_543; // @[executor.scala 470:55]
  wire [7:0] _GEN_1024 = opcode_1 != 4'h0 ? _GEN_768 : _GEN_544; // @[executor.scala 470:55]
  wire [7:0] _GEN_1025 = opcode_1 != 4'h0 ? _GEN_769 : _GEN_545; // @[executor.scala 470:55]
  wire [7:0] _GEN_1026 = opcode_1 != 4'h0 ? _GEN_774 : _GEN_546; // @[executor.scala 470:55]
  wire [7:0] _GEN_1027 = opcode_1 != 4'h0 ? _GEN_775 : _GEN_547; // @[executor.scala 470:55]
  wire [7:0] _GEN_1028 = opcode_1 != 4'h0 ? _GEN_776 : _GEN_548; // @[executor.scala 470:55]
  wire [7:0] _GEN_1029 = opcode_1 != 4'h0 ? _GEN_777 : _GEN_549; // @[executor.scala 470:55]
  wire [7:0] _GEN_1030 = opcode_1 != 4'h0 ? _GEN_782 : _GEN_550; // @[executor.scala 470:55]
  wire [7:0] _GEN_1031 = opcode_1 != 4'h0 ? _GEN_783 : _GEN_551; // @[executor.scala 470:55]
  wire [7:0] _GEN_1032 = opcode_1 != 4'h0 ? _GEN_784 : _GEN_552; // @[executor.scala 470:55]
  wire [7:0] _GEN_1033 = opcode_1 != 4'h0 ? _GEN_785 : _GEN_553; // @[executor.scala 470:55]
  wire [7:0] _GEN_1034 = opcode_1 != 4'h0 ? _GEN_790 : _GEN_554; // @[executor.scala 470:55]
  wire [7:0] _GEN_1035 = opcode_1 != 4'h0 ? _GEN_791 : _GEN_555; // @[executor.scala 470:55]
  wire [7:0] _GEN_1036 = opcode_1 != 4'h0 ? _GEN_792 : _GEN_556; // @[executor.scala 470:55]
  wire [7:0] _GEN_1037 = opcode_1 != 4'h0 ? _GEN_793 : _GEN_557; // @[executor.scala 470:55]
  wire [7:0] _GEN_1038 = opcode_1 != 4'h0 ? _GEN_798 : _GEN_558; // @[executor.scala 470:55]
  wire [7:0] _GEN_1039 = opcode_1 != 4'h0 ? _GEN_799 : _GEN_559; // @[executor.scala 470:55]
  wire [7:0] _GEN_1040 = opcode_1 != 4'h0 ? _GEN_800 : _GEN_560; // @[executor.scala 470:55]
  wire [7:0] _GEN_1041 = opcode_1 != 4'h0 ? _GEN_801 : _GEN_561; // @[executor.scala 470:55]
  wire [7:0] _GEN_1042 = opcode_1 != 4'h0 ? _GEN_806 : _GEN_562; // @[executor.scala 470:55]
  wire [7:0] _GEN_1043 = opcode_1 != 4'h0 ? _GEN_807 : _GEN_563; // @[executor.scala 470:55]
  wire [7:0] _GEN_1044 = opcode_1 != 4'h0 ? _GEN_808 : _GEN_564; // @[executor.scala 470:55]
  wire [7:0] _GEN_1045 = opcode_1 != 4'h0 ? _GEN_809 : _GEN_565; // @[executor.scala 470:55]
  wire [7:0] _GEN_1046 = opcode_1 != 4'h0 ? _GEN_814 : _GEN_566; // @[executor.scala 470:55]
  wire [7:0] _GEN_1047 = opcode_1 != 4'h0 ? _GEN_815 : _GEN_567; // @[executor.scala 470:55]
  wire [7:0] _GEN_1048 = opcode_1 != 4'h0 ? _GEN_816 : _GEN_568; // @[executor.scala 470:55]
  wire [7:0] _GEN_1049 = opcode_1 != 4'h0 ? _GEN_817 : _GEN_569; // @[executor.scala 470:55]
  wire [7:0] _GEN_1050 = opcode_1 != 4'h0 ? _GEN_822 : _GEN_570; // @[executor.scala 470:55]
  wire [7:0] _GEN_1051 = opcode_1 != 4'h0 ? _GEN_823 : _GEN_571; // @[executor.scala 470:55]
  wire [7:0] _GEN_1052 = opcode_1 != 4'h0 ? _GEN_824 : _GEN_572; // @[executor.scala 470:55]
  wire [7:0] _GEN_1053 = opcode_1 != 4'h0 ? _GEN_825 : _GEN_573; // @[executor.scala 470:55]
  wire [7:0] _GEN_1054 = opcode_1 != 4'h0 ? _GEN_830 : _GEN_574; // @[executor.scala 470:55]
  wire [7:0] _GEN_1055 = opcode_1 != 4'h0 ? _GEN_831 : _GEN_575; // @[executor.scala 470:55]
  wire [7:0] _GEN_1056 = opcode_1 != 4'h0 ? _GEN_832 : _GEN_576; // @[executor.scala 470:55]
  wire [7:0] _GEN_1057 = opcode_1 != 4'h0 ? _GEN_833 : _GEN_577; // @[executor.scala 470:55]
  wire [7:0] _GEN_1058 = opcode_1 != 4'h0 ? _GEN_838 : _GEN_578; // @[executor.scala 470:55]
  wire [7:0] _GEN_1059 = opcode_1 != 4'h0 ? _GEN_839 : _GEN_579; // @[executor.scala 470:55]
  wire [7:0] _GEN_1060 = opcode_1 != 4'h0 ? _GEN_840 : _GEN_580; // @[executor.scala 470:55]
  wire [7:0] _GEN_1061 = opcode_1 != 4'h0 ? _GEN_841 : _GEN_581; // @[executor.scala 470:55]
  wire [7:0] _GEN_1062 = opcode_1 != 4'h0 ? _GEN_846 : _GEN_582; // @[executor.scala 470:55]
  wire [7:0] _GEN_1063 = opcode_1 != 4'h0 ? _GEN_847 : _GEN_583; // @[executor.scala 470:55]
  wire [7:0] _GEN_1064 = opcode_1 != 4'h0 ? _GEN_848 : _GEN_584; // @[executor.scala 470:55]
  wire [7:0] _GEN_1065 = opcode_1 != 4'h0 ? _GEN_849 : _GEN_585; // @[executor.scala 470:55]
  wire [7:0] _GEN_1066 = opcode_1 != 4'h0 ? _GEN_854 : _GEN_586; // @[executor.scala 470:55]
  wire [7:0] _GEN_1067 = opcode_1 != 4'h0 ? _GEN_855 : _GEN_587; // @[executor.scala 470:55]
  wire [7:0] _GEN_1068 = opcode_1 != 4'h0 ? _GEN_856 : _GEN_588; // @[executor.scala 470:55]
  wire [7:0] _GEN_1069 = opcode_1 != 4'h0 ? _GEN_857 : _GEN_589; // @[executor.scala 470:55]
  wire [7:0] _GEN_1070 = opcode_1 != 4'h0 ? _GEN_862 : _GEN_590; // @[executor.scala 470:55]
  wire [7:0] _GEN_1071 = opcode_1 != 4'h0 ? _GEN_863 : _GEN_591; // @[executor.scala 470:55]
  wire [7:0] _GEN_1072 = opcode_1 != 4'h0 ? _GEN_864 : _GEN_592; // @[executor.scala 470:55]
  wire [7:0] _GEN_1073 = opcode_1 != 4'h0 ? _GEN_865 : _GEN_593; // @[executor.scala 470:55]
  wire [7:0] _GEN_1074 = opcode_1 != 4'h0 ? _GEN_870 : _GEN_594; // @[executor.scala 470:55]
  wire [7:0] _GEN_1075 = opcode_1 != 4'h0 ? _GEN_871 : _GEN_595; // @[executor.scala 470:55]
  wire [7:0] _GEN_1076 = opcode_1 != 4'h0 ? _GEN_872 : _GEN_596; // @[executor.scala 470:55]
  wire [7:0] _GEN_1077 = opcode_1 != 4'h0 ? _GEN_873 : _GEN_597; // @[executor.scala 470:55]
  wire [7:0] _GEN_1078 = opcode_1 != 4'h0 ? _GEN_878 : _GEN_598; // @[executor.scala 470:55]
  wire [7:0] _GEN_1079 = opcode_1 != 4'h0 ? _GEN_879 : _GEN_599; // @[executor.scala 470:55]
  wire [7:0] _GEN_1080 = opcode_1 != 4'h0 ? _GEN_880 : _GEN_600; // @[executor.scala 470:55]
  wire [7:0] _GEN_1081 = opcode_1 != 4'h0 ? _GEN_881 : _GEN_601; // @[executor.scala 470:55]
  wire [7:0] _GEN_1082 = opcode_1 != 4'h0 ? _GEN_886 : _GEN_602; // @[executor.scala 470:55]
  wire [7:0] _GEN_1083 = opcode_1 != 4'h0 ? _GEN_887 : _GEN_603; // @[executor.scala 470:55]
  wire [7:0] _GEN_1084 = opcode_1 != 4'h0 ? _GEN_888 : _GEN_604; // @[executor.scala 470:55]
  wire [7:0] _GEN_1085 = opcode_1 != 4'h0 ? _GEN_889 : _GEN_605; // @[executor.scala 470:55]
  wire [7:0] _GEN_1086 = opcode_1 != 4'h0 ? _GEN_894 : _GEN_606; // @[executor.scala 470:55]
  wire [7:0] _GEN_1087 = opcode_1 != 4'h0 ? _GEN_895 : _GEN_607; // @[executor.scala 470:55]
  wire [7:0] _GEN_1088 = opcode_1 != 4'h0 ? _GEN_896 : _GEN_608; // @[executor.scala 470:55]
  wire [7:0] _GEN_1089 = opcode_1 != 4'h0 ? _GEN_897 : _GEN_609; // @[executor.scala 470:55]
  wire [7:0] _GEN_1090 = opcode_1 != 4'h0 ? _GEN_902 : _GEN_610; // @[executor.scala 470:55]
  wire [7:0] _GEN_1091 = opcode_1 != 4'h0 ? _GEN_903 : _GEN_611; // @[executor.scala 470:55]
  wire [7:0] _GEN_1092 = opcode_1 != 4'h0 ? _GEN_904 : _GEN_612; // @[executor.scala 470:55]
  wire [7:0] _GEN_1093 = opcode_1 != 4'h0 ? _GEN_905 : _GEN_613; // @[executor.scala 470:55]
  wire [7:0] _GEN_1094 = opcode_1 != 4'h0 ? _GEN_910 : _GEN_614; // @[executor.scala 470:55]
  wire [7:0] _GEN_1095 = opcode_1 != 4'h0 ? _GEN_911 : _GEN_615; // @[executor.scala 470:55]
  wire [7:0] _GEN_1096 = opcode_1 != 4'h0 ? _GEN_912 : _GEN_616; // @[executor.scala 470:55]
  wire [7:0] _GEN_1097 = opcode_1 != 4'h0 ? _GEN_913 : _GEN_617; // @[executor.scala 470:55]
  wire [7:0] _GEN_1098 = opcode_1 != 4'h0 ? _GEN_918 : _GEN_618; // @[executor.scala 470:55]
  wire [7:0] _GEN_1099 = opcode_1 != 4'h0 ? _GEN_919 : _GEN_619; // @[executor.scala 470:55]
  wire [7:0] _GEN_1100 = opcode_1 != 4'h0 ? _GEN_920 : _GEN_620; // @[executor.scala 470:55]
  wire [7:0] _GEN_1101 = opcode_1 != 4'h0 ? _GEN_921 : _GEN_621; // @[executor.scala 470:55]
  wire [7:0] _GEN_1102 = opcode_1 != 4'h0 ? _GEN_926 : _GEN_622; // @[executor.scala 470:55]
  wire [7:0] _GEN_1103 = opcode_1 != 4'h0 ? _GEN_927 : _GEN_623; // @[executor.scala 470:55]
  wire [7:0] _GEN_1104 = opcode_1 != 4'h0 ? _GEN_928 : _GEN_624; // @[executor.scala 470:55]
  wire [7:0] _GEN_1105 = opcode_1 != 4'h0 ? _GEN_929 : _GEN_625; // @[executor.scala 470:55]
  wire [7:0] _GEN_1106 = opcode_1 != 4'h0 ? _GEN_934 : _GEN_626; // @[executor.scala 470:55]
  wire [7:0] _GEN_1107 = opcode_1 != 4'h0 ? _GEN_935 : _GEN_627; // @[executor.scala 470:55]
  wire [7:0] _GEN_1108 = opcode_1 != 4'h0 ? _GEN_936 : _GEN_628; // @[executor.scala 470:55]
  wire [7:0] _GEN_1109 = opcode_1 != 4'h0 ? _GEN_937 : _GEN_629; // @[executor.scala 470:55]
  wire [7:0] _GEN_1110 = opcode_1 != 4'h0 ? _GEN_942 : _GEN_630; // @[executor.scala 470:55]
  wire [7:0] _GEN_1111 = opcode_1 != 4'h0 ? _GEN_943 : _GEN_631; // @[executor.scala 470:55]
  wire [7:0] _GEN_1112 = opcode_1 != 4'h0 ? _GEN_944 : _GEN_632; // @[executor.scala 470:55]
  wire [7:0] _GEN_1113 = opcode_1 != 4'h0 ? _GEN_945 : _GEN_633; // @[executor.scala 470:55]
  wire [7:0] _GEN_1114 = opcode_1 != 4'h0 ? _GEN_950 : _GEN_634; // @[executor.scala 470:55]
  wire [7:0] _GEN_1115 = opcode_1 != 4'h0 ? _GEN_951 : _GEN_635; // @[executor.scala 470:55]
  wire [7:0] _GEN_1116 = opcode_1 != 4'h0 ? _GEN_952 : _GEN_636; // @[executor.scala 470:55]
  wire [7:0] _GEN_1117 = opcode_1 != 4'h0 ? _GEN_953 : _GEN_637; // @[executor.scala 470:55]
  wire [7:0] _GEN_1118 = opcode_1 != 4'h0 ? _GEN_958 : _GEN_638; // @[executor.scala 470:55]
  wire [7:0] _GEN_1119 = opcode_1 != 4'h0 ? _GEN_959 : _GEN_639; // @[executor.scala 470:55]
  wire [7:0] _GEN_1120 = opcode_1 != 4'h0 ? _GEN_960 : _GEN_640; // @[executor.scala 470:55]
  wire [7:0] _GEN_1121 = opcode_1 != 4'h0 ? _GEN_961 : _GEN_641; // @[executor.scala 470:55]
  wire [3:0] _GEN_1122 = opcode_1 == 4'hf ? parameter_2_1[13:10] : _GEN_480; // @[executor.scala 466:52 executor.scala 467:55]
  wire  _GEN_1123 = opcode_1 == 4'hf ? parameter_2_1[0] : _GEN_481; // @[executor.scala 466:52 executor.scala 468:55]
  wire [7:0] _GEN_1124 = opcode_1 == 4'hf ? _GEN_482 : _GEN_962; // @[executor.scala 466:52]
  wire [7:0] _GEN_1125 = opcode_1 == 4'hf ? _GEN_483 : _GEN_963; // @[executor.scala 466:52]
  wire [7:0] _GEN_1126 = opcode_1 == 4'hf ? _GEN_484 : _GEN_964; // @[executor.scala 466:52]
  wire [7:0] _GEN_1127 = opcode_1 == 4'hf ? _GEN_485 : _GEN_965; // @[executor.scala 466:52]
  wire [7:0] _GEN_1128 = opcode_1 == 4'hf ? _GEN_486 : _GEN_966; // @[executor.scala 466:52]
  wire [7:0] _GEN_1129 = opcode_1 == 4'hf ? _GEN_487 : _GEN_967; // @[executor.scala 466:52]
  wire [7:0] _GEN_1130 = opcode_1 == 4'hf ? _GEN_488 : _GEN_968; // @[executor.scala 466:52]
  wire [7:0] _GEN_1131 = opcode_1 == 4'hf ? _GEN_489 : _GEN_969; // @[executor.scala 466:52]
  wire [7:0] _GEN_1132 = opcode_1 == 4'hf ? _GEN_490 : _GEN_970; // @[executor.scala 466:52]
  wire [7:0] _GEN_1133 = opcode_1 == 4'hf ? _GEN_491 : _GEN_971; // @[executor.scala 466:52]
  wire [7:0] _GEN_1134 = opcode_1 == 4'hf ? _GEN_492 : _GEN_972; // @[executor.scala 466:52]
  wire [7:0] _GEN_1135 = opcode_1 == 4'hf ? _GEN_493 : _GEN_973; // @[executor.scala 466:52]
  wire [7:0] _GEN_1136 = opcode_1 == 4'hf ? _GEN_494 : _GEN_974; // @[executor.scala 466:52]
  wire [7:0] _GEN_1137 = opcode_1 == 4'hf ? _GEN_495 : _GEN_975; // @[executor.scala 466:52]
  wire [7:0] _GEN_1138 = opcode_1 == 4'hf ? _GEN_496 : _GEN_976; // @[executor.scala 466:52]
  wire [7:0] _GEN_1139 = opcode_1 == 4'hf ? _GEN_497 : _GEN_977; // @[executor.scala 466:52]
  wire [7:0] _GEN_1140 = opcode_1 == 4'hf ? _GEN_498 : _GEN_978; // @[executor.scala 466:52]
  wire [7:0] _GEN_1141 = opcode_1 == 4'hf ? _GEN_499 : _GEN_979; // @[executor.scala 466:52]
  wire [7:0] _GEN_1142 = opcode_1 == 4'hf ? _GEN_500 : _GEN_980; // @[executor.scala 466:52]
  wire [7:0] _GEN_1143 = opcode_1 == 4'hf ? _GEN_501 : _GEN_981; // @[executor.scala 466:52]
  wire [7:0] _GEN_1144 = opcode_1 == 4'hf ? _GEN_502 : _GEN_982; // @[executor.scala 466:52]
  wire [7:0] _GEN_1145 = opcode_1 == 4'hf ? _GEN_503 : _GEN_983; // @[executor.scala 466:52]
  wire [7:0] _GEN_1146 = opcode_1 == 4'hf ? _GEN_504 : _GEN_984; // @[executor.scala 466:52]
  wire [7:0] _GEN_1147 = opcode_1 == 4'hf ? _GEN_505 : _GEN_985; // @[executor.scala 466:52]
  wire [7:0] _GEN_1148 = opcode_1 == 4'hf ? _GEN_506 : _GEN_986; // @[executor.scala 466:52]
  wire [7:0] _GEN_1149 = opcode_1 == 4'hf ? _GEN_507 : _GEN_987; // @[executor.scala 466:52]
  wire [7:0] _GEN_1150 = opcode_1 == 4'hf ? _GEN_508 : _GEN_988; // @[executor.scala 466:52]
  wire [7:0] _GEN_1151 = opcode_1 == 4'hf ? _GEN_509 : _GEN_989; // @[executor.scala 466:52]
  wire [7:0] _GEN_1152 = opcode_1 == 4'hf ? _GEN_510 : _GEN_990; // @[executor.scala 466:52]
  wire [7:0] _GEN_1153 = opcode_1 == 4'hf ? _GEN_511 : _GEN_991; // @[executor.scala 466:52]
  wire [7:0] _GEN_1154 = opcode_1 == 4'hf ? _GEN_512 : _GEN_992; // @[executor.scala 466:52]
  wire [7:0] _GEN_1155 = opcode_1 == 4'hf ? _GEN_513 : _GEN_993; // @[executor.scala 466:52]
  wire [7:0] _GEN_1156 = opcode_1 == 4'hf ? _GEN_514 : _GEN_994; // @[executor.scala 466:52]
  wire [7:0] _GEN_1157 = opcode_1 == 4'hf ? _GEN_515 : _GEN_995; // @[executor.scala 466:52]
  wire [7:0] _GEN_1158 = opcode_1 == 4'hf ? _GEN_516 : _GEN_996; // @[executor.scala 466:52]
  wire [7:0] _GEN_1159 = opcode_1 == 4'hf ? _GEN_517 : _GEN_997; // @[executor.scala 466:52]
  wire [7:0] _GEN_1160 = opcode_1 == 4'hf ? _GEN_518 : _GEN_998; // @[executor.scala 466:52]
  wire [7:0] _GEN_1161 = opcode_1 == 4'hf ? _GEN_519 : _GEN_999; // @[executor.scala 466:52]
  wire [7:0] _GEN_1162 = opcode_1 == 4'hf ? _GEN_520 : _GEN_1000; // @[executor.scala 466:52]
  wire [7:0] _GEN_1163 = opcode_1 == 4'hf ? _GEN_521 : _GEN_1001; // @[executor.scala 466:52]
  wire [7:0] _GEN_1164 = opcode_1 == 4'hf ? _GEN_522 : _GEN_1002; // @[executor.scala 466:52]
  wire [7:0] _GEN_1165 = opcode_1 == 4'hf ? _GEN_523 : _GEN_1003; // @[executor.scala 466:52]
  wire [7:0] _GEN_1166 = opcode_1 == 4'hf ? _GEN_524 : _GEN_1004; // @[executor.scala 466:52]
  wire [7:0] _GEN_1167 = opcode_1 == 4'hf ? _GEN_525 : _GEN_1005; // @[executor.scala 466:52]
  wire [7:0] _GEN_1168 = opcode_1 == 4'hf ? _GEN_526 : _GEN_1006; // @[executor.scala 466:52]
  wire [7:0] _GEN_1169 = opcode_1 == 4'hf ? _GEN_527 : _GEN_1007; // @[executor.scala 466:52]
  wire [7:0] _GEN_1170 = opcode_1 == 4'hf ? _GEN_528 : _GEN_1008; // @[executor.scala 466:52]
  wire [7:0] _GEN_1171 = opcode_1 == 4'hf ? _GEN_529 : _GEN_1009; // @[executor.scala 466:52]
  wire [7:0] _GEN_1172 = opcode_1 == 4'hf ? _GEN_530 : _GEN_1010; // @[executor.scala 466:52]
  wire [7:0] _GEN_1173 = opcode_1 == 4'hf ? _GEN_531 : _GEN_1011; // @[executor.scala 466:52]
  wire [7:0] _GEN_1174 = opcode_1 == 4'hf ? _GEN_532 : _GEN_1012; // @[executor.scala 466:52]
  wire [7:0] _GEN_1175 = opcode_1 == 4'hf ? _GEN_533 : _GEN_1013; // @[executor.scala 466:52]
  wire [7:0] _GEN_1176 = opcode_1 == 4'hf ? _GEN_534 : _GEN_1014; // @[executor.scala 466:52]
  wire [7:0] _GEN_1177 = opcode_1 == 4'hf ? _GEN_535 : _GEN_1015; // @[executor.scala 466:52]
  wire [7:0] _GEN_1178 = opcode_1 == 4'hf ? _GEN_536 : _GEN_1016; // @[executor.scala 466:52]
  wire [7:0] _GEN_1179 = opcode_1 == 4'hf ? _GEN_537 : _GEN_1017; // @[executor.scala 466:52]
  wire [7:0] _GEN_1180 = opcode_1 == 4'hf ? _GEN_538 : _GEN_1018; // @[executor.scala 466:52]
  wire [7:0] _GEN_1181 = opcode_1 == 4'hf ? _GEN_539 : _GEN_1019; // @[executor.scala 466:52]
  wire [7:0] _GEN_1182 = opcode_1 == 4'hf ? _GEN_540 : _GEN_1020; // @[executor.scala 466:52]
  wire [7:0] _GEN_1183 = opcode_1 == 4'hf ? _GEN_541 : _GEN_1021; // @[executor.scala 466:52]
  wire [7:0] _GEN_1184 = opcode_1 == 4'hf ? _GEN_542 : _GEN_1022; // @[executor.scala 466:52]
  wire [7:0] _GEN_1185 = opcode_1 == 4'hf ? _GEN_543 : _GEN_1023; // @[executor.scala 466:52]
  wire [7:0] _GEN_1186 = opcode_1 == 4'hf ? _GEN_544 : _GEN_1024; // @[executor.scala 466:52]
  wire [7:0] _GEN_1187 = opcode_1 == 4'hf ? _GEN_545 : _GEN_1025; // @[executor.scala 466:52]
  wire [7:0] _GEN_1188 = opcode_1 == 4'hf ? _GEN_546 : _GEN_1026; // @[executor.scala 466:52]
  wire [7:0] _GEN_1189 = opcode_1 == 4'hf ? _GEN_547 : _GEN_1027; // @[executor.scala 466:52]
  wire [7:0] _GEN_1190 = opcode_1 == 4'hf ? _GEN_548 : _GEN_1028; // @[executor.scala 466:52]
  wire [7:0] _GEN_1191 = opcode_1 == 4'hf ? _GEN_549 : _GEN_1029; // @[executor.scala 466:52]
  wire [7:0] _GEN_1192 = opcode_1 == 4'hf ? _GEN_550 : _GEN_1030; // @[executor.scala 466:52]
  wire [7:0] _GEN_1193 = opcode_1 == 4'hf ? _GEN_551 : _GEN_1031; // @[executor.scala 466:52]
  wire [7:0] _GEN_1194 = opcode_1 == 4'hf ? _GEN_552 : _GEN_1032; // @[executor.scala 466:52]
  wire [7:0] _GEN_1195 = opcode_1 == 4'hf ? _GEN_553 : _GEN_1033; // @[executor.scala 466:52]
  wire [7:0] _GEN_1196 = opcode_1 == 4'hf ? _GEN_554 : _GEN_1034; // @[executor.scala 466:52]
  wire [7:0] _GEN_1197 = opcode_1 == 4'hf ? _GEN_555 : _GEN_1035; // @[executor.scala 466:52]
  wire [7:0] _GEN_1198 = opcode_1 == 4'hf ? _GEN_556 : _GEN_1036; // @[executor.scala 466:52]
  wire [7:0] _GEN_1199 = opcode_1 == 4'hf ? _GEN_557 : _GEN_1037; // @[executor.scala 466:52]
  wire [7:0] _GEN_1200 = opcode_1 == 4'hf ? _GEN_558 : _GEN_1038; // @[executor.scala 466:52]
  wire [7:0] _GEN_1201 = opcode_1 == 4'hf ? _GEN_559 : _GEN_1039; // @[executor.scala 466:52]
  wire [7:0] _GEN_1202 = opcode_1 == 4'hf ? _GEN_560 : _GEN_1040; // @[executor.scala 466:52]
  wire [7:0] _GEN_1203 = opcode_1 == 4'hf ? _GEN_561 : _GEN_1041; // @[executor.scala 466:52]
  wire [7:0] _GEN_1204 = opcode_1 == 4'hf ? _GEN_562 : _GEN_1042; // @[executor.scala 466:52]
  wire [7:0] _GEN_1205 = opcode_1 == 4'hf ? _GEN_563 : _GEN_1043; // @[executor.scala 466:52]
  wire [7:0] _GEN_1206 = opcode_1 == 4'hf ? _GEN_564 : _GEN_1044; // @[executor.scala 466:52]
  wire [7:0] _GEN_1207 = opcode_1 == 4'hf ? _GEN_565 : _GEN_1045; // @[executor.scala 466:52]
  wire [7:0] _GEN_1208 = opcode_1 == 4'hf ? _GEN_566 : _GEN_1046; // @[executor.scala 466:52]
  wire [7:0] _GEN_1209 = opcode_1 == 4'hf ? _GEN_567 : _GEN_1047; // @[executor.scala 466:52]
  wire [7:0] _GEN_1210 = opcode_1 == 4'hf ? _GEN_568 : _GEN_1048; // @[executor.scala 466:52]
  wire [7:0] _GEN_1211 = opcode_1 == 4'hf ? _GEN_569 : _GEN_1049; // @[executor.scala 466:52]
  wire [7:0] _GEN_1212 = opcode_1 == 4'hf ? _GEN_570 : _GEN_1050; // @[executor.scala 466:52]
  wire [7:0] _GEN_1213 = opcode_1 == 4'hf ? _GEN_571 : _GEN_1051; // @[executor.scala 466:52]
  wire [7:0] _GEN_1214 = opcode_1 == 4'hf ? _GEN_572 : _GEN_1052; // @[executor.scala 466:52]
  wire [7:0] _GEN_1215 = opcode_1 == 4'hf ? _GEN_573 : _GEN_1053; // @[executor.scala 466:52]
  wire [7:0] _GEN_1216 = opcode_1 == 4'hf ? _GEN_574 : _GEN_1054; // @[executor.scala 466:52]
  wire [7:0] _GEN_1217 = opcode_1 == 4'hf ? _GEN_575 : _GEN_1055; // @[executor.scala 466:52]
  wire [7:0] _GEN_1218 = opcode_1 == 4'hf ? _GEN_576 : _GEN_1056; // @[executor.scala 466:52]
  wire [7:0] _GEN_1219 = opcode_1 == 4'hf ? _GEN_577 : _GEN_1057; // @[executor.scala 466:52]
  wire [7:0] _GEN_1220 = opcode_1 == 4'hf ? _GEN_578 : _GEN_1058; // @[executor.scala 466:52]
  wire [7:0] _GEN_1221 = opcode_1 == 4'hf ? _GEN_579 : _GEN_1059; // @[executor.scala 466:52]
  wire [7:0] _GEN_1222 = opcode_1 == 4'hf ? _GEN_580 : _GEN_1060; // @[executor.scala 466:52]
  wire [7:0] _GEN_1223 = opcode_1 == 4'hf ? _GEN_581 : _GEN_1061; // @[executor.scala 466:52]
  wire [7:0] _GEN_1224 = opcode_1 == 4'hf ? _GEN_582 : _GEN_1062; // @[executor.scala 466:52]
  wire [7:0] _GEN_1225 = opcode_1 == 4'hf ? _GEN_583 : _GEN_1063; // @[executor.scala 466:52]
  wire [7:0] _GEN_1226 = opcode_1 == 4'hf ? _GEN_584 : _GEN_1064; // @[executor.scala 466:52]
  wire [7:0] _GEN_1227 = opcode_1 == 4'hf ? _GEN_585 : _GEN_1065; // @[executor.scala 466:52]
  wire [7:0] _GEN_1228 = opcode_1 == 4'hf ? _GEN_586 : _GEN_1066; // @[executor.scala 466:52]
  wire [7:0] _GEN_1229 = opcode_1 == 4'hf ? _GEN_587 : _GEN_1067; // @[executor.scala 466:52]
  wire [7:0] _GEN_1230 = opcode_1 == 4'hf ? _GEN_588 : _GEN_1068; // @[executor.scala 466:52]
  wire [7:0] _GEN_1231 = opcode_1 == 4'hf ? _GEN_589 : _GEN_1069; // @[executor.scala 466:52]
  wire [7:0] _GEN_1232 = opcode_1 == 4'hf ? _GEN_590 : _GEN_1070; // @[executor.scala 466:52]
  wire [7:0] _GEN_1233 = opcode_1 == 4'hf ? _GEN_591 : _GEN_1071; // @[executor.scala 466:52]
  wire [7:0] _GEN_1234 = opcode_1 == 4'hf ? _GEN_592 : _GEN_1072; // @[executor.scala 466:52]
  wire [7:0] _GEN_1235 = opcode_1 == 4'hf ? _GEN_593 : _GEN_1073; // @[executor.scala 466:52]
  wire [7:0] _GEN_1236 = opcode_1 == 4'hf ? _GEN_594 : _GEN_1074; // @[executor.scala 466:52]
  wire [7:0] _GEN_1237 = opcode_1 == 4'hf ? _GEN_595 : _GEN_1075; // @[executor.scala 466:52]
  wire [7:0] _GEN_1238 = opcode_1 == 4'hf ? _GEN_596 : _GEN_1076; // @[executor.scala 466:52]
  wire [7:0] _GEN_1239 = opcode_1 == 4'hf ? _GEN_597 : _GEN_1077; // @[executor.scala 466:52]
  wire [7:0] _GEN_1240 = opcode_1 == 4'hf ? _GEN_598 : _GEN_1078; // @[executor.scala 466:52]
  wire [7:0] _GEN_1241 = opcode_1 == 4'hf ? _GEN_599 : _GEN_1079; // @[executor.scala 466:52]
  wire [7:0] _GEN_1242 = opcode_1 == 4'hf ? _GEN_600 : _GEN_1080; // @[executor.scala 466:52]
  wire [7:0] _GEN_1243 = opcode_1 == 4'hf ? _GEN_601 : _GEN_1081; // @[executor.scala 466:52]
  wire [7:0] _GEN_1244 = opcode_1 == 4'hf ? _GEN_602 : _GEN_1082; // @[executor.scala 466:52]
  wire [7:0] _GEN_1245 = opcode_1 == 4'hf ? _GEN_603 : _GEN_1083; // @[executor.scala 466:52]
  wire [7:0] _GEN_1246 = opcode_1 == 4'hf ? _GEN_604 : _GEN_1084; // @[executor.scala 466:52]
  wire [7:0] _GEN_1247 = opcode_1 == 4'hf ? _GEN_605 : _GEN_1085; // @[executor.scala 466:52]
  wire [7:0] _GEN_1248 = opcode_1 == 4'hf ? _GEN_606 : _GEN_1086; // @[executor.scala 466:52]
  wire [7:0] _GEN_1249 = opcode_1 == 4'hf ? _GEN_607 : _GEN_1087; // @[executor.scala 466:52]
  wire [7:0] _GEN_1250 = opcode_1 == 4'hf ? _GEN_608 : _GEN_1088; // @[executor.scala 466:52]
  wire [7:0] _GEN_1251 = opcode_1 == 4'hf ? _GEN_609 : _GEN_1089; // @[executor.scala 466:52]
  wire [7:0] _GEN_1252 = opcode_1 == 4'hf ? _GEN_610 : _GEN_1090; // @[executor.scala 466:52]
  wire [7:0] _GEN_1253 = opcode_1 == 4'hf ? _GEN_611 : _GEN_1091; // @[executor.scala 466:52]
  wire [7:0] _GEN_1254 = opcode_1 == 4'hf ? _GEN_612 : _GEN_1092; // @[executor.scala 466:52]
  wire [7:0] _GEN_1255 = opcode_1 == 4'hf ? _GEN_613 : _GEN_1093; // @[executor.scala 466:52]
  wire [7:0] _GEN_1256 = opcode_1 == 4'hf ? _GEN_614 : _GEN_1094; // @[executor.scala 466:52]
  wire [7:0] _GEN_1257 = opcode_1 == 4'hf ? _GEN_615 : _GEN_1095; // @[executor.scala 466:52]
  wire [7:0] _GEN_1258 = opcode_1 == 4'hf ? _GEN_616 : _GEN_1096; // @[executor.scala 466:52]
  wire [7:0] _GEN_1259 = opcode_1 == 4'hf ? _GEN_617 : _GEN_1097; // @[executor.scala 466:52]
  wire [7:0] _GEN_1260 = opcode_1 == 4'hf ? _GEN_618 : _GEN_1098; // @[executor.scala 466:52]
  wire [7:0] _GEN_1261 = opcode_1 == 4'hf ? _GEN_619 : _GEN_1099; // @[executor.scala 466:52]
  wire [7:0] _GEN_1262 = opcode_1 == 4'hf ? _GEN_620 : _GEN_1100; // @[executor.scala 466:52]
  wire [7:0] _GEN_1263 = opcode_1 == 4'hf ? _GEN_621 : _GEN_1101; // @[executor.scala 466:52]
  wire [7:0] _GEN_1264 = opcode_1 == 4'hf ? _GEN_622 : _GEN_1102; // @[executor.scala 466:52]
  wire [7:0] _GEN_1265 = opcode_1 == 4'hf ? _GEN_623 : _GEN_1103; // @[executor.scala 466:52]
  wire [7:0] _GEN_1266 = opcode_1 == 4'hf ? _GEN_624 : _GEN_1104; // @[executor.scala 466:52]
  wire [7:0] _GEN_1267 = opcode_1 == 4'hf ? _GEN_625 : _GEN_1105; // @[executor.scala 466:52]
  wire [7:0] _GEN_1268 = opcode_1 == 4'hf ? _GEN_626 : _GEN_1106; // @[executor.scala 466:52]
  wire [7:0] _GEN_1269 = opcode_1 == 4'hf ? _GEN_627 : _GEN_1107; // @[executor.scala 466:52]
  wire [7:0] _GEN_1270 = opcode_1 == 4'hf ? _GEN_628 : _GEN_1108; // @[executor.scala 466:52]
  wire [7:0] _GEN_1271 = opcode_1 == 4'hf ? _GEN_629 : _GEN_1109; // @[executor.scala 466:52]
  wire [7:0] _GEN_1272 = opcode_1 == 4'hf ? _GEN_630 : _GEN_1110; // @[executor.scala 466:52]
  wire [7:0] _GEN_1273 = opcode_1 == 4'hf ? _GEN_631 : _GEN_1111; // @[executor.scala 466:52]
  wire [7:0] _GEN_1274 = opcode_1 == 4'hf ? _GEN_632 : _GEN_1112; // @[executor.scala 466:52]
  wire [7:0] _GEN_1275 = opcode_1 == 4'hf ? _GEN_633 : _GEN_1113; // @[executor.scala 466:52]
  wire [7:0] _GEN_1276 = opcode_1 == 4'hf ? _GEN_634 : _GEN_1114; // @[executor.scala 466:52]
  wire [7:0] _GEN_1277 = opcode_1 == 4'hf ? _GEN_635 : _GEN_1115; // @[executor.scala 466:52]
  wire [7:0] _GEN_1278 = opcode_1 == 4'hf ? _GEN_636 : _GEN_1116; // @[executor.scala 466:52]
  wire [7:0] _GEN_1279 = opcode_1 == 4'hf ? _GEN_637 : _GEN_1117; // @[executor.scala 466:52]
  wire [7:0] _GEN_1280 = opcode_1 == 4'hf ? _GEN_638 : _GEN_1118; // @[executor.scala 466:52]
  wire [7:0] _GEN_1281 = opcode_1 == 4'hf ? _GEN_639 : _GEN_1119; // @[executor.scala 466:52]
  wire [7:0] _GEN_1282 = opcode_1 == 4'hf ? _GEN_640 : _GEN_1120; // @[executor.scala 466:52]
  wire [7:0] _GEN_1283 = opcode_1 == 4'hf ? _GEN_641 : _GEN_1121; // @[executor.scala 466:52]
  wire [3:0] opcode_2 = vliw_2[31:28]; // @[primitive.scala 9:44]
  wire [13:0] parameter_2_2 = vliw_2[13:0]; // @[primitive.scala 11:44]
  wire [7:0] _GEN_2810 = {{2'd0}, dst_offset_2}; // @[executor.scala 473:49]
  wire [7:0] byte_320 = field_2[7:0]; // @[executor.scala 475:56]
  wire [7:0] _GEN_1284 = mask_2[0] ? byte_320 : _GEN_1124; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] byte_321 = field_2[15:8]; // @[executor.scala 475:56]
  wire [7:0] _GEN_1285 = mask_2[1] ? byte_321 : _GEN_1125; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] byte_322 = field_2[23:16]; // @[executor.scala 475:56]
  wire [7:0] _GEN_1286 = mask_2[2] ? byte_322 : _GEN_1126; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] byte_323 = field_2[31:24]; // @[executor.scala 475:56]
  wire [7:0] _GEN_1287 = mask_2[3] ? byte_323 : _GEN_1127; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1288 = _GEN_2810 == 8'h0 ? _GEN_1284 : _GEN_1124; // @[executor.scala 473:84]
  wire [7:0] _GEN_1289 = _GEN_2810 == 8'h0 ? _GEN_1285 : _GEN_1125; // @[executor.scala 473:84]
  wire [7:0] _GEN_1290 = _GEN_2810 == 8'h0 ? _GEN_1286 : _GEN_1126; // @[executor.scala 473:84]
  wire [7:0] _GEN_1291 = _GEN_2810 == 8'h0 ? _GEN_1287 : _GEN_1127; // @[executor.scala 473:84]
  wire [7:0] _GEN_1292 = mask_2[0] ? byte_320 : _GEN_1128; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1293 = mask_2[1] ? byte_321 : _GEN_1129; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1294 = mask_2[2] ? byte_322 : _GEN_1130; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1295 = mask_2[3] ? byte_323 : _GEN_1131; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1296 = _GEN_2810 == 8'h1 ? _GEN_1292 : _GEN_1128; // @[executor.scala 473:84]
  wire [7:0] _GEN_1297 = _GEN_2810 == 8'h1 ? _GEN_1293 : _GEN_1129; // @[executor.scala 473:84]
  wire [7:0] _GEN_1298 = _GEN_2810 == 8'h1 ? _GEN_1294 : _GEN_1130; // @[executor.scala 473:84]
  wire [7:0] _GEN_1299 = _GEN_2810 == 8'h1 ? _GEN_1295 : _GEN_1131; // @[executor.scala 473:84]
  wire [7:0] _GEN_1300 = mask_2[0] ? byte_320 : _GEN_1132; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1301 = mask_2[1] ? byte_321 : _GEN_1133; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1302 = mask_2[2] ? byte_322 : _GEN_1134; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1303 = mask_2[3] ? byte_323 : _GEN_1135; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1304 = _GEN_2810 == 8'h2 ? _GEN_1300 : _GEN_1132; // @[executor.scala 473:84]
  wire [7:0] _GEN_1305 = _GEN_2810 == 8'h2 ? _GEN_1301 : _GEN_1133; // @[executor.scala 473:84]
  wire [7:0] _GEN_1306 = _GEN_2810 == 8'h2 ? _GEN_1302 : _GEN_1134; // @[executor.scala 473:84]
  wire [7:0] _GEN_1307 = _GEN_2810 == 8'h2 ? _GEN_1303 : _GEN_1135; // @[executor.scala 473:84]
  wire [7:0] _GEN_1308 = mask_2[0] ? byte_320 : _GEN_1136; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1309 = mask_2[1] ? byte_321 : _GEN_1137; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1310 = mask_2[2] ? byte_322 : _GEN_1138; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1311 = mask_2[3] ? byte_323 : _GEN_1139; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1312 = _GEN_2810 == 8'h3 ? _GEN_1308 : _GEN_1136; // @[executor.scala 473:84]
  wire [7:0] _GEN_1313 = _GEN_2810 == 8'h3 ? _GEN_1309 : _GEN_1137; // @[executor.scala 473:84]
  wire [7:0] _GEN_1314 = _GEN_2810 == 8'h3 ? _GEN_1310 : _GEN_1138; // @[executor.scala 473:84]
  wire [7:0] _GEN_1315 = _GEN_2810 == 8'h3 ? _GEN_1311 : _GEN_1139; // @[executor.scala 473:84]
  wire [7:0] _GEN_1316 = mask_2[0] ? byte_320 : _GEN_1140; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1317 = mask_2[1] ? byte_321 : _GEN_1141; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1318 = mask_2[2] ? byte_322 : _GEN_1142; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1319 = mask_2[3] ? byte_323 : _GEN_1143; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1320 = _GEN_2810 == 8'h4 ? _GEN_1316 : _GEN_1140; // @[executor.scala 473:84]
  wire [7:0] _GEN_1321 = _GEN_2810 == 8'h4 ? _GEN_1317 : _GEN_1141; // @[executor.scala 473:84]
  wire [7:0] _GEN_1322 = _GEN_2810 == 8'h4 ? _GEN_1318 : _GEN_1142; // @[executor.scala 473:84]
  wire [7:0] _GEN_1323 = _GEN_2810 == 8'h4 ? _GEN_1319 : _GEN_1143; // @[executor.scala 473:84]
  wire [7:0] _GEN_1324 = mask_2[0] ? byte_320 : _GEN_1144; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1325 = mask_2[1] ? byte_321 : _GEN_1145; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1326 = mask_2[2] ? byte_322 : _GEN_1146; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1327 = mask_2[3] ? byte_323 : _GEN_1147; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1328 = _GEN_2810 == 8'h5 ? _GEN_1324 : _GEN_1144; // @[executor.scala 473:84]
  wire [7:0] _GEN_1329 = _GEN_2810 == 8'h5 ? _GEN_1325 : _GEN_1145; // @[executor.scala 473:84]
  wire [7:0] _GEN_1330 = _GEN_2810 == 8'h5 ? _GEN_1326 : _GEN_1146; // @[executor.scala 473:84]
  wire [7:0] _GEN_1331 = _GEN_2810 == 8'h5 ? _GEN_1327 : _GEN_1147; // @[executor.scala 473:84]
  wire [7:0] _GEN_1332 = mask_2[0] ? byte_320 : _GEN_1148; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1333 = mask_2[1] ? byte_321 : _GEN_1149; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1334 = mask_2[2] ? byte_322 : _GEN_1150; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1335 = mask_2[3] ? byte_323 : _GEN_1151; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1336 = _GEN_2810 == 8'h6 ? _GEN_1332 : _GEN_1148; // @[executor.scala 473:84]
  wire [7:0] _GEN_1337 = _GEN_2810 == 8'h6 ? _GEN_1333 : _GEN_1149; // @[executor.scala 473:84]
  wire [7:0] _GEN_1338 = _GEN_2810 == 8'h6 ? _GEN_1334 : _GEN_1150; // @[executor.scala 473:84]
  wire [7:0] _GEN_1339 = _GEN_2810 == 8'h6 ? _GEN_1335 : _GEN_1151; // @[executor.scala 473:84]
  wire [7:0] _GEN_1340 = mask_2[0] ? byte_320 : _GEN_1152; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1341 = mask_2[1] ? byte_321 : _GEN_1153; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1342 = mask_2[2] ? byte_322 : _GEN_1154; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1343 = mask_2[3] ? byte_323 : _GEN_1155; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1344 = _GEN_2810 == 8'h7 ? _GEN_1340 : _GEN_1152; // @[executor.scala 473:84]
  wire [7:0] _GEN_1345 = _GEN_2810 == 8'h7 ? _GEN_1341 : _GEN_1153; // @[executor.scala 473:84]
  wire [7:0] _GEN_1346 = _GEN_2810 == 8'h7 ? _GEN_1342 : _GEN_1154; // @[executor.scala 473:84]
  wire [7:0] _GEN_1347 = _GEN_2810 == 8'h7 ? _GEN_1343 : _GEN_1155; // @[executor.scala 473:84]
  wire [7:0] _GEN_1348 = mask_2[0] ? byte_320 : _GEN_1156; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1349 = mask_2[1] ? byte_321 : _GEN_1157; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1350 = mask_2[2] ? byte_322 : _GEN_1158; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1351 = mask_2[3] ? byte_323 : _GEN_1159; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1352 = _GEN_2810 == 8'h8 ? _GEN_1348 : _GEN_1156; // @[executor.scala 473:84]
  wire [7:0] _GEN_1353 = _GEN_2810 == 8'h8 ? _GEN_1349 : _GEN_1157; // @[executor.scala 473:84]
  wire [7:0] _GEN_1354 = _GEN_2810 == 8'h8 ? _GEN_1350 : _GEN_1158; // @[executor.scala 473:84]
  wire [7:0] _GEN_1355 = _GEN_2810 == 8'h8 ? _GEN_1351 : _GEN_1159; // @[executor.scala 473:84]
  wire [7:0] _GEN_1356 = mask_2[0] ? byte_320 : _GEN_1160; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1357 = mask_2[1] ? byte_321 : _GEN_1161; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1358 = mask_2[2] ? byte_322 : _GEN_1162; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1359 = mask_2[3] ? byte_323 : _GEN_1163; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1360 = _GEN_2810 == 8'h9 ? _GEN_1356 : _GEN_1160; // @[executor.scala 473:84]
  wire [7:0] _GEN_1361 = _GEN_2810 == 8'h9 ? _GEN_1357 : _GEN_1161; // @[executor.scala 473:84]
  wire [7:0] _GEN_1362 = _GEN_2810 == 8'h9 ? _GEN_1358 : _GEN_1162; // @[executor.scala 473:84]
  wire [7:0] _GEN_1363 = _GEN_2810 == 8'h9 ? _GEN_1359 : _GEN_1163; // @[executor.scala 473:84]
  wire [7:0] _GEN_1364 = mask_2[0] ? byte_320 : _GEN_1164; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1365 = mask_2[1] ? byte_321 : _GEN_1165; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1366 = mask_2[2] ? byte_322 : _GEN_1166; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1367 = mask_2[3] ? byte_323 : _GEN_1167; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1368 = _GEN_2810 == 8'ha ? _GEN_1364 : _GEN_1164; // @[executor.scala 473:84]
  wire [7:0] _GEN_1369 = _GEN_2810 == 8'ha ? _GEN_1365 : _GEN_1165; // @[executor.scala 473:84]
  wire [7:0] _GEN_1370 = _GEN_2810 == 8'ha ? _GEN_1366 : _GEN_1166; // @[executor.scala 473:84]
  wire [7:0] _GEN_1371 = _GEN_2810 == 8'ha ? _GEN_1367 : _GEN_1167; // @[executor.scala 473:84]
  wire [7:0] _GEN_1372 = mask_2[0] ? byte_320 : _GEN_1168; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1373 = mask_2[1] ? byte_321 : _GEN_1169; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1374 = mask_2[2] ? byte_322 : _GEN_1170; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1375 = mask_2[3] ? byte_323 : _GEN_1171; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1376 = _GEN_2810 == 8'hb ? _GEN_1372 : _GEN_1168; // @[executor.scala 473:84]
  wire [7:0] _GEN_1377 = _GEN_2810 == 8'hb ? _GEN_1373 : _GEN_1169; // @[executor.scala 473:84]
  wire [7:0] _GEN_1378 = _GEN_2810 == 8'hb ? _GEN_1374 : _GEN_1170; // @[executor.scala 473:84]
  wire [7:0] _GEN_1379 = _GEN_2810 == 8'hb ? _GEN_1375 : _GEN_1171; // @[executor.scala 473:84]
  wire [7:0] _GEN_1380 = mask_2[0] ? byte_320 : _GEN_1172; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1381 = mask_2[1] ? byte_321 : _GEN_1173; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1382 = mask_2[2] ? byte_322 : _GEN_1174; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1383 = mask_2[3] ? byte_323 : _GEN_1175; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1384 = _GEN_2810 == 8'hc ? _GEN_1380 : _GEN_1172; // @[executor.scala 473:84]
  wire [7:0] _GEN_1385 = _GEN_2810 == 8'hc ? _GEN_1381 : _GEN_1173; // @[executor.scala 473:84]
  wire [7:0] _GEN_1386 = _GEN_2810 == 8'hc ? _GEN_1382 : _GEN_1174; // @[executor.scala 473:84]
  wire [7:0] _GEN_1387 = _GEN_2810 == 8'hc ? _GEN_1383 : _GEN_1175; // @[executor.scala 473:84]
  wire [7:0] _GEN_1388 = mask_2[0] ? byte_320 : _GEN_1176; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1389 = mask_2[1] ? byte_321 : _GEN_1177; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1390 = mask_2[2] ? byte_322 : _GEN_1178; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1391 = mask_2[3] ? byte_323 : _GEN_1179; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1392 = _GEN_2810 == 8'hd ? _GEN_1388 : _GEN_1176; // @[executor.scala 473:84]
  wire [7:0] _GEN_1393 = _GEN_2810 == 8'hd ? _GEN_1389 : _GEN_1177; // @[executor.scala 473:84]
  wire [7:0] _GEN_1394 = _GEN_2810 == 8'hd ? _GEN_1390 : _GEN_1178; // @[executor.scala 473:84]
  wire [7:0] _GEN_1395 = _GEN_2810 == 8'hd ? _GEN_1391 : _GEN_1179; // @[executor.scala 473:84]
  wire [7:0] _GEN_1396 = mask_2[0] ? byte_320 : _GEN_1180; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1397 = mask_2[1] ? byte_321 : _GEN_1181; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1398 = mask_2[2] ? byte_322 : _GEN_1182; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1399 = mask_2[3] ? byte_323 : _GEN_1183; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1400 = _GEN_2810 == 8'he ? _GEN_1396 : _GEN_1180; // @[executor.scala 473:84]
  wire [7:0] _GEN_1401 = _GEN_2810 == 8'he ? _GEN_1397 : _GEN_1181; // @[executor.scala 473:84]
  wire [7:0] _GEN_1402 = _GEN_2810 == 8'he ? _GEN_1398 : _GEN_1182; // @[executor.scala 473:84]
  wire [7:0] _GEN_1403 = _GEN_2810 == 8'he ? _GEN_1399 : _GEN_1183; // @[executor.scala 473:84]
  wire [7:0] _GEN_1404 = mask_2[0] ? byte_320 : _GEN_1184; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1405 = mask_2[1] ? byte_321 : _GEN_1185; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1406 = mask_2[2] ? byte_322 : _GEN_1186; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1407 = mask_2[3] ? byte_323 : _GEN_1187; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1408 = _GEN_2810 == 8'hf ? _GEN_1404 : _GEN_1184; // @[executor.scala 473:84]
  wire [7:0] _GEN_1409 = _GEN_2810 == 8'hf ? _GEN_1405 : _GEN_1185; // @[executor.scala 473:84]
  wire [7:0] _GEN_1410 = _GEN_2810 == 8'hf ? _GEN_1406 : _GEN_1186; // @[executor.scala 473:84]
  wire [7:0] _GEN_1411 = _GEN_2810 == 8'hf ? _GEN_1407 : _GEN_1187; // @[executor.scala 473:84]
  wire [7:0] _GEN_1412 = mask_2[0] ? byte_320 : _GEN_1188; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1413 = mask_2[1] ? byte_321 : _GEN_1189; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1414 = mask_2[2] ? byte_322 : _GEN_1190; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1415 = mask_2[3] ? byte_323 : _GEN_1191; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1416 = _GEN_2810 == 8'h10 ? _GEN_1412 : _GEN_1188; // @[executor.scala 473:84]
  wire [7:0] _GEN_1417 = _GEN_2810 == 8'h10 ? _GEN_1413 : _GEN_1189; // @[executor.scala 473:84]
  wire [7:0] _GEN_1418 = _GEN_2810 == 8'h10 ? _GEN_1414 : _GEN_1190; // @[executor.scala 473:84]
  wire [7:0] _GEN_1419 = _GEN_2810 == 8'h10 ? _GEN_1415 : _GEN_1191; // @[executor.scala 473:84]
  wire [7:0] _GEN_1420 = mask_2[0] ? byte_320 : _GEN_1192; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1421 = mask_2[1] ? byte_321 : _GEN_1193; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1422 = mask_2[2] ? byte_322 : _GEN_1194; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1423 = mask_2[3] ? byte_323 : _GEN_1195; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1424 = _GEN_2810 == 8'h11 ? _GEN_1420 : _GEN_1192; // @[executor.scala 473:84]
  wire [7:0] _GEN_1425 = _GEN_2810 == 8'h11 ? _GEN_1421 : _GEN_1193; // @[executor.scala 473:84]
  wire [7:0] _GEN_1426 = _GEN_2810 == 8'h11 ? _GEN_1422 : _GEN_1194; // @[executor.scala 473:84]
  wire [7:0] _GEN_1427 = _GEN_2810 == 8'h11 ? _GEN_1423 : _GEN_1195; // @[executor.scala 473:84]
  wire [7:0] _GEN_1428 = mask_2[0] ? byte_320 : _GEN_1196; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1429 = mask_2[1] ? byte_321 : _GEN_1197; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1430 = mask_2[2] ? byte_322 : _GEN_1198; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1431 = mask_2[3] ? byte_323 : _GEN_1199; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1432 = _GEN_2810 == 8'h12 ? _GEN_1428 : _GEN_1196; // @[executor.scala 473:84]
  wire [7:0] _GEN_1433 = _GEN_2810 == 8'h12 ? _GEN_1429 : _GEN_1197; // @[executor.scala 473:84]
  wire [7:0] _GEN_1434 = _GEN_2810 == 8'h12 ? _GEN_1430 : _GEN_1198; // @[executor.scala 473:84]
  wire [7:0] _GEN_1435 = _GEN_2810 == 8'h12 ? _GEN_1431 : _GEN_1199; // @[executor.scala 473:84]
  wire [7:0] _GEN_1436 = mask_2[0] ? byte_320 : _GEN_1200; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1437 = mask_2[1] ? byte_321 : _GEN_1201; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1438 = mask_2[2] ? byte_322 : _GEN_1202; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1439 = mask_2[3] ? byte_323 : _GEN_1203; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1440 = _GEN_2810 == 8'h13 ? _GEN_1436 : _GEN_1200; // @[executor.scala 473:84]
  wire [7:0] _GEN_1441 = _GEN_2810 == 8'h13 ? _GEN_1437 : _GEN_1201; // @[executor.scala 473:84]
  wire [7:0] _GEN_1442 = _GEN_2810 == 8'h13 ? _GEN_1438 : _GEN_1202; // @[executor.scala 473:84]
  wire [7:0] _GEN_1443 = _GEN_2810 == 8'h13 ? _GEN_1439 : _GEN_1203; // @[executor.scala 473:84]
  wire [7:0] _GEN_1444 = mask_2[0] ? byte_320 : _GEN_1204; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1445 = mask_2[1] ? byte_321 : _GEN_1205; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1446 = mask_2[2] ? byte_322 : _GEN_1206; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1447 = mask_2[3] ? byte_323 : _GEN_1207; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1448 = _GEN_2810 == 8'h14 ? _GEN_1444 : _GEN_1204; // @[executor.scala 473:84]
  wire [7:0] _GEN_1449 = _GEN_2810 == 8'h14 ? _GEN_1445 : _GEN_1205; // @[executor.scala 473:84]
  wire [7:0] _GEN_1450 = _GEN_2810 == 8'h14 ? _GEN_1446 : _GEN_1206; // @[executor.scala 473:84]
  wire [7:0] _GEN_1451 = _GEN_2810 == 8'h14 ? _GEN_1447 : _GEN_1207; // @[executor.scala 473:84]
  wire [7:0] _GEN_1452 = mask_2[0] ? byte_320 : _GEN_1208; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1453 = mask_2[1] ? byte_321 : _GEN_1209; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1454 = mask_2[2] ? byte_322 : _GEN_1210; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1455 = mask_2[3] ? byte_323 : _GEN_1211; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1456 = _GEN_2810 == 8'h15 ? _GEN_1452 : _GEN_1208; // @[executor.scala 473:84]
  wire [7:0] _GEN_1457 = _GEN_2810 == 8'h15 ? _GEN_1453 : _GEN_1209; // @[executor.scala 473:84]
  wire [7:0] _GEN_1458 = _GEN_2810 == 8'h15 ? _GEN_1454 : _GEN_1210; // @[executor.scala 473:84]
  wire [7:0] _GEN_1459 = _GEN_2810 == 8'h15 ? _GEN_1455 : _GEN_1211; // @[executor.scala 473:84]
  wire [7:0] _GEN_1460 = mask_2[0] ? byte_320 : _GEN_1212; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1461 = mask_2[1] ? byte_321 : _GEN_1213; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1462 = mask_2[2] ? byte_322 : _GEN_1214; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1463 = mask_2[3] ? byte_323 : _GEN_1215; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1464 = _GEN_2810 == 8'h16 ? _GEN_1460 : _GEN_1212; // @[executor.scala 473:84]
  wire [7:0] _GEN_1465 = _GEN_2810 == 8'h16 ? _GEN_1461 : _GEN_1213; // @[executor.scala 473:84]
  wire [7:0] _GEN_1466 = _GEN_2810 == 8'h16 ? _GEN_1462 : _GEN_1214; // @[executor.scala 473:84]
  wire [7:0] _GEN_1467 = _GEN_2810 == 8'h16 ? _GEN_1463 : _GEN_1215; // @[executor.scala 473:84]
  wire [7:0] _GEN_1468 = mask_2[0] ? byte_320 : _GEN_1216; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1469 = mask_2[1] ? byte_321 : _GEN_1217; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1470 = mask_2[2] ? byte_322 : _GEN_1218; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1471 = mask_2[3] ? byte_323 : _GEN_1219; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1472 = _GEN_2810 == 8'h17 ? _GEN_1468 : _GEN_1216; // @[executor.scala 473:84]
  wire [7:0] _GEN_1473 = _GEN_2810 == 8'h17 ? _GEN_1469 : _GEN_1217; // @[executor.scala 473:84]
  wire [7:0] _GEN_1474 = _GEN_2810 == 8'h17 ? _GEN_1470 : _GEN_1218; // @[executor.scala 473:84]
  wire [7:0] _GEN_1475 = _GEN_2810 == 8'h17 ? _GEN_1471 : _GEN_1219; // @[executor.scala 473:84]
  wire [7:0] _GEN_1476 = mask_2[0] ? byte_320 : _GEN_1220; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1477 = mask_2[1] ? byte_321 : _GEN_1221; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1478 = mask_2[2] ? byte_322 : _GEN_1222; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1479 = mask_2[3] ? byte_323 : _GEN_1223; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1480 = _GEN_2810 == 8'h18 ? _GEN_1476 : _GEN_1220; // @[executor.scala 473:84]
  wire [7:0] _GEN_1481 = _GEN_2810 == 8'h18 ? _GEN_1477 : _GEN_1221; // @[executor.scala 473:84]
  wire [7:0] _GEN_1482 = _GEN_2810 == 8'h18 ? _GEN_1478 : _GEN_1222; // @[executor.scala 473:84]
  wire [7:0] _GEN_1483 = _GEN_2810 == 8'h18 ? _GEN_1479 : _GEN_1223; // @[executor.scala 473:84]
  wire [7:0] _GEN_1484 = mask_2[0] ? byte_320 : _GEN_1224; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1485 = mask_2[1] ? byte_321 : _GEN_1225; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1486 = mask_2[2] ? byte_322 : _GEN_1226; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1487 = mask_2[3] ? byte_323 : _GEN_1227; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1488 = _GEN_2810 == 8'h19 ? _GEN_1484 : _GEN_1224; // @[executor.scala 473:84]
  wire [7:0] _GEN_1489 = _GEN_2810 == 8'h19 ? _GEN_1485 : _GEN_1225; // @[executor.scala 473:84]
  wire [7:0] _GEN_1490 = _GEN_2810 == 8'h19 ? _GEN_1486 : _GEN_1226; // @[executor.scala 473:84]
  wire [7:0] _GEN_1491 = _GEN_2810 == 8'h19 ? _GEN_1487 : _GEN_1227; // @[executor.scala 473:84]
  wire [7:0] _GEN_1492 = mask_2[0] ? byte_320 : _GEN_1228; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1493 = mask_2[1] ? byte_321 : _GEN_1229; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1494 = mask_2[2] ? byte_322 : _GEN_1230; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1495 = mask_2[3] ? byte_323 : _GEN_1231; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1496 = _GEN_2810 == 8'h1a ? _GEN_1492 : _GEN_1228; // @[executor.scala 473:84]
  wire [7:0] _GEN_1497 = _GEN_2810 == 8'h1a ? _GEN_1493 : _GEN_1229; // @[executor.scala 473:84]
  wire [7:0] _GEN_1498 = _GEN_2810 == 8'h1a ? _GEN_1494 : _GEN_1230; // @[executor.scala 473:84]
  wire [7:0] _GEN_1499 = _GEN_2810 == 8'h1a ? _GEN_1495 : _GEN_1231; // @[executor.scala 473:84]
  wire [7:0] _GEN_1500 = mask_2[0] ? byte_320 : _GEN_1232; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1501 = mask_2[1] ? byte_321 : _GEN_1233; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1502 = mask_2[2] ? byte_322 : _GEN_1234; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1503 = mask_2[3] ? byte_323 : _GEN_1235; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1504 = _GEN_2810 == 8'h1b ? _GEN_1500 : _GEN_1232; // @[executor.scala 473:84]
  wire [7:0] _GEN_1505 = _GEN_2810 == 8'h1b ? _GEN_1501 : _GEN_1233; // @[executor.scala 473:84]
  wire [7:0] _GEN_1506 = _GEN_2810 == 8'h1b ? _GEN_1502 : _GEN_1234; // @[executor.scala 473:84]
  wire [7:0] _GEN_1507 = _GEN_2810 == 8'h1b ? _GEN_1503 : _GEN_1235; // @[executor.scala 473:84]
  wire [7:0] _GEN_1508 = mask_2[0] ? byte_320 : _GEN_1236; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1509 = mask_2[1] ? byte_321 : _GEN_1237; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1510 = mask_2[2] ? byte_322 : _GEN_1238; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1511 = mask_2[3] ? byte_323 : _GEN_1239; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1512 = _GEN_2810 == 8'h1c ? _GEN_1508 : _GEN_1236; // @[executor.scala 473:84]
  wire [7:0] _GEN_1513 = _GEN_2810 == 8'h1c ? _GEN_1509 : _GEN_1237; // @[executor.scala 473:84]
  wire [7:0] _GEN_1514 = _GEN_2810 == 8'h1c ? _GEN_1510 : _GEN_1238; // @[executor.scala 473:84]
  wire [7:0] _GEN_1515 = _GEN_2810 == 8'h1c ? _GEN_1511 : _GEN_1239; // @[executor.scala 473:84]
  wire [7:0] _GEN_1516 = mask_2[0] ? byte_320 : _GEN_1240; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1517 = mask_2[1] ? byte_321 : _GEN_1241; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1518 = mask_2[2] ? byte_322 : _GEN_1242; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1519 = mask_2[3] ? byte_323 : _GEN_1243; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1520 = _GEN_2810 == 8'h1d ? _GEN_1516 : _GEN_1240; // @[executor.scala 473:84]
  wire [7:0] _GEN_1521 = _GEN_2810 == 8'h1d ? _GEN_1517 : _GEN_1241; // @[executor.scala 473:84]
  wire [7:0] _GEN_1522 = _GEN_2810 == 8'h1d ? _GEN_1518 : _GEN_1242; // @[executor.scala 473:84]
  wire [7:0] _GEN_1523 = _GEN_2810 == 8'h1d ? _GEN_1519 : _GEN_1243; // @[executor.scala 473:84]
  wire [7:0] _GEN_1524 = mask_2[0] ? byte_320 : _GEN_1244; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1525 = mask_2[1] ? byte_321 : _GEN_1245; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1526 = mask_2[2] ? byte_322 : _GEN_1246; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1527 = mask_2[3] ? byte_323 : _GEN_1247; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1528 = _GEN_2810 == 8'h1e ? _GEN_1524 : _GEN_1244; // @[executor.scala 473:84]
  wire [7:0] _GEN_1529 = _GEN_2810 == 8'h1e ? _GEN_1525 : _GEN_1245; // @[executor.scala 473:84]
  wire [7:0] _GEN_1530 = _GEN_2810 == 8'h1e ? _GEN_1526 : _GEN_1246; // @[executor.scala 473:84]
  wire [7:0] _GEN_1531 = _GEN_2810 == 8'h1e ? _GEN_1527 : _GEN_1247; // @[executor.scala 473:84]
  wire [7:0] _GEN_1532 = mask_2[0] ? byte_320 : _GEN_1248; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1533 = mask_2[1] ? byte_321 : _GEN_1249; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1534 = mask_2[2] ? byte_322 : _GEN_1250; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1535 = mask_2[3] ? byte_323 : _GEN_1251; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1536 = _GEN_2810 == 8'h1f ? _GEN_1532 : _GEN_1248; // @[executor.scala 473:84]
  wire [7:0] _GEN_1537 = _GEN_2810 == 8'h1f ? _GEN_1533 : _GEN_1249; // @[executor.scala 473:84]
  wire [7:0] _GEN_1538 = _GEN_2810 == 8'h1f ? _GEN_1534 : _GEN_1250; // @[executor.scala 473:84]
  wire [7:0] _GEN_1539 = _GEN_2810 == 8'h1f ? _GEN_1535 : _GEN_1251; // @[executor.scala 473:84]
  wire [7:0] _GEN_1540 = mask_2[0] ? byte_320 : _GEN_1252; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1541 = mask_2[1] ? byte_321 : _GEN_1253; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1542 = mask_2[2] ? byte_322 : _GEN_1254; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1543 = mask_2[3] ? byte_323 : _GEN_1255; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1544 = _GEN_2810 == 8'h20 ? _GEN_1540 : _GEN_1252; // @[executor.scala 473:84]
  wire [7:0] _GEN_1545 = _GEN_2810 == 8'h20 ? _GEN_1541 : _GEN_1253; // @[executor.scala 473:84]
  wire [7:0] _GEN_1546 = _GEN_2810 == 8'h20 ? _GEN_1542 : _GEN_1254; // @[executor.scala 473:84]
  wire [7:0] _GEN_1547 = _GEN_2810 == 8'h20 ? _GEN_1543 : _GEN_1255; // @[executor.scala 473:84]
  wire [7:0] _GEN_1548 = mask_2[0] ? byte_320 : _GEN_1256; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1549 = mask_2[1] ? byte_321 : _GEN_1257; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1550 = mask_2[2] ? byte_322 : _GEN_1258; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1551 = mask_2[3] ? byte_323 : _GEN_1259; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1552 = _GEN_2810 == 8'h21 ? _GEN_1548 : _GEN_1256; // @[executor.scala 473:84]
  wire [7:0] _GEN_1553 = _GEN_2810 == 8'h21 ? _GEN_1549 : _GEN_1257; // @[executor.scala 473:84]
  wire [7:0] _GEN_1554 = _GEN_2810 == 8'h21 ? _GEN_1550 : _GEN_1258; // @[executor.scala 473:84]
  wire [7:0] _GEN_1555 = _GEN_2810 == 8'h21 ? _GEN_1551 : _GEN_1259; // @[executor.scala 473:84]
  wire [7:0] _GEN_1556 = mask_2[0] ? byte_320 : _GEN_1260; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1557 = mask_2[1] ? byte_321 : _GEN_1261; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1558 = mask_2[2] ? byte_322 : _GEN_1262; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1559 = mask_2[3] ? byte_323 : _GEN_1263; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1560 = _GEN_2810 == 8'h22 ? _GEN_1556 : _GEN_1260; // @[executor.scala 473:84]
  wire [7:0] _GEN_1561 = _GEN_2810 == 8'h22 ? _GEN_1557 : _GEN_1261; // @[executor.scala 473:84]
  wire [7:0] _GEN_1562 = _GEN_2810 == 8'h22 ? _GEN_1558 : _GEN_1262; // @[executor.scala 473:84]
  wire [7:0] _GEN_1563 = _GEN_2810 == 8'h22 ? _GEN_1559 : _GEN_1263; // @[executor.scala 473:84]
  wire [7:0] _GEN_1564 = mask_2[0] ? byte_320 : _GEN_1264; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1565 = mask_2[1] ? byte_321 : _GEN_1265; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1566 = mask_2[2] ? byte_322 : _GEN_1266; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1567 = mask_2[3] ? byte_323 : _GEN_1267; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1568 = _GEN_2810 == 8'h23 ? _GEN_1564 : _GEN_1264; // @[executor.scala 473:84]
  wire [7:0] _GEN_1569 = _GEN_2810 == 8'h23 ? _GEN_1565 : _GEN_1265; // @[executor.scala 473:84]
  wire [7:0] _GEN_1570 = _GEN_2810 == 8'h23 ? _GEN_1566 : _GEN_1266; // @[executor.scala 473:84]
  wire [7:0] _GEN_1571 = _GEN_2810 == 8'h23 ? _GEN_1567 : _GEN_1267; // @[executor.scala 473:84]
  wire [7:0] _GEN_1572 = mask_2[0] ? byte_320 : _GEN_1268; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1573 = mask_2[1] ? byte_321 : _GEN_1269; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1574 = mask_2[2] ? byte_322 : _GEN_1270; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1575 = mask_2[3] ? byte_323 : _GEN_1271; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1576 = _GEN_2810 == 8'h24 ? _GEN_1572 : _GEN_1268; // @[executor.scala 473:84]
  wire [7:0] _GEN_1577 = _GEN_2810 == 8'h24 ? _GEN_1573 : _GEN_1269; // @[executor.scala 473:84]
  wire [7:0] _GEN_1578 = _GEN_2810 == 8'h24 ? _GEN_1574 : _GEN_1270; // @[executor.scala 473:84]
  wire [7:0] _GEN_1579 = _GEN_2810 == 8'h24 ? _GEN_1575 : _GEN_1271; // @[executor.scala 473:84]
  wire [7:0] _GEN_1580 = mask_2[0] ? byte_320 : _GEN_1272; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1581 = mask_2[1] ? byte_321 : _GEN_1273; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1582 = mask_2[2] ? byte_322 : _GEN_1274; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1583 = mask_2[3] ? byte_323 : _GEN_1275; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1584 = _GEN_2810 == 8'h25 ? _GEN_1580 : _GEN_1272; // @[executor.scala 473:84]
  wire [7:0] _GEN_1585 = _GEN_2810 == 8'h25 ? _GEN_1581 : _GEN_1273; // @[executor.scala 473:84]
  wire [7:0] _GEN_1586 = _GEN_2810 == 8'h25 ? _GEN_1582 : _GEN_1274; // @[executor.scala 473:84]
  wire [7:0] _GEN_1587 = _GEN_2810 == 8'h25 ? _GEN_1583 : _GEN_1275; // @[executor.scala 473:84]
  wire [7:0] _GEN_1588 = mask_2[0] ? byte_320 : _GEN_1276; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1589 = mask_2[1] ? byte_321 : _GEN_1277; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1590 = mask_2[2] ? byte_322 : _GEN_1278; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1591 = mask_2[3] ? byte_323 : _GEN_1279; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1592 = _GEN_2810 == 8'h26 ? _GEN_1588 : _GEN_1276; // @[executor.scala 473:84]
  wire [7:0] _GEN_1593 = _GEN_2810 == 8'h26 ? _GEN_1589 : _GEN_1277; // @[executor.scala 473:84]
  wire [7:0] _GEN_1594 = _GEN_2810 == 8'h26 ? _GEN_1590 : _GEN_1278; // @[executor.scala 473:84]
  wire [7:0] _GEN_1595 = _GEN_2810 == 8'h26 ? _GEN_1591 : _GEN_1279; // @[executor.scala 473:84]
  wire [7:0] _GEN_1596 = mask_2[0] ? byte_320 : _GEN_1280; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1597 = mask_2[1] ? byte_321 : _GEN_1281; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1598 = mask_2[2] ? byte_322 : _GEN_1282; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1599 = mask_2[3] ? byte_323 : _GEN_1283; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1600 = _GEN_2810 == 8'h27 ? _GEN_1596 : _GEN_1280; // @[executor.scala 473:84]
  wire [7:0] _GEN_1601 = _GEN_2810 == 8'h27 ? _GEN_1597 : _GEN_1281; // @[executor.scala 473:84]
  wire [7:0] _GEN_1602 = _GEN_2810 == 8'h27 ? _GEN_1598 : _GEN_1282; // @[executor.scala 473:84]
  wire [7:0] _GEN_1603 = _GEN_2810 == 8'h27 ? _GEN_1599 : _GEN_1283; // @[executor.scala 473:84]
  wire [7:0] _GEN_1604 = opcode_2 != 4'h0 ? _GEN_1288 : _GEN_1124; // @[executor.scala 470:55]
  wire [7:0] _GEN_1605 = opcode_2 != 4'h0 ? _GEN_1289 : _GEN_1125; // @[executor.scala 470:55]
  wire [7:0] _GEN_1606 = opcode_2 != 4'h0 ? _GEN_1290 : _GEN_1126; // @[executor.scala 470:55]
  wire [7:0] _GEN_1607 = opcode_2 != 4'h0 ? _GEN_1291 : _GEN_1127; // @[executor.scala 470:55]
  wire [7:0] _GEN_1608 = opcode_2 != 4'h0 ? _GEN_1296 : _GEN_1128; // @[executor.scala 470:55]
  wire [7:0] _GEN_1609 = opcode_2 != 4'h0 ? _GEN_1297 : _GEN_1129; // @[executor.scala 470:55]
  wire [7:0] _GEN_1610 = opcode_2 != 4'h0 ? _GEN_1298 : _GEN_1130; // @[executor.scala 470:55]
  wire [7:0] _GEN_1611 = opcode_2 != 4'h0 ? _GEN_1299 : _GEN_1131; // @[executor.scala 470:55]
  wire [7:0] _GEN_1612 = opcode_2 != 4'h0 ? _GEN_1304 : _GEN_1132; // @[executor.scala 470:55]
  wire [7:0] _GEN_1613 = opcode_2 != 4'h0 ? _GEN_1305 : _GEN_1133; // @[executor.scala 470:55]
  wire [7:0] _GEN_1614 = opcode_2 != 4'h0 ? _GEN_1306 : _GEN_1134; // @[executor.scala 470:55]
  wire [7:0] _GEN_1615 = opcode_2 != 4'h0 ? _GEN_1307 : _GEN_1135; // @[executor.scala 470:55]
  wire [7:0] _GEN_1616 = opcode_2 != 4'h0 ? _GEN_1312 : _GEN_1136; // @[executor.scala 470:55]
  wire [7:0] _GEN_1617 = opcode_2 != 4'h0 ? _GEN_1313 : _GEN_1137; // @[executor.scala 470:55]
  wire [7:0] _GEN_1618 = opcode_2 != 4'h0 ? _GEN_1314 : _GEN_1138; // @[executor.scala 470:55]
  wire [7:0] _GEN_1619 = opcode_2 != 4'h0 ? _GEN_1315 : _GEN_1139; // @[executor.scala 470:55]
  wire [7:0] _GEN_1620 = opcode_2 != 4'h0 ? _GEN_1320 : _GEN_1140; // @[executor.scala 470:55]
  wire [7:0] _GEN_1621 = opcode_2 != 4'h0 ? _GEN_1321 : _GEN_1141; // @[executor.scala 470:55]
  wire [7:0] _GEN_1622 = opcode_2 != 4'h0 ? _GEN_1322 : _GEN_1142; // @[executor.scala 470:55]
  wire [7:0] _GEN_1623 = opcode_2 != 4'h0 ? _GEN_1323 : _GEN_1143; // @[executor.scala 470:55]
  wire [7:0] _GEN_1624 = opcode_2 != 4'h0 ? _GEN_1328 : _GEN_1144; // @[executor.scala 470:55]
  wire [7:0] _GEN_1625 = opcode_2 != 4'h0 ? _GEN_1329 : _GEN_1145; // @[executor.scala 470:55]
  wire [7:0] _GEN_1626 = opcode_2 != 4'h0 ? _GEN_1330 : _GEN_1146; // @[executor.scala 470:55]
  wire [7:0] _GEN_1627 = opcode_2 != 4'h0 ? _GEN_1331 : _GEN_1147; // @[executor.scala 470:55]
  wire [7:0] _GEN_1628 = opcode_2 != 4'h0 ? _GEN_1336 : _GEN_1148; // @[executor.scala 470:55]
  wire [7:0] _GEN_1629 = opcode_2 != 4'h0 ? _GEN_1337 : _GEN_1149; // @[executor.scala 470:55]
  wire [7:0] _GEN_1630 = opcode_2 != 4'h0 ? _GEN_1338 : _GEN_1150; // @[executor.scala 470:55]
  wire [7:0] _GEN_1631 = opcode_2 != 4'h0 ? _GEN_1339 : _GEN_1151; // @[executor.scala 470:55]
  wire [7:0] _GEN_1632 = opcode_2 != 4'h0 ? _GEN_1344 : _GEN_1152; // @[executor.scala 470:55]
  wire [7:0] _GEN_1633 = opcode_2 != 4'h0 ? _GEN_1345 : _GEN_1153; // @[executor.scala 470:55]
  wire [7:0] _GEN_1634 = opcode_2 != 4'h0 ? _GEN_1346 : _GEN_1154; // @[executor.scala 470:55]
  wire [7:0] _GEN_1635 = opcode_2 != 4'h0 ? _GEN_1347 : _GEN_1155; // @[executor.scala 470:55]
  wire [7:0] _GEN_1636 = opcode_2 != 4'h0 ? _GEN_1352 : _GEN_1156; // @[executor.scala 470:55]
  wire [7:0] _GEN_1637 = opcode_2 != 4'h0 ? _GEN_1353 : _GEN_1157; // @[executor.scala 470:55]
  wire [7:0] _GEN_1638 = opcode_2 != 4'h0 ? _GEN_1354 : _GEN_1158; // @[executor.scala 470:55]
  wire [7:0] _GEN_1639 = opcode_2 != 4'h0 ? _GEN_1355 : _GEN_1159; // @[executor.scala 470:55]
  wire [7:0] _GEN_1640 = opcode_2 != 4'h0 ? _GEN_1360 : _GEN_1160; // @[executor.scala 470:55]
  wire [7:0] _GEN_1641 = opcode_2 != 4'h0 ? _GEN_1361 : _GEN_1161; // @[executor.scala 470:55]
  wire [7:0] _GEN_1642 = opcode_2 != 4'h0 ? _GEN_1362 : _GEN_1162; // @[executor.scala 470:55]
  wire [7:0] _GEN_1643 = opcode_2 != 4'h0 ? _GEN_1363 : _GEN_1163; // @[executor.scala 470:55]
  wire [7:0] _GEN_1644 = opcode_2 != 4'h0 ? _GEN_1368 : _GEN_1164; // @[executor.scala 470:55]
  wire [7:0] _GEN_1645 = opcode_2 != 4'h0 ? _GEN_1369 : _GEN_1165; // @[executor.scala 470:55]
  wire [7:0] _GEN_1646 = opcode_2 != 4'h0 ? _GEN_1370 : _GEN_1166; // @[executor.scala 470:55]
  wire [7:0] _GEN_1647 = opcode_2 != 4'h0 ? _GEN_1371 : _GEN_1167; // @[executor.scala 470:55]
  wire [7:0] _GEN_1648 = opcode_2 != 4'h0 ? _GEN_1376 : _GEN_1168; // @[executor.scala 470:55]
  wire [7:0] _GEN_1649 = opcode_2 != 4'h0 ? _GEN_1377 : _GEN_1169; // @[executor.scala 470:55]
  wire [7:0] _GEN_1650 = opcode_2 != 4'h0 ? _GEN_1378 : _GEN_1170; // @[executor.scala 470:55]
  wire [7:0] _GEN_1651 = opcode_2 != 4'h0 ? _GEN_1379 : _GEN_1171; // @[executor.scala 470:55]
  wire [7:0] _GEN_1652 = opcode_2 != 4'h0 ? _GEN_1384 : _GEN_1172; // @[executor.scala 470:55]
  wire [7:0] _GEN_1653 = opcode_2 != 4'h0 ? _GEN_1385 : _GEN_1173; // @[executor.scala 470:55]
  wire [7:0] _GEN_1654 = opcode_2 != 4'h0 ? _GEN_1386 : _GEN_1174; // @[executor.scala 470:55]
  wire [7:0] _GEN_1655 = opcode_2 != 4'h0 ? _GEN_1387 : _GEN_1175; // @[executor.scala 470:55]
  wire [7:0] _GEN_1656 = opcode_2 != 4'h0 ? _GEN_1392 : _GEN_1176; // @[executor.scala 470:55]
  wire [7:0] _GEN_1657 = opcode_2 != 4'h0 ? _GEN_1393 : _GEN_1177; // @[executor.scala 470:55]
  wire [7:0] _GEN_1658 = opcode_2 != 4'h0 ? _GEN_1394 : _GEN_1178; // @[executor.scala 470:55]
  wire [7:0] _GEN_1659 = opcode_2 != 4'h0 ? _GEN_1395 : _GEN_1179; // @[executor.scala 470:55]
  wire [7:0] _GEN_1660 = opcode_2 != 4'h0 ? _GEN_1400 : _GEN_1180; // @[executor.scala 470:55]
  wire [7:0] _GEN_1661 = opcode_2 != 4'h0 ? _GEN_1401 : _GEN_1181; // @[executor.scala 470:55]
  wire [7:0] _GEN_1662 = opcode_2 != 4'h0 ? _GEN_1402 : _GEN_1182; // @[executor.scala 470:55]
  wire [7:0] _GEN_1663 = opcode_2 != 4'h0 ? _GEN_1403 : _GEN_1183; // @[executor.scala 470:55]
  wire [7:0] _GEN_1664 = opcode_2 != 4'h0 ? _GEN_1408 : _GEN_1184; // @[executor.scala 470:55]
  wire [7:0] _GEN_1665 = opcode_2 != 4'h0 ? _GEN_1409 : _GEN_1185; // @[executor.scala 470:55]
  wire [7:0] _GEN_1666 = opcode_2 != 4'h0 ? _GEN_1410 : _GEN_1186; // @[executor.scala 470:55]
  wire [7:0] _GEN_1667 = opcode_2 != 4'h0 ? _GEN_1411 : _GEN_1187; // @[executor.scala 470:55]
  wire [7:0] _GEN_1668 = opcode_2 != 4'h0 ? _GEN_1416 : _GEN_1188; // @[executor.scala 470:55]
  wire [7:0] _GEN_1669 = opcode_2 != 4'h0 ? _GEN_1417 : _GEN_1189; // @[executor.scala 470:55]
  wire [7:0] _GEN_1670 = opcode_2 != 4'h0 ? _GEN_1418 : _GEN_1190; // @[executor.scala 470:55]
  wire [7:0] _GEN_1671 = opcode_2 != 4'h0 ? _GEN_1419 : _GEN_1191; // @[executor.scala 470:55]
  wire [7:0] _GEN_1672 = opcode_2 != 4'h0 ? _GEN_1424 : _GEN_1192; // @[executor.scala 470:55]
  wire [7:0] _GEN_1673 = opcode_2 != 4'h0 ? _GEN_1425 : _GEN_1193; // @[executor.scala 470:55]
  wire [7:0] _GEN_1674 = opcode_2 != 4'h0 ? _GEN_1426 : _GEN_1194; // @[executor.scala 470:55]
  wire [7:0] _GEN_1675 = opcode_2 != 4'h0 ? _GEN_1427 : _GEN_1195; // @[executor.scala 470:55]
  wire [7:0] _GEN_1676 = opcode_2 != 4'h0 ? _GEN_1432 : _GEN_1196; // @[executor.scala 470:55]
  wire [7:0] _GEN_1677 = opcode_2 != 4'h0 ? _GEN_1433 : _GEN_1197; // @[executor.scala 470:55]
  wire [7:0] _GEN_1678 = opcode_2 != 4'h0 ? _GEN_1434 : _GEN_1198; // @[executor.scala 470:55]
  wire [7:0] _GEN_1679 = opcode_2 != 4'h0 ? _GEN_1435 : _GEN_1199; // @[executor.scala 470:55]
  wire [7:0] _GEN_1680 = opcode_2 != 4'h0 ? _GEN_1440 : _GEN_1200; // @[executor.scala 470:55]
  wire [7:0] _GEN_1681 = opcode_2 != 4'h0 ? _GEN_1441 : _GEN_1201; // @[executor.scala 470:55]
  wire [7:0] _GEN_1682 = opcode_2 != 4'h0 ? _GEN_1442 : _GEN_1202; // @[executor.scala 470:55]
  wire [7:0] _GEN_1683 = opcode_2 != 4'h0 ? _GEN_1443 : _GEN_1203; // @[executor.scala 470:55]
  wire [7:0] _GEN_1684 = opcode_2 != 4'h0 ? _GEN_1448 : _GEN_1204; // @[executor.scala 470:55]
  wire [7:0] _GEN_1685 = opcode_2 != 4'h0 ? _GEN_1449 : _GEN_1205; // @[executor.scala 470:55]
  wire [7:0] _GEN_1686 = opcode_2 != 4'h0 ? _GEN_1450 : _GEN_1206; // @[executor.scala 470:55]
  wire [7:0] _GEN_1687 = opcode_2 != 4'h0 ? _GEN_1451 : _GEN_1207; // @[executor.scala 470:55]
  wire [7:0] _GEN_1688 = opcode_2 != 4'h0 ? _GEN_1456 : _GEN_1208; // @[executor.scala 470:55]
  wire [7:0] _GEN_1689 = opcode_2 != 4'h0 ? _GEN_1457 : _GEN_1209; // @[executor.scala 470:55]
  wire [7:0] _GEN_1690 = opcode_2 != 4'h0 ? _GEN_1458 : _GEN_1210; // @[executor.scala 470:55]
  wire [7:0] _GEN_1691 = opcode_2 != 4'h0 ? _GEN_1459 : _GEN_1211; // @[executor.scala 470:55]
  wire [7:0] _GEN_1692 = opcode_2 != 4'h0 ? _GEN_1464 : _GEN_1212; // @[executor.scala 470:55]
  wire [7:0] _GEN_1693 = opcode_2 != 4'h0 ? _GEN_1465 : _GEN_1213; // @[executor.scala 470:55]
  wire [7:0] _GEN_1694 = opcode_2 != 4'h0 ? _GEN_1466 : _GEN_1214; // @[executor.scala 470:55]
  wire [7:0] _GEN_1695 = opcode_2 != 4'h0 ? _GEN_1467 : _GEN_1215; // @[executor.scala 470:55]
  wire [7:0] _GEN_1696 = opcode_2 != 4'h0 ? _GEN_1472 : _GEN_1216; // @[executor.scala 470:55]
  wire [7:0] _GEN_1697 = opcode_2 != 4'h0 ? _GEN_1473 : _GEN_1217; // @[executor.scala 470:55]
  wire [7:0] _GEN_1698 = opcode_2 != 4'h0 ? _GEN_1474 : _GEN_1218; // @[executor.scala 470:55]
  wire [7:0] _GEN_1699 = opcode_2 != 4'h0 ? _GEN_1475 : _GEN_1219; // @[executor.scala 470:55]
  wire [7:0] _GEN_1700 = opcode_2 != 4'h0 ? _GEN_1480 : _GEN_1220; // @[executor.scala 470:55]
  wire [7:0] _GEN_1701 = opcode_2 != 4'h0 ? _GEN_1481 : _GEN_1221; // @[executor.scala 470:55]
  wire [7:0] _GEN_1702 = opcode_2 != 4'h0 ? _GEN_1482 : _GEN_1222; // @[executor.scala 470:55]
  wire [7:0] _GEN_1703 = opcode_2 != 4'h0 ? _GEN_1483 : _GEN_1223; // @[executor.scala 470:55]
  wire [7:0] _GEN_1704 = opcode_2 != 4'h0 ? _GEN_1488 : _GEN_1224; // @[executor.scala 470:55]
  wire [7:0] _GEN_1705 = opcode_2 != 4'h0 ? _GEN_1489 : _GEN_1225; // @[executor.scala 470:55]
  wire [7:0] _GEN_1706 = opcode_2 != 4'h0 ? _GEN_1490 : _GEN_1226; // @[executor.scala 470:55]
  wire [7:0] _GEN_1707 = opcode_2 != 4'h0 ? _GEN_1491 : _GEN_1227; // @[executor.scala 470:55]
  wire [7:0] _GEN_1708 = opcode_2 != 4'h0 ? _GEN_1496 : _GEN_1228; // @[executor.scala 470:55]
  wire [7:0] _GEN_1709 = opcode_2 != 4'h0 ? _GEN_1497 : _GEN_1229; // @[executor.scala 470:55]
  wire [7:0] _GEN_1710 = opcode_2 != 4'h0 ? _GEN_1498 : _GEN_1230; // @[executor.scala 470:55]
  wire [7:0] _GEN_1711 = opcode_2 != 4'h0 ? _GEN_1499 : _GEN_1231; // @[executor.scala 470:55]
  wire [7:0] _GEN_1712 = opcode_2 != 4'h0 ? _GEN_1504 : _GEN_1232; // @[executor.scala 470:55]
  wire [7:0] _GEN_1713 = opcode_2 != 4'h0 ? _GEN_1505 : _GEN_1233; // @[executor.scala 470:55]
  wire [7:0] _GEN_1714 = opcode_2 != 4'h0 ? _GEN_1506 : _GEN_1234; // @[executor.scala 470:55]
  wire [7:0] _GEN_1715 = opcode_2 != 4'h0 ? _GEN_1507 : _GEN_1235; // @[executor.scala 470:55]
  wire [7:0] _GEN_1716 = opcode_2 != 4'h0 ? _GEN_1512 : _GEN_1236; // @[executor.scala 470:55]
  wire [7:0] _GEN_1717 = opcode_2 != 4'h0 ? _GEN_1513 : _GEN_1237; // @[executor.scala 470:55]
  wire [7:0] _GEN_1718 = opcode_2 != 4'h0 ? _GEN_1514 : _GEN_1238; // @[executor.scala 470:55]
  wire [7:0] _GEN_1719 = opcode_2 != 4'h0 ? _GEN_1515 : _GEN_1239; // @[executor.scala 470:55]
  wire [7:0] _GEN_1720 = opcode_2 != 4'h0 ? _GEN_1520 : _GEN_1240; // @[executor.scala 470:55]
  wire [7:0] _GEN_1721 = opcode_2 != 4'h0 ? _GEN_1521 : _GEN_1241; // @[executor.scala 470:55]
  wire [7:0] _GEN_1722 = opcode_2 != 4'h0 ? _GEN_1522 : _GEN_1242; // @[executor.scala 470:55]
  wire [7:0] _GEN_1723 = opcode_2 != 4'h0 ? _GEN_1523 : _GEN_1243; // @[executor.scala 470:55]
  wire [7:0] _GEN_1724 = opcode_2 != 4'h0 ? _GEN_1528 : _GEN_1244; // @[executor.scala 470:55]
  wire [7:0] _GEN_1725 = opcode_2 != 4'h0 ? _GEN_1529 : _GEN_1245; // @[executor.scala 470:55]
  wire [7:0] _GEN_1726 = opcode_2 != 4'h0 ? _GEN_1530 : _GEN_1246; // @[executor.scala 470:55]
  wire [7:0] _GEN_1727 = opcode_2 != 4'h0 ? _GEN_1531 : _GEN_1247; // @[executor.scala 470:55]
  wire [7:0] _GEN_1728 = opcode_2 != 4'h0 ? _GEN_1536 : _GEN_1248; // @[executor.scala 470:55]
  wire [7:0] _GEN_1729 = opcode_2 != 4'h0 ? _GEN_1537 : _GEN_1249; // @[executor.scala 470:55]
  wire [7:0] _GEN_1730 = opcode_2 != 4'h0 ? _GEN_1538 : _GEN_1250; // @[executor.scala 470:55]
  wire [7:0] _GEN_1731 = opcode_2 != 4'h0 ? _GEN_1539 : _GEN_1251; // @[executor.scala 470:55]
  wire [7:0] _GEN_1732 = opcode_2 != 4'h0 ? _GEN_1544 : _GEN_1252; // @[executor.scala 470:55]
  wire [7:0] _GEN_1733 = opcode_2 != 4'h0 ? _GEN_1545 : _GEN_1253; // @[executor.scala 470:55]
  wire [7:0] _GEN_1734 = opcode_2 != 4'h0 ? _GEN_1546 : _GEN_1254; // @[executor.scala 470:55]
  wire [7:0] _GEN_1735 = opcode_2 != 4'h0 ? _GEN_1547 : _GEN_1255; // @[executor.scala 470:55]
  wire [7:0] _GEN_1736 = opcode_2 != 4'h0 ? _GEN_1552 : _GEN_1256; // @[executor.scala 470:55]
  wire [7:0] _GEN_1737 = opcode_2 != 4'h0 ? _GEN_1553 : _GEN_1257; // @[executor.scala 470:55]
  wire [7:0] _GEN_1738 = opcode_2 != 4'h0 ? _GEN_1554 : _GEN_1258; // @[executor.scala 470:55]
  wire [7:0] _GEN_1739 = opcode_2 != 4'h0 ? _GEN_1555 : _GEN_1259; // @[executor.scala 470:55]
  wire [7:0] _GEN_1740 = opcode_2 != 4'h0 ? _GEN_1560 : _GEN_1260; // @[executor.scala 470:55]
  wire [7:0] _GEN_1741 = opcode_2 != 4'h0 ? _GEN_1561 : _GEN_1261; // @[executor.scala 470:55]
  wire [7:0] _GEN_1742 = opcode_2 != 4'h0 ? _GEN_1562 : _GEN_1262; // @[executor.scala 470:55]
  wire [7:0] _GEN_1743 = opcode_2 != 4'h0 ? _GEN_1563 : _GEN_1263; // @[executor.scala 470:55]
  wire [7:0] _GEN_1744 = opcode_2 != 4'h0 ? _GEN_1568 : _GEN_1264; // @[executor.scala 470:55]
  wire [7:0] _GEN_1745 = opcode_2 != 4'h0 ? _GEN_1569 : _GEN_1265; // @[executor.scala 470:55]
  wire [7:0] _GEN_1746 = opcode_2 != 4'h0 ? _GEN_1570 : _GEN_1266; // @[executor.scala 470:55]
  wire [7:0] _GEN_1747 = opcode_2 != 4'h0 ? _GEN_1571 : _GEN_1267; // @[executor.scala 470:55]
  wire [7:0] _GEN_1748 = opcode_2 != 4'h0 ? _GEN_1576 : _GEN_1268; // @[executor.scala 470:55]
  wire [7:0] _GEN_1749 = opcode_2 != 4'h0 ? _GEN_1577 : _GEN_1269; // @[executor.scala 470:55]
  wire [7:0] _GEN_1750 = opcode_2 != 4'h0 ? _GEN_1578 : _GEN_1270; // @[executor.scala 470:55]
  wire [7:0] _GEN_1751 = opcode_2 != 4'h0 ? _GEN_1579 : _GEN_1271; // @[executor.scala 470:55]
  wire [7:0] _GEN_1752 = opcode_2 != 4'h0 ? _GEN_1584 : _GEN_1272; // @[executor.scala 470:55]
  wire [7:0] _GEN_1753 = opcode_2 != 4'h0 ? _GEN_1585 : _GEN_1273; // @[executor.scala 470:55]
  wire [7:0] _GEN_1754 = opcode_2 != 4'h0 ? _GEN_1586 : _GEN_1274; // @[executor.scala 470:55]
  wire [7:0] _GEN_1755 = opcode_2 != 4'h0 ? _GEN_1587 : _GEN_1275; // @[executor.scala 470:55]
  wire [7:0] _GEN_1756 = opcode_2 != 4'h0 ? _GEN_1592 : _GEN_1276; // @[executor.scala 470:55]
  wire [7:0] _GEN_1757 = opcode_2 != 4'h0 ? _GEN_1593 : _GEN_1277; // @[executor.scala 470:55]
  wire [7:0] _GEN_1758 = opcode_2 != 4'h0 ? _GEN_1594 : _GEN_1278; // @[executor.scala 470:55]
  wire [7:0] _GEN_1759 = opcode_2 != 4'h0 ? _GEN_1595 : _GEN_1279; // @[executor.scala 470:55]
  wire [7:0] _GEN_1760 = opcode_2 != 4'h0 ? _GEN_1600 : _GEN_1280; // @[executor.scala 470:55]
  wire [7:0] _GEN_1761 = opcode_2 != 4'h0 ? _GEN_1601 : _GEN_1281; // @[executor.scala 470:55]
  wire [7:0] _GEN_1762 = opcode_2 != 4'h0 ? _GEN_1602 : _GEN_1282; // @[executor.scala 470:55]
  wire [7:0] _GEN_1763 = opcode_2 != 4'h0 ? _GEN_1603 : _GEN_1283; // @[executor.scala 470:55]
  wire [3:0] _GEN_1764 = opcode_2 == 4'hf ? parameter_2_2[13:10] : _GEN_1122; // @[executor.scala 466:52 executor.scala 467:55]
  wire  _GEN_1765 = opcode_2 == 4'hf ? parameter_2_2[0] : _GEN_1123; // @[executor.scala 466:52 executor.scala 468:55]
  wire [7:0] _GEN_1766 = opcode_2 == 4'hf ? _GEN_1124 : _GEN_1604; // @[executor.scala 466:52]
  wire [7:0] _GEN_1767 = opcode_2 == 4'hf ? _GEN_1125 : _GEN_1605; // @[executor.scala 466:52]
  wire [7:0] _GEN_1768 = opcode_2 == 4'hf ? _GEN_1126 : _GEN_1606; // @[executor.scala 466:52]
  wire [7:0] _GEN_1769 = opcode_2 == 4'hf ? _GEN_1127 : _GEN_1607; // @[executor.scala 466:52]
  wire [7:0] _GEN_1770 = opcode_2 == 4'hf ? _GEN_1128 : _GEN_1608; // @[executor.scala 466:52]
  wire [7:0] _GEN_1771 = opcode_2 == 4'hf ? _GEN_1129 : _GEN_1609; // @[executor.scala 466:52]
  wire [7:0] _GEN_1772 = opcode_2 == 4'hf ? _GEN_1130 : _GEN_1610; // @[executor.scala 466:52]
  wire [7:0] _GEN_1773 = opcode_2 == 4'hf ? _GEN_1131 : _GEN_1611; // @[executor.scala 466:52]
  wire [7:0] _GEN_1774 = opcode_2 == 4'hf ? _GEN_1132 : _GEN_1612; // @[executor.scala 466:52]
  wire [7:0] _GEN_1775 = opcode_2 == 4'hf ? _GEN_1133 : _GEN_1613; // @[executor.scala 466:52]
  wire [7:0] _GEN_1776 = opcode_2 == 4'hf ? _GEN_1134 : _GEN_1614; // @[executor.scala 466:52]
  wire [7:0] _GEN_1777 = opcode_2 == 4'hf ? _GEN_1135 : _GEN_1615; // @[executor.scala 466:52]
  wire [7:0] _GEN_1778 = opcode_2 == 4'hf ? _GEN_1136 : _GEN_1616; // @[executor.scala 466:52]
  wire [7:0] _GEN_1779 = opcode_2 == 4'hf ? _GEN_1137 : _GEN_1617; // @[executor.scala 466:52]
  wire [7:0] _GEN_1780 = opcode_2 == 4'hf ? _GEN_1138 : _GEN_1618; // @[executor.scala 466:52]
  wire [7:0] _GEN_1781 = opcode_2 == 4'hf ? _GEN_1139 : _GEN_1619; // @[executor.scala 466:52]
  wire [7:0] _GEN_1782 = opcode_2 == 4'hf ? _GEN_1140 : _GEN_1620; // @[executor.scala 466:52]
  wire [7:0] _GEN_1783 = opcode_2 == 4'hf ? _GEN_1141 : _GEN_1621; // @[executor.scala 466:52]
  wire [7:0] _GEN_1784 = opcode_2 == 4'hf ? _GEN_1142 : _GEN_1622; // @[executor.scala 466:52]
  wire [7:0] _GEN_1785 = opcode_2 == 4'hf ? _GEN_1143 : _GEN_1623; // @[executor.scala 466:52]
  wire [7:0] _GEN_1786 = opcode_2 == 4'hf ? _GEN_1144 : _GEN_1624; // @[executor.scala 466:52]
  wire [7:0] _GEN_1787 = opcode_2 == 4'hf ? _GEN_1145 : _GEN_1625; // @[executor.scala 466:52]
  wire [7:0] _GEN_1788 = opcode_2 == 4'hf ? _GEN_1146 : _GEN_1626; // @[executor.scala 466:52]
  wire [7:0] _GEN_1789 = opcode_2 == 4'hf ? _GEN_1147 : _GEN_1627; // @[executor.scala 466:52]
  wire [7:0] _GEN_1790 = opcode_2 == 4'hf ? _GEN_1148 : _GEN_1628; // @[executor.scala 466:52]
  wire [7:0] _GEN_1791 = opcode_2 == 4'hf ? _GEN_1149 : _GEN_1629; // @[executor.scala 466:52]
  wire [7:0] _GEN_1792 = opcode_2 == 4'hf ? _GEN_1150 : _GEN_1630; // @[executor.scala 466:52]
  wire [7:0] _GEN_1793 = opcode_2 == 4'hf ? _GEN_1151 : _GEN_1631; // @[executor.scala 466:52]
  wire [7:0] _GEN_1794 = opcode_2 == 4'hf ? _GEN_1152 : _GEN_1632; // @[executor.scala 466:52]
  wire [7:0] _GEN_1795 = opcode_2 == 4'hf ? _GEN_1153 : _GEN_1633; // @[executor.scala 466:52]
  wire [7:0] _GEN_1796 = opcode_2 == 4'hf ? _GEN_1154 : _GEN_1634; // @[executor.scala 466:52]
  wire [7:0] _GEN_1797 = opcode_2 == 4'hf ? _GEN_1155 : _GEN_1635; // @[executor.scala 466:52]
  wire [7:0] _GEN_1798 = opcode_2 == 4'hf ? _GEN_1156 : _GEN_1636; // @[executor.scala 466:52]
  wire [7:0] _GEN_1799 = opcode_2 == 4'hf ? _GEN_1157 : _GEN_1637; // @[executor.scala 466:52]
  wire [7:0] _GEN_1800 = opcode_2 == 4'hf ? _GEN_1158 : _GEN_1638; // @[executor.scala 466:52]
  wire [7:0] _GEN_1801 = opcode_2 == 4'hf ? _GEN_1159 : _GEN_1639; // @[executor.scala 466:52]
  wire [7:0] _GEN_1802 = opcode_2 == 4'hf ? _GEN_1160 : _GEN_1640; // @[executor.scala 466:52]
  wire [7:0] _GEN_1803 = opcode_2 == 4'hf ? _GEN_1161 : _GEN_1641; // @[executor.scala 466:52]
  wire [7:0] _GEN_1804 = opcode_2 == 4'hf ? _GEN_1162 : _GEN_1642; // @[executor.scala 466:52]
  wire [7:0] _GEN_1805 = opcode_2 == 4'hf ? _GEN_1163 : _GEN_1643; // @[executor.scala 466:52]
  wire [7:0] _GEN_1806 = opcode_2 == 4'hf ? _GEN_1164 : _GEN_1644; // @[executor.scala 466:52]
  wire [7:0] _GEN_1807 = opcode_2 == 4'hf ? _GEN_1165 : _GEN_1645; // @[executor.scala 466:52]
  wire [7:0] _GEN_1808 = opcode_2 == 4'hf ? _GEN_1166 : _GEN_1646; // @[executor.scala 466:52]
  wire [7:0] _GEN_1809 = opcode_2 == 4'hf ? _GEN_1167 : _GEN_1647; // @[executor.scala 466:52]
  wire [7:0] _GEN_1810 = opcode_2 == 4'hf ? _GEN_1168 : _GEN_1648; // @[executor.scala 466:52]
  wire [7:0] _GEN_1811 = opcode_2 == 4'hf ? _GEN_1169 : _GEN_1649; // @[executor.scala 466:52]
  wire [7:0] _GEN_1812 = opcode_2 == 4'hf ? _GEN_1170 : _GEN_1650; // @[executor.scala 466:52]
  wire [7:0] _GEN_1813 = opcode_2 == 4'hf ? _GEN_1171 : _GEN_1651; // @[executor.scala 466:52]
  wire [7:0] _GEN_1814 = opcode_2 == 4'hf ? _GEN_1172 : _GEN_1652; // @[executor.scala 466:52]
  wire [7:0] _GEN_1815 = opcode_2 == 4'hf ? _GEN_1173 : _GEN_1653; // @[executor.scala 466:52]
  wire [7:0] _GEN_1816 = opcode_2 == 4'hf ? _GEN_1174 : _GEN_1654; // @[executor.scala 466:52]
  wire [7:0] _GEN_1817 = opcode_2 == 4'hf ? _GEN_1175 : _GEN_1655; // @[executor.scala 466:52]
  wire [7:0] _GEN_1818 = opcode_2 == 4'hf ? _GEN_1176 : _GEN_1656; // @[executor.scala 466:52]
  wire [7:0] _GEN_1819 = opcode_2 == 4'hf ? _GEN_1177 : _GEN_1657; // @[executor.scala 466:52]
  wire [7:0] _GEN_1820 = opcode_2 == 4'hf ? _GEN_1178 : _GEN_1658; // @[executor.scala 466:52]
  wire [7:0] _GEN_1821 = opcode_2 == 4'hf ? _GEN_1179 : _GEN_1659; // @[executor.scala 466:52]
  wire [7:0] _GEN_1822 = opcode_2 == 4'hf ? _GEN_1180 : _GEN_1660; // @[executor.scala 466:52]
  wire [7:0] _GEN_1823 = opcode_2 == 4'hf ? _GEN_1181 : _GEN_1661; // @[executor.scala 466:52]
  wire [7:0] _GEN_1824 = opcode_2 == 4'hf ? _GEN_1182 : _GEN_1662; // @[executor.scala 466:52]
  wire [7:0] _GEN_1825 = opcode_2 == 4'hf ? _GEN_1183 : _GEN_1663; // @[executor.scala 466:52]
  wire [7:0] _GEN_1826 = opcode_2 == 4'hf ? _GEN_1184 : _GEN_1664; // @[executor.scala 466:52]
  wire [7:0] _GEN_1827 = opcode_2 == 4'hf ? _GEN_1185 : _GEN_1665; // @[executor.scala 466:52]
  wire [7:0] _GEN_1828 = opcode_2 == 4'hf ? _GEN_1186 : _GEN_1666; // @[executor.scala 466:52]
  wire [7:0] _GEN_1829 = opcode_2 == 4'hf ? _GEN_1187 : _GEN_1667; // @[executor.scala 466:52]
  wire [7:0] _GEN_1830 = opcode_2 == 4'hf ? _GEN_1188 : _GEN_1668; // @[executor.scala 466:52]
  wire [7:0] _GEN_1831 = opcode_2 == 4'hf ? _GEN_1189 : _GEN_1669; // @[executor.scala 466:52]
  wire [7:0] _GEN_1832 = opcode_2 == 4'hf ? _GEN_1190 : _GEN_1670; // @[executor.scala 466:52]
  wire [7:0] _GEN_1833 = opcode_2 == 4'hf ? _GEN_1191 : _GEN_1671; // @[executor.scala 466:52]
  wire [7:0] _GEN_1834 = opcode_2 == 4'hf ? _GEN_1192 : _GEN_1672; // @[executor.scala 466:52]
  wire [7:0] _GEN_1835 = opcode_2 == 4'hf ? _GEN_1193 : _GEN_1673; // @[executor.scala 466:52]
  wire [7:0] _GEN_1836 = opcode_2 == 4'hf ? _GEN_1194 : _GEN_1674; // @[executor.scala 466:52]
  wire [7:0] _GEN_1837 = opcode_2 == 4'hf ? _GEN_1195 : _GEN_1675; // @[executor.scala 466:52]
  wire [7:0] _GEN_1838 = opcode_2 == 4'hf ? _GEN_1196 : _GEN_1676; // @[executor.scala 466:52]
  wire [7:0] _GEN_1839 = opcode_2 == 4'hf ? _GEN_1197 : _GEN_1677; // @[executor.scala 466:52]
  wire [7:0] _GEN_1840 = opcode_2 == 4'hf ? _GEN_1198 : _GEN_1678; // @[executor.scala 466:52]
  wire [7:0] _GEN_1841 = opcode_2 == 4'hf ? _GEN_1199 : _GEN_1679; // @[executor.scala 466:52]
  wire [7:0] _GEN_1842 = opcode_2 == 4'hf ? _GEN_1200 : _GEN_1680; // @[executor.scala 466:52]
  wire [7:0] _GEN_1843 = opcode_2 == 4'hf ? _GEN_1201 : _GEN_1681; // @[executor.scala 466:52]
  wire [7:0] _GEN_1844 = opcode_2 == 4'hf ? _GEN_1202 : _GEN_1682; // @[executor.scala 466:52]
  wire [7:0] _GEN_1845 = opcode_2 == 4'hf ? _GEN_1203 : _GEN_1683; // @[executor.scala 466:52]
  wire [7:0] _GEN_1846 = opcode_2 == 4'hf ? _GEN_1204 : _GEN_1684; // @[executor.scala 466:52]
  wire [7:0] _GEN_1847 = opcode_2 == 4'hf ? _GEN_1205 : _GEN_1685; // @[executor.scala 466:52]
  wire [7:0] _GEN_1848 = opcode_2 == 4'hf ? _GEN_1206 : _GEN_1686; // @[executor.scala 466:52]
  wire [7:0] _GEN_1849 = opcode_2 == 4'hf ? _GEN_1207 : _GEN_1687; // @[executor.scala 466:52]
  wire [7:0] _GEN_1850 = opcode_2 == 4'hf ? _GEN_1208 : _GEN_1688; // @[executor.scala 466:52]
  wire [7:0] _GEN_1851 = opcode_2 == 4'hf ? _GEN_1209 : _GEN_1689; // @[executor.scala 466:52]
  wire [7:0] _GEN_1852 = opcode_2 == 4'hf ? _GEN_1210 : _GEN_1690; // @[executor.scala 466:52]
  wire [7:0] _GEN_1853 = opcode_2 == 4'hf ? _GEN_1211 : _GEN_1691; // @[executor.scala 466:52]
  wire [7:0] _GEN_1854 = opcode_2 == 4'hf ? _GEN_1212 : _GEN_1692; // @[executor.scala 466:52]
  wire [7:0] _GEN_1855 = opcode_2 == 4'hf ? _GEN_1213 : _GEN_1693; // @[executor.scala 466:52]
  wire [7:0] _GEN_1856 = opcode_2 == 4'hf ? _GEN_1214 : _GEN_1694; // @[executor.scala 466:52]
  wire [7:0] _GEN_1857 = opcode_2 == 4'hf ? _GEN_1215 : _GEN_1695; // @[executor.scala 466:52]
  wire [7:0] _GEN_1858 = opcode_2 == 4'hf ? _GEN_1216 : _GEN_1696; // @[executor.scala 466:52]
  wire [7:0] _GEN_1859 = opcode_2 == 4'hf ? _GEN_1217 : _GEN_1697; // @[executor.scala 466:52]
  wire [7:0] _GEN_1860 = opcode_2 == 4'hf ? _GEN_1218 : _GEN_1698; // @[executor.scala 466:52]
  wire [7:0] _GEN_1861 = opcode_2 == 4'hf ? _GEN_1219 : _GEN_1699; // @[executor.scala 466:52]
  wire [7:0] _GEN_1862 = opcode_2 == 4'hf ? _GEN_1220 : _GEN_1700; // @[executor.scala 466:52]
  wire [7:0] _GEN_1863 = opcode_2 == 4'hf ? _GEN_1221 : _GEN_1701; // @[executor.scala 466:52]
  wire [7:0] _GEN_1864 = opcode_2 == 4'hf ? _GEN_1222 : _GEN_1702; // @[executor.scala 466:52]
  wire [7:0] _GEN_1865 = opcode_2 == 4'hf ? _GEN_1223 : _GEN_1703; // @[executor.scala 466:52]
  wire [7:0] _GEN_1866 = opcode_2 == 4'hf ? _GEN_1224 : _GEN_1704; // @[executor.scala 466:52]
  wire [7:0] _GEN_1867 = opcode_2 == 4'hf ? _GEN_1225 : _GEN_1705; // @[executor.scala 466:52]
  wire [7:0] _GEN_1868 = opcode_2 == 4'hf ? _GEN_1226 : _GEN_1706; // @[executor.scala 466:52]
  wire [7:0] _GEN_1869 = opcode_2 == 4'hf ? _GEN_1227 : _GEN_1707; // @[executor.scala 466:52]
  wire [7:0] _GEN_1870 = opcode_2 == 4'hf ? _GEN_1228 : _GEN_1708; // @[executor.scala 466:52]
  wire [7:0] _GEN_1871 = opcode_2 == 4'hf ? _GEN_1229 : _GEN_1709; // @[executor.scala 466:52]
  wire [7:0] _GEN_1872 = opcode_2 == 4'hf ? _GEN_1230 : _GEN_1710; // @[executor.scala 466:52]
  wire [7:0] _GEN_1873 = opcode_2 == 4'hf ? _GEN_1231 : _GEN_1711; // @[executor.scala 466:52]
  wire [7:0] _GEN_1874 = opcode_2 == 4'hf ? _GEN_1232 : _GEN_1712; // @[executor.scala 466:52]
  wire [7:0] _GEN_1875 = opcode_2 == 4'hf ? _GEN_1233 : _GEN_1713; // @[executor.scala 466:52]
  wire [7:0] _GEN_1876 = opcode_2 == 4'hf ? _GEN_1234 : _GEN_1714; // @[executor.scala 466:52]
  wire [7:0] _GEN_1877 = opcode_2 == 4'hf ? _GEN_1235 : _GEN_1715; // @[executor.scala 466:52]
  wire [7:0] _GEN_1878 = opcode_2 == 4'hf ? _GEN_1236 : _GEN_1716; // @[executor.scala 466:52]
  wire [7:0] _GEN_1879 = opcode_2 == 4'hf ? _GEN_1237 : _GEN_1717; // @[executor.scala 466:52]
  wire [7:0] _GEN_1880 = opcode_2 == 4'hf ? _GEN_1238 : _GEN_1718; // @[executor.scala 466:52]
  wire [7:0] _GEN_1881 = opcode_2 == 4'hf ? _GEN_1239 : _GEN_1719; // @[executor.scala 466:52]
  wire [7:0] _GEN_1882 = opcode_2 == 4'hf ? _GEN_1240 : _GEN_1720; // @[executor.scala 466:52]
  wire [7:0] _GEN_1883 = opcode_2 == 4'hf ? _GEN_1241 : _GEN_1721; // @[executor.scala 466:52]
  wire [7:0] _GEN_1884 = opcode_2 == 4'hf ? _GEN_1242 : _GEN_1722; // @[executor.scala 466:52]
  wire [7:0] _GEN_1885 = opcode_2 == 4'hf ? _GEN_1243 : _GEN_1723; // @[executor.scala 466:52]
  wire [7:0] _GEN_1886 = opcode_2 == 4'hf ? _GEN_1244 : _GEN_1724; // @[executor.scala 466:52]
  wire [7:0] _GEN_1887 = opcode_2 == 4'hf ? _GEN_1245 : _GEN_1725; // @[executor.scala 466:52]
  wire [7:0] _GEN_1888 = opcode_2 == 4'hf ? _GEN_1246 : _GEN_1726; // @[executor.scala 466:52]
  wire [7:0] _GEN_1889 = opcode_2 == 4'hf ? _GEN_1247 : _GEN_1727; // @[executor.scala 466:52]
  wire [7:0] _GEN_1890 = opcode_2 == 4'hf ? _GEN_1248 : _GEN_1728; // @[executor.scala 466:52]
  wire [7:0] _GEN_1891 = opcode_2 == 4'hf ? _GEN_1249 : _GEN_1729; // @[executor.scala 466:52]
  wire [7:0] _GEN_1892 = opcode_2 == 4'hf ? _GEN_1250 : _GEN_1730; // @[executor.scala 466:52]
  wire [7:0] _GEN_1893 = opcode_2 == 4'hf ? _GEN_1251 : _GEN_1731; // @[executor.scala 466:52]
  wire [7:0] _GEN_1894 = opcode_2 == 4'hf ? _GEN_1252 : _GEN_1732; // @[executor.scala 466:52]
  wire [7:0] _GEN_1895 = opcode_2 == 4'hf ? _GEN_1253 : _GEN_1733; // @[executor.scala 466:52]
  wire [7:0] _GEN_1896 = opcode_2 == 4'hf ? _GEN_1254 : _GEN_1734; // @[executor.scala 466:52]
  wire [7:0] _GEN_1897 = opcode_2 == 4'hf ? _GEN_1255 : _GEN_1735; // @[executor.scala 466:52]
  wire [7:0] _GEN_1898 = opcode_2 == 4'hf ? _GEN_1256 : _GEN_1736; // @[executor.scala 466:52]
  wire [7:0] _GEN_1899 = opcode_2 == 4'hf ? _GEN_1257 : _GEN_1737; // @[executor.scala 466:52]
  wire [7:0] _GEN_1900 = opcode_2 == 4'hf ? _GEN_1258 : _GEN_1738; // @[executor.scala 466:52]
  wire [7:0] _GEN_1901 = opcode_2 == 4'hf ? _GEN_1259 : _GEN_1739; // @[executor.scala 466:52]
  wire [7:0] _GEN_1902 = opcode_2 == 4'hf ? _GEN_1260 : _GEN_1740; // @[executor.scala 466:52]
  wire [7:0] _GEN_1903 = opcode_2 == 4'hf ? _GEN_1261 : _GEN_1741; // @[executor.scala 466:52]
  wire [7:0] _GEN_1904 = opcode_2 == 4'hf ? _GEN_1262 : _GEN_1742; // @[executor.scala 466:52]
  wire [7:0] _GEN_1905 = opcode_2 == 4'hf ? _GEN_1263 : _GEN_1743; // @[executor.scala 466:52]
  wire [7:0] _GEN_1906 = opcode_2 == 4'hf ? _GEN_1264 : _GEN_1744; // @[executor.scala 466:52]
  wire [7:0] _GEN_1907 = opcode_2 == 4'hf ? _GEN_1265 : _GEN_1745; // @[executor.scala 466:52]
  wire [7:0] _GEN_1908 = opcode_2 == 4'hf ? _GEN_1266 : _GEN_1746; // @[executor.scala 466:52]
  wire [7:0] _GEN_1909 = opcode_2 == 4'hf ? _GEN_1267 : _GEN_1747; // @[executor.scala 466:52]
  wire [7:0] _GEN_1910 = opcode_2 == 4'hf ? _GEN_1268 : _GEN_1748; // @[executor.scala 466:52]
  wire [7:0] _GEN_1911 = opcode_2 == 4'hf ? _GEN_1269 : _GEN_1749; // @[executor.scala 466:52]
  wire [7:0] _GEN_1912 = opcode_2 == 4'hf ? _GEN_1270 : _GEN_1750; // @[executor.scala 466:52]
  wire [7:0] _GEN_1913 = opcode_2 == 4'hf ? _GEN_1271 : _GEN_1751; // @[executor.scala 466:52]
  wire [7:0] _GEN_1914 = opcode_2 == 4'hf ? _GEN_1272 : _GEN_1752; // @[executor.scala 466:52]
  wire [7:0] _GEN_1915 = opcode_2 == 4'hf ? _GEN_1273 : _GEN_1753; // @[executor.scala 466:52]
  wire [7:0] _GEN_1916 = opcode_2 == 4'hf ? _GEN_1274 : _GEN_1754; // @[executor.scala 466:52]
  wire [7:0] _GEN_1917 = opcode_2 == 4'hf ? _GEN_1275 : _GEN_1755; // @[executor.scala 466:52]
  wire [7:0] _GEN_1918 = opcode_2 == 4'hf ? _GEN_1276 : _GEN_1756; // @[executor.scala 466:52]
  wire [7:0] _GEN_1919 = opcode_2 == 4'hf ? _GEN_1277 : _GEN_1757; // @[executor.scala 466:52]
  wire [7:0] _GEN_1920 = opcode_2 == 4'hf ? _GEN_1278 : _GEN_1758; // @[executor.scala 466:52]
  wire [7:0] _GEN_1921 = opcode_2 == 4'hf ? _GEN_1279 : _GEN_1759; // @[executor.scala 466:52]
  wire [7:0] _GEN_1922 = opcode_2 == 4'hf ? _GEN_1280 : _GEN_1760; // @[executor.scala 466:52]
  wire [7:0] _GEN_1923 = opcode_2 == 4'hf ? _GEN_1281 : _GEN_1761; // @[executor.scala 466:52]
  wire [7:0] _GEN_1924 = opcode_2 == 4'hf ? _GEN_1282 : _GEN_1762; // @[executor.scala 466:52]
  wire [7:0] _GEN_1925 = opcode_2 == 4'hf ? _GEN_1283 : _GEN_1763; // @[executor.scala 466:52]
  wire [3:0] opcode_3 = vliw_3[31:28]; // @[primitive.scala 9:44]
  wire [13:0] parameter_2_3 = vliw_3[13:0]; // @[primitive.scala 11:44]
  wire [7:0] _GEN_2850 = {{2'd0}, dst_offset_3}; // @[executor.scala 473:49]
  wire [7:0] byte_480 = field_3[7:0]; // @[executor.scala 475:56]
  wire [7:0] _GEN_1926 = mask_3[0] ? byte_480 : _GEN_1766; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] byte_481 = field_3[15:8]; // @[executor.scala 475:56]
  wire [7:0] _GEN_1927 = mask_3[1] ? byte_481 : _GEN_1767; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] byte_482 = field_3[23:16]; // @[executor.scala 475:56]
  wire [7:0] _GEN_1928 = mask_3[2] ? byte_482 : _GEN_1768; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] byte_483 = field_3[31:24]; // @[executor.scala 475:56]
  wire [7:0] _GEN_1929 = mask_3[3] ? byte_483 : _GEN_1769; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1930 = _GEN_2850 == 8'h0 ? _GEN_1926 : _GEN_1766; // @[executor.scala 473:84]
  wire [7:0] _GEN_1931 = _GEN_2850 == 8'h0 ? _GEN_1927 : _GEN_1767; // @[executor.scala 473:84]
  wire [7:0] _GEN_1932 = _GEN_2850 == 8'h0 ? _GEN_1928 : _GEN_1768; // @[executor.scala 473:84]
  wire [7:0] _GEN_1933 = _GEN_2850 == 8'h0 ? _GEN_1929 : _GEN_1769; // @[executor.scala 473:84]
  wire [7:0] _GEN_1934 = mask_3[0] ? byte_480 : _GEN_1770; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1935 = mask_3[1] ? byte_481 : _GEN_1771; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1936 = mask_3[2] ? byte_482 : _GEN_1772; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1937 = mask_3[3] ? byte_483 : _GEN_1773; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1938 = _GEN_2850 == 8'h1 ? _GEN_1934 : _GEN_1770; // @[executor.scala 473:84]
  wire [7:0] _GEN_1939 = _GEN_2850 == 8'h1 ? _GEN_1935 : _GEN_1771; // @[executor.scala 473:84]
  wire [7:0] _GEN_1940 = _GEN_2850 == 8'h1 ? _GEN_1936 : _GEN_1772; // @[executor.scala 473:84]
  wire [7:0] _GEN_1941 = _GEN_2850 == 8'h1 ? _GEN_1937 : _GEN_1773; // @[executor.scala 473:84]
  wire [7:0] _GEN_1942 = mask_3[0] ? byte_480 : _GEN_1774; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1943 = mask_3[1] ? byte_481 : _GEN_1775; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1944 = mask_3[2] ? byte_482 : _GEN_1776; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1945 = mask_3[3] ? byte_483 : _GEN_1777; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1946 = _GEN_2850 == 8'h2 ? _GEN_1942 : _GEN_1774; // @[executor.scala 473:84]
  wire [7:0] _GEN_1947 = _GEN_2850 == 8'h2 ? _GEN_1943 : _GEN_1775; // @[executor.scala 473:84]
  wire [7:0] _GEN_1948 = _GEN_2850 == 8'h2 ? _GEN_1944 : _GEN_1776; // @[executor.scala 473:84]
  wire [7:0] _GEN_1949 = _GEN_2850 == 8'h2 ? _GEN_1945 : _GEN_1777; // @[executor.scala 473:84]
  wire [7:0] _GEN_1950 = mask_3[0] ? byte_480 : _GEN_1778; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1951 = mask_3[1] ? byte_481 : _GEN_1779; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1952 = mask_3[2] ? byte_482 : _GEN_1780; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1953 = mask_3[3] ? byte_483 : _GEN_1781; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1954 = _GEN_2850 == 8'h3 ? _GEN_1950 : _GEN_1778; // @[executor.scala 473:84]
  wire [7:0] _GEN_1955 = _GEN_2850 == 8'h3 ? _GEN_1951 : _GEN_1779; // @[executor.scala 473:84]
  wire [7:0] _GEN_1956 = _GEN_2850 == 8'h3 ? _GEN_1952 : _GEN_1780; // @[executor.scala 473:84]
  wire [7:0] _GEN_1957 = _GEN_2850 == 8'h3 ? _GEN_1953 : _GEN_1781; // @[executor.scala 473:84]
  wire [7:0] _GEN_1958 = mask_3[0] ? byte_480 : _GEN_1782; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1959 = mask_3[1] ? byte_481 : _GEN_1783; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1960 = mask_3[2] ? byte_482 : _GEN_1784; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1961 = mask_3[3] ? byte_483 : _GEN_1785; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1962 = _GEN_2850 == 8'h4 ? _GEN_1958 : _GEN_1782; // @[executor.scala 473:84]
  wire [7:0] _GEN_1963 = _GEN_2850 == 8'h4 ? _GEN_1959 : _GEN_1783; // @[executor.scala 473:84]
  wire [7:0] _GEN_1964 = _GEN_2850 == 8'h4 ? _GEN_1960 : _GEN_1784; // @[executor.scala 473:84]
  wire [7:0] _GEN_1965 = _GEN_2850 == 8'h4 ? _GEN_1961 : _GEN_1785; // @[executor.scala 473:84]
  wire [7:0] _GEN_1966 = mask_3[0] ? byte_480 : _GEN_1786; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1967 = mask_3[1] ? byte_481 : _GEN_1787; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1968 = mask_3[2] ? byte_482 : _GEN_1788; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1969 = mask_3[3] ? byte_483 : _GEN_1789; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1970 = _GEN_2850 == 8'h5 ? _GEN_1966 : _GEN_1786; // @[executor.scala 473:84]
  wire [7:0] _GEN_1971 = _GEN_2850 == 8'h5 ? _GEN_1967 : _GEN_1787; // @[executor.scala 473:84]
  wire [7:0] _GEN_1972 = _GEN_2850 == 8'h5 ? _GEN_1968 : _GEN_1788; // @[executor.scala 473:84]
  wire [7:0] _GEN_1973 = _GEN_2850 == 8'h5 ? _GEN_1969 : _GEN_1789; // @[executor.scala 473:84]
  wire [7:0] _GEN_1974 = mask_3[0] ? byte_480 : _GEN_1790; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1975 = mask_3[1] ? byte_481 : _GEN_1791; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1976 = mask_3[2] ? byte_482 : _GEN_1792; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1977 = mask_3[3] ? byte_483 : _GEN_1793; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1978 = _GEN_2850 == 8'h6 ? _GEN_1974 : _GEN_1790; // @[executor.scala 473:84]
  wire [7:0] _GEN_1979 = _GEN_2850 == 8'h6 ? _GEN_1975 : _GEN_1791; // @[executor.scala 473:84]
  wire [7:0] _GEN_1980 = _GEN_2850 == 8'h6 ? _GEN_1976 : _GEN_1792; // @[executor.scala 473:84]
  wire [7:0] _GEN_1981 = _GEN_2850 == 8'h6 ? _GEN_1977 : _GEN_1793; // @[executor.scala 473:84]
  wire [7:0] _GEN_1982 = mask_3[0] ? byte_480 : _GEN_1794; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1983 = mask_3[1] ? byte_481 : _GEN_1795; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1984 = mask_3[2] ? byte_482 : _GEN_1796; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1985 = mask_3[3] ? byte_483 : _GEN_1797; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1986 = _GEN_2850 == 8'h7 ? _GEN_1982 : _GEN_1794; // @[executor.scala 473:84]
  wire [7:0] _GEN_1987 = _GEN_2850 == 8'h7 ? _GEN_1983 : _GEN_1795; // @[executor.scala 473:84]
  wire [7:0] _GEN_1988 = _GEN_2850 == 8'h7 ? _GEN_1984 : _GEN_1796; // @[executor.scala 473:84]
  wire [7:0] _GEN_1989 = _GEN_2850 == 8'h7 ? _GEN_1985 : _GEN_1797; // @[executor.scala 473:84]
  wire [7:0] _GEN_1990 = mask_3[0] ? byte_480 : _GEN_1798; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1991 = mask_3[1] ? byte_481 : _GEN_1799; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1992 = mask_3[2] ? byte_482 : _GEN_1800; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1993 = mask_3[3] ? byte_483 : _GEN_1801; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1994 = _GEN_2850 == 8'h8 ? _GEN_1990 : _GEN_1798; // @[executor.scala 473:84]
  wire [7:0] _GEN_1995 = _GEN_2850 == 8'h8 ? _GEN_1991 : _GEN_1799; // @[executor.scala 473:84]
  wire [7:0] _GEN_1996 = _GEN_2850 == 8'h8 ? _GEN_1992 : _GEN_1800; // @[executor.scala 473:84]
  wire [7:0] _GEN_1997 = _GEN_2850 == 8'h8 ? _GEN_1993 : _GEN_1801; // @[executor.scala 473:84]
  wire [7:0] _GEN_1998 = mask_3[0] ? byte_480 : _GEN_1802; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1999 = mask_3[1] ? byte_481 : _GEN_1803; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2000 = mask_3[2] ? byte_482 : _GEN_1804; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2001 = mask_3[3] ? byte_483 : _GEN_1805; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2002 = _GEN_2850 == 8'h9 ? _GEN_1998 : _GEN_1802; // @[executor.scala 473:84]
  wire [7:0] _GEN_2003 = _GEN_2850 == 8'h9 ? _GEN_1999 : _GEN_1803; // @[executor.scala 473:84]
  wire [7:0] _GEN_2004 = _GEN_2850 == 8'h9 ? _GEN_2000 : _GEN_1804; // @[executor.scala 473:84]
  wire [7:0] _GEN_2005 = _GEN_2850 == 8'h9 ? _GEN_2001 : _GEN_1805; // @[executor.scala 473:84]
  wire [7:0] _GEN_2006 = mask_3[0] ? byte_480 : _GEN_1806; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2007 = mask_3[1] ? byte_481 : _GEN_1807; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2008 = mask_3[2] ? byte_482 : _GEN_1808; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2009 = mask_3[3] ? byte_483 : _GEN_1809; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2010 = _GEN_2850 == 8'ha ? _GEN_2006 : _GEN_1806; // @[executor.scala 473:84]
  wire [7:0] _GEN_2011 = _GEN_2850 == 8'ha ? _GEN_2007 : _GEN_1807; // @[executor.scala 473:84]
  wire [7:0] _GEN_2012 = _GEN_2850 == 8'ha ? _GEN_2008 : _GEN_1808; // @[executor.scala 473:84]
  wire [7:0] _GEN_2013 = _GEN_2850 == 8'ha ? _GEN_2009 : _GEN_1809; // @[executor.scala 473:84]
  wire [7:0] _GEN_2014 = mask_3[0] ? byte_480 : _GEN_1810; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2015 = mask_3[1] ? byte_481 : _GEN_1811; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2016 = mask_3[2] ? byte_482 : _GEN_1812; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2017 = mask_3[3] ? byte_483 : _GEN_1813; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2018 = _GEN_2850 == 8'hb ? _GEN_2014 : _GEN_1810; // @[executor.scala 473:84]
  wire [7:0] _GEN_2019 = _GEN_2850 == 8'hb ? _GEN_2015 : _GEN_1811; // @[executor.scala 473:84]
  wire [7:0] _GEN_2020 = _GEN_2850 == 8'hb ? _GEN_2016 : _GEN_1812; // @[executor.scala 473:84]
  wire [7:0] _GEN_2021 = _GEN_2850 == 8'hb ? _GEN_2017 : _GEN_1813; // @[executor.scala 473:84]
  wire [7:0] _GEN_2022 = mask_3[0] ? byte_480 : _GEN_1814; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2023 = mask_3[1] ? byte_481 : _GEN_1815; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2024 = mask_3[2] ? byte_482 : _GEN_1816; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2025 = mask_3[3] ? byte_483 : _GEN_1817; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2026 = _GEN_2850 == 8'hc ? _GEN_2022 : _GEN_1814; // @[executor.scala 473:84]
  wire [7:0] _GEN_2027 = _GEN_2850 == 8'hc ? _GEN_2023 : _GEN_1815; // @[executor.scala 473:84]
  wire [7:0] _GEN_2028 = _GEN_2850 == 8'hc ? _GEN_2024 : _GEN_1816; // @[executor.scala 473:84]
  wire [7:0] _GEN_2029 = _GEN_2850 == 8'hc ? _GEN_2025 : _GEN_1817; // @[executor.scala 473:84]
  wire [7:0] _GEN_2030 = mask_3[0] ? byte_480 : _GEN_1818; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2031 = mask_3[1] ? byte_481 : _GEN_1819; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2032 = mask_3[2] ? byte_482 : _GEN_1820; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2033 = mask_3[3] ? byte_483 : _GEN_1821; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2034 = _GEN_2850 == 8'hd ? _GEN_2030 : _GEN_1818; // @[executor.scala 473:84]
  wire [7:0] _GEN_2035 = _GEN_2850 == 8'hd ? _GEN_2031 : _GEN_1819; // @[executor.scala 473:84]
  wire [7:0] _GEN_2036 = _GEN_2850 == 8'hd ? _GEN_2032 : _GEN_1820; // @[executor.scala 473:84]
  wire [7:0] _GEN_2037 = _GEN_2850 == 8'hd ? _GEN_2033 : _GEN_1821; // @[executor.scala 473:84]
  wire [7:0] _GEN_2038 = mask_3[0] ? byte_480 : _GEN_1822; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2039 = mask_3[1] ? byte_481 : _GEN_1823; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2040 = mask_3[2] ? byte_482 : _GEN_1824; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2041 = mask_3[3] ? byte_483 : _GEN_1825; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2042 = _GEN_2850 == 8'he ? _GEN_2038 : _GEN_1822; // @[executor.scala 473:84]
  wire [7:0] _GEN_2043 = _GEN_2850 == 8'he ? _GEN_2039 : _GEN_1823; // @[executor.scala 473:84]
  wire [7:0] _GEN_2044 = _GEN_2850 == 8'he ? _GEN_2040 : _GEN_1824; // @[executor.scala 473:84]
  wire [7:0] _GEN_2045 = _GEN_2850 == 8'he ? _GEN_2041 : _GEN_1825; // @[executor.scala 473:84]
  wire [7:0] _GEN_2046 = mask_3[0] ? byte_480 : _GEN_1826; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2047 = mask_3[1] ? byte_481 : _GEN_1827; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2048 = mask_3[2] ? byte_482 : _GEN_1828; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2049 = mask_3[3] ? byte_483 : _GEN_1829; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2050 = _GEN_2850 == 8'hf ? _GEN_2046 : _GEN_1826; // @[executor.scala 473:84]
  wire [7:0] _GEN_2051 = _GEN_2850 == 8'hf ? _GEN_2047 : _GEN_1827; // @[executor.scala 473:84]
  wire [7:0] _GEN_2052 = _GEN_2850 == 8'hf ? _GEN_2048 : _GEN_1828; // @[executor.scala 473:84]
  wire [7:0] _GEN_2053 = _GEN_2850 == 8'hf ? _GEN_2049 : _GEN_1829; // @[executor.scala 473:84]
  wire [7:0] _GEN_2054 = mask_3[0] ? byte_480 : _GEN_1830; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2055 = mask_3[1] ? byte_481 : _GEN_1831; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2056 = mask_3[2] ? byte_482 : _GEN_1832; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2057 = mask_3[3] ? byte_483 : _GEN_1833; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2058 = _GEN_2850 == 8'h10 ? _GEN_2054 : _GEN_1830; // @[executor.scala 473:84]
  wire [7:0] _GEN_2059 = _GEN_2850 == 8'h10 ? _GEN_2055 : _GEN_1831; // @[executor.scala 473:84]
  wire [7:0] _GEN_2060 = _GEN_2850 == 8'h10 ? _GEN_2056 : _GEN_1832; // @[executor.scala 473:84]
  wire [7:0] _GEN_2061 = _GEN_2850 == 8'h10 ? _GEN_2057 : _GEN_1833; // @[executor.scala 473:84]
  wire [7:0] _GEN_2062 = mask_3[0] ? byte_480 : _GEN_1834; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2063 = mask_3[1] ? byte_481 : _GEN_1835; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2064 = mask_3[2] ? byte_482 : _GEN_1836; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2065 = mask_3[3] ? byte_483 : _GEN_1837; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2066 = _GEN_2850 == 8'h11 ? _GEN_2062 : _GEN_1834; // @[executor.scala 473:84]
  wire [7:0] _GEN_2067 = _GEN_2850 == 8'h11 ? _GEN_2063 : _GEN_1835; // @[executor.scala 473:84]
  wire [7:0] _GEN_2068 = _GEN_2850 == 8'h11 ? _GEN_2064 : _GEN_1836; // @[executor.scala 473:84]
  wire [7:0] _GEN_2069 = _GEN_2850 == 8'h11 ? _GEN_2065 : _GEN_1837; // @[executor.scala 473:84]
  wire [7:0] _GEN_2070 = mask_3[0] ? byte_480 : _GEN_1838; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2071 = mask_3[1] ? byte_481 : _GEN_1839; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2072 = mask_3[2] ? byte_482 : _GEN_1840; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2073 = mask_3[3] ? byte_483 : _GEN_1841; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2074 = _GEN_2850 == 8'h12 ? _GEN_2070 : _GEN_1838; // @[executor.scala 473:84]
  wire [7:0] _GEN_2075 = _GEN_2850 == 8'h12 ? _GEN_2071 : _GEN_1839; // @[executor.scala 473:84]
  wire [7:0] _GEN_2076 = _GEN_2850 == 8'h12 ? _GEN_2072 : _GEN_1840; // @[executor.scala 473:84]
  wire [7:0] _GEN_2077 = _GEN_2850 == 8'h12 ? _GEN_2073 : _GEN_1841; // @[executor.scala 473:84]
  wire [7:0] _GEN_2078 = mask_3[0] ? byte_480 : _GEN_1842; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2079 = mask_3[1] ? byte_481 : _GEN_1843; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2080 = mask_3[2] ? byte_482 : _GEN_1844; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2081 = mask_3[3] ? byte_483 : _GEN_1845; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2082 = _GEN_2850 == 8'h13 ? _GEN_2078 : _GEN_1842; // @[executor.scala 473:84]
  wire [7:0] _GEN_2083 = _GEN_2850 == 8'h13 ? _GEN_2079 : _GEN_1843; // @[executor.scala 473:84]
  wire [7:0] _GEN_2084 = _GEN_2850 == 8'h13 ? _GEN_2080 : _GEN_1844; // @[executor.scala 473:84]
  wire [7:0] _GEN_2085 = _GEN_2850 == 8'h13 ? _GEN_2081 : _GEN_1845; // @[executor.scala 473:84]
  wire [7:0] _GEN_2086 = mask_3[0] ? byte_480 : _GEN_1846; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2087 = mask_3[1] ? byte_481 : _GEN_1847; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2088 = mask_3[2] ? byte_482 : _GEN_1848; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2089 = mask_3[3] ? byte_483 : _GEN_1849; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2090 = _GEN_2850 == 8'h14 ? _GEN_2086 : _GEN_1846; // @[executor.scala 473:84]
  wire [7:0] _GEN_2091 = _GEN_2850 == 8'h14 ? _GEN_2087 : _GEN_1847; // @[executor.scala 473:84]
  wire [7:0] _GEN_2092 = _GEN_2850 == 8'h14 ? _GEN_2088 : _GEN_1848; // @[executor.scala 473:84]
  wire [7:0] _GEN_2093 = _GEN_2850 == 8'h14 ? _GEN_2089 : _GEN_1849; // @[executor.scala 473:84]
  wire [7:0] _GEN_2094 = mask_3[0] ? byte_480 : _GEN_1850; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2095 = mask_3[1] ? byte_481 : _GEN_1851; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2096 = mask_3[2] ? byte_482 : _GEN_1852; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2097 = mask_3[3] ? byte_483 : _GEN_1853; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2098 = _GEN_2850 == 8'h15 ? _GEN_2094 : _GEN_1850; // @[executor.scala 473:84]
  wire [7:0] _GEN_2099 = _GEN_2850 == 8'h15 ? _GEN_2095 : _GEN_1851; // @[executor.scala 473:84]
  wire [7:0] _GEN_2100 = _GEN_2850 == 8'h15 ? _GEN_2096 : _GEN_1852; // @[executor.scala 473:84]
  wire [7:0] _GEN_2101 = _GEN_2850 == 8'h15 ? _GEN_2097 : _GEN_1853; // @[executor.scala 473:84]
  wire [7:0] _GEN_2102 = mask_3[0] ? byte_480 : _GEN_1854; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2103 = mask_3[1] ? byte_481 : _GEN_1855; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2104 = mask_3[2] ? byte_482 : _GEN_1856; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2105 = mask_3[3] ? byte_483 : _GEN_1857; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2106 = _GEN_2850 == 8'h16 ? _GEN_2102 : _GEN_1854; // @[executor.scala 473:84]
  wire [7:0] _GEN_2107 = _GEN_2850 == 8'h16 ? _GEN_2103 : _GEN_1855; // @[executor.scala 473:84]
  wire [7:0] _GEN_2108 = _GEN_2850 == 8'h16 ? _GEN_2104 : _GEN_1856; // @[executor.scala 473:84]
  wire [7:0] _GEN_2109 = _GEN_2850 == 8'h16 ? _GEN_2105 : _GEN_1857; // @[executor.scala 473:84]
  wire [7:0] _GEN_2110 = mask_3[0] ? byte_480 : _GEN_1858; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2111 = mask_3[1] ? byte_481 : _GEN_1859; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2112 = mask_3[2] ? byte_482 : _GEN_1860; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2113 = mask_3[3] ? byte_483 : _GEN_1861; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2114 = _GEN_2850 == 8'h17 ? _GEN_2110 : _GEN_1858; // @[executor.scala 473:84]
  wire [7:0] _GEN_2115 = _GEN_2850 == 8'h17 ? _GEN_2111 : _GEN_1859; // @[executor.scala 473:84]
  wire [7:0] _GEN_2116 = _GEN_2850 == 8'h17 ? _GEN_2112 : _GEN_1860; // @[executor.scala 473:84]
  wire [7:0] _GEN_2117 = _GEN_2850 == 8'h17 ? _GEN_2113 : _GEN_1861; // @[executor.scala 473:84]
  wire [7:0] _GEN_2118 = mask_3[0] ? byte_480 : _GEN_1862; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2119 = mask_3[1] ? byte_481 : _GEN_1863; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2120 = mask_3[2] ? byte_482 : _GEN_1864; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2121 = mask_3[3] ? byte_483 : _GEN_1865; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2122 = _GEN_2850 == 8'h18 ? _GEN_2118 : _GEN_1862; // @[executor.scala 473:84]
  wire [7:0] _GEN_2123 = _GEN_2850 == 8'h18 ? _GEN_2119 : _GEN_1863; // @[executor.scala 473:84]
  wire [7:0] _GEN_2124 = _GEN_2850 == 8'h18 ? _GEN_2120 : _GEN_1864; // @[executor.scala 473:84]
  wire [7:0] _GEN_2125 = _GEN_2850 == 8'h18 ? _GEN_2121 : _GEN_1865; // @[executor.scala 473:84]
  wire [7:0] _GEN_2126 = mask_3[0] ? byte_480 : _GEN_1866; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2127 = mask_3[1] ? byte_481 : _GEN_1867; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2128 = mask_3[2] ? byte_482 : _GEN_1868; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2129 = mask_3[3] ? byte_483 : _GEN_1869; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2130 = _GEN_2850 == 8'h19 ? _GEN_2126 : _GEN_1866; // @[executor.scala 473:84]
  wire [7:0] _GEN_2131 = _GEN_2850 == 8'h19 ? _GEN_2127 : _GEN_1867; // @[executor.scala 473:84]
  wire [7:0] _GEN_2132 = _GEN_2850 == 8'h19 ? _GEN_2128 : _GEN_1868; // @[executor.scala 473:84]
  wire [7:0] _GEN_2133 = _GEN_2850 == 8'h19 ? _GEN_2129 : _GEN_1869; // @[executor.scala 473:84]
  wire [7:0] _GEN_2134 = mask_3[0] ? byte_480 : _GEN_1870; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2135 = mask_3[1] ? byte_481 : _GEN_1871; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2136 = mask_3[2] ? byte_482 : _GEN_1872; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2137 = mask_3[3] ? byte_483 : _GEN_1873; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2138 = _GEN_2850 == 8'h1a ? _GEN_2134 : _GEN_1870; // @[executor.scala 473:84]
  wire [7:0] _GEN_2139 = _GEN_2850 == 8'h1a ? _GEN_2135 : _GEN_1871; // @[executor.scala 473:84]
  wire [7:0] _GEN_2140 = _GEN_2850 == 8'h1a ? _GEN_2136 : _GEN_1872; // @[executor.scala 473:84]
  wire [7:0] _GEN_2141 = _GEN_2850 == 8'h1a ? _GEN_2137 : _GEN_1873; // @[executor.scala 473:84]
  wire [7:0] _GEN_2142 = mask_3[0] ? byte_480 : _GEN_1874; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2143 = mask_3[1] ? byte_481 : _GEN_1875; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2144 = mask_3[2] ? byte_482 : _GEN_1876; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2145 = mask_3[3] ? byte_483 : _GEN_1877; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2146 = _GEN_2850 == 8'h1b ? _GEN_2142 : _GEN_1874; // @[executor.scala 473:84]
  wire [7:0] _GEN_2147 = _GEN_2850 == 8'h1b ? _GEN_2143 : _GEN_1875; // @[executor.scala 473:84]
  wire [7:0] _GEN_2148 = _GEN_2850 == 8'h1b ? _GEN_2144 : _GEN_1876; // @[executor.scala 473:84]
  wire [7:0] _GEN_2149 = _GEN_2850 == 8'h1b ? _GEN_2145 : _GEN_1877; // @[executor.scala 473:84]
  wire [7:0] _GEN_2150 = mask_3[0] ? byte_480 : _GEN_1878; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2151 = mask_3[1] ? byte_481 : _GEN_1879; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2152 = mask_3[2] ? byte_482 : _GEN_1880; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2153 = mask_3[3] ? byte_483 : _GEN_1881; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2154 = _GEN_2850 == 8'h1c ? _GEN_2150 : _GEN_1878; // @[executor.scala 473:84]
  wire [7:0] _GEN_2155 = _GEN_2850 == 8'h1c ? _GEN_2151 : _GEN_1879; // @[executor.scala 473:84]
  wire [7:0] _GEN_2156 = _GEN_2850 == 8'h1c ? _GEN_2152 : _GEN_1880; // @[executor.scala 473:84]
  wire [7:0] _GEN_2157 = _GEN_2850 == 8'h1c ? _GEN_2153 : _GEN_1881; // @[executor.scala 473:84]
  wire [7:0] _GEN_2158 = mask_3[0] ? byte_480 : _GEN_1882; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2159 = mask_3[1] ? byte_481 : _GEN_1883; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2160 = mask_3[2] ? byte_482 : _GEN_1884; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2161 = mask_3[3] ? byte_483 : _GEN_1885; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2162 = _GEN_2850 == 8'h1d ? _GEN_2158 : _GEN_1882; // @[executor.scala 473:84]
  wire [7:0] _GEN_2163 = _GEN_2850 == 8'h1d ? _GEN_2159 : _GEN_1883; // @[executor.scala 473:84]
  wire [7:0] _GEN_2164 = _GEN_2850 == 8'h1d ? _GEN_2160 : _GEN_1884; // @[executor.scala 473:84]
  wire [7:0] _GEN_2165 = _GEN_2850 == 8'h1d ? _GEN_2161 : _GEN_1885; // @[executor.scala 473:84]
  wire [7:0] _GEN_2166 = mask_3[0] ? byte_480 : _GEN_1886; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2167 = mask_3[1] ? byte_481 : _GEN_1887; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2168 = mask_3[2] ? byte_482 : _GEN_1888; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2169 = mask_3[3] ? byte_483 : _GEN_1889; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2170 = _GEN_2850 == 8'h1e ? _GEN_2166 : _GEN_1886; // @[executor.scala 473:84]
  wire [7:0] _GEN_2171 = _GEN_2850 == 8'h1e ? _GEN_2167 : _GEN_1887; // @[executor.scala 473:84]
  wire [7:0] _GEN_2172 = _GEN_2850 == 8'h1e ? _GEN_2168 : _GEN_1888; // @[executor.scala 473:84]
  wire [7:0] _GEN_2173 = _GEN_2850 == 8'h1e ? _GEN_2169 : _GEN_1889; // @[executor.scala 473:84]
  wire [7:0] _GEN_2174 = mask_3[0] ? byte_480 : _GEN_1890; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2175 = mask_3[1] ? byte_481 : _GEN_1891; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2176 = mask_3[2] ? byte_482 : _GEN_1892; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2177 = mask_3[3] ? byte_483 : _GEN_1893; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2178 = _GEN_2850 == 8'h1f ? _GEN_2174 : _GEN_1890; // @[executor.scala 473:84]
  wire [7:0] _GEN_2179 = _GEN_2850 == 8'h1f ? _GEN_2175 : _GEN_1891; // @[executor.scala 473:84]
  wire [7:0] _GEN_2180 = _GEN_2850 == 8'h1f ? _GEN_2176 : _GEN_1892; // @[executor.scala 473:84]
  wire [7:0] _GEN_2181 = _GEN_2850 == 8'h1f ? _GEN_2177 : _GEN_1893; // @[executor.scala 473:84]
  wire [7:0] _GEN_2182 = mask_3[0] ? byte_480 : _GEN_1894; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2183 = mask_3[1] ? byte_481 : _GEN_1895; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2184 = mask_3[2] ? byte_482 : _GEN_1896; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2185 = mask_3[3] ? byte_483 : _GEN_1897; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2186 = _GEN_2850 == 8'h20 ? _GEN_2182 : _GEN_1894; // @[executor.scala 473:84]
  wire [7:0] _GEN_2187 = _GEN_2850 == 8'h20 ? _GEN_2183 : _GEN_1895; // @[executor.scala 473:84]
  wire [7:0] _GEN_2188 = _GEN_2850 == 8'h20 ? _GEN_2184 : _GEN_1896; // @[executor.scala 473:84]
  wire [7:0] _GEN_2189 = _GEN_2850 == 8'h20 ? _GEN_2185 : _GEN_1897; // @[executor.scala 473:84]
  wire [7:0] _GEN_2190 = mask_3[0] ? byte_480 : _GEN_1898; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2191 = mask_3[1] ? byte_481 : _GEN_1899; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2192 = mask_3[2] ? byte_482 : _GEN_1900; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2193 = mask_3[3] ? byte_483 : _GEN_1901; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2194 = _GEN_2850 == 8'h21 ? _GEN_2190 : _GEN_1898; // @[executor.scala 473:84]
  wire [7:0] _GEN_2195 = _GEN_2850 == 8'h21 ? _GEN_2191 : _GEN_1899; // @[executor.scala 473:84]
  wire [7:0] _GEN_2196 = _GEN_2850 == 8'h21 ? _GEN_2192 : _GEN_1900; // @[executor.scala 473:84]
  wire [7:0] _GEN_2197 = _GEN_2850 == 8'h21 ? _GEN_2193 : _GEN_1901; // @[executor.scala 473:84]
  wire [7:0] _GEN_2198 = mask_3[0] ? byte_480 : _GEN_1902; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2199 = mask_3[1] ? byte_481 : _GEN_1903; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2200 = mask_3[2] ? byte_482 : _GEN_1904; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2201 = mask_3[3] ? byte_483 : _GEN_1905; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2202 = _GEN_2850 == 8'h22 ? _GEN_2198 : _GEN_1902; // @[executor.scala 473:84]
  wire [7:0] _GEN_2203 = _GEN_2850 == 8'h22 ? _GEN_2199 : _GEN_1903; // @[executor.scala 473:84]
  wire [7:0] _GEN_2204 = _GEN_2850 == 8'h22 ? _GEN_2200 : _GEN_1904; // @[executor.scala 473:84]
  wire [7:0] _GEN_2205 = _GEN_2850 == 8'h22 ? _GEN_2201 : _GEN_1905; // @[executor.scala 473:84]
  wire [7:0] _GEN_2206 = mask_3[0] ? byte_480 : _GEN_1906; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2207 = mask_3[1] ? byte_481 : _GEN_1907; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2208 = mask_3[2] ? byte_482 : _GEN_1908; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2209 = mask_3[3] ? byte_483 : _GEN_1909; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2210 = _GEN_2850 == 8'h23 ? _GEN_2206 : _GEN_1906; // @[executor.scala 473:84]
  wire [7:0] _GEN_2211 = _GEN_2850 == 8'h23 ? _GEN_2207 : _GEN_1907; // @[executor.scala 473:84]
  wire [7:0] _GEN_2212 = _GEN_2850 == 8'h23 ? _GEN_2208 : _GEN_1908; // @[executor.scala 473:84]
  wire [7:0] _GEN_2213 = _GEN_2850 == 8'h23 ? _GEN_2209 : _GEN_1909; // @[executor.scala 473:84]
  wire [7:0] _GEN_2214 = mask_3[0] ? byte_480 : _GEN_1910; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2215 = mask_3[1] ? byte_481 : _GEN_1911; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2216 = mask_3[2] ? byte_482 : _GEN_1912; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2217 = mask_3[3] ? byte_483 : _GEN_1913; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2218 = _GEN_2850 == 8'h24 ? _GEN_2214 : _GEN_1910; // @[executor.scala 473:84]
  wire [7:0] _GEN_2219 = _GEN_2850 == 8'h24 ? _GEN_2215 : _GEN_1911; // @[executor.scala 473:84]
  wire [7:0] _GEN_2220 = _GEN_2850 == 8'h24 ? _GEN_2216 : _GEN_1912; // @[executor.scala 473:84]
  wire [7:0] _GEN_2221 = _GEN_2850 == 8'h24 ? _GEN_2217 : _GEN_1913; // @[executor.scala 473:84]
  wire [7:0] _GEN_2222 = mask_3[0] ? byte_480 : _GEN_1914; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2223 = mask_3[1] ? byte_481 : _GEN_1915; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2224 = mask_3[2] ? byte_482 : _GEN_1916; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2225 = mask_3[3] ? byte_483 : _GEN_1917; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2226 = _GEN_2850 == 8'h25 ? _GEN_2222 : _GEN_1914; // @[executor.scala 473:84]
  wire [7:0] _GEN_2227 = _GEN_2850 == 8'h25 ? _GEN_2223 : _GEN_1915; // @[executor.scala 473:84]
  wire [7:0] _GEN_2228 = _GEN_2850 == 8'h25 ? _GEN_2224 : _GEN_1916; // @[executor.scala 473:84]
  wire [7:0] _GEN_2229 = _GEN_2850 == 8'h25 ? _GEN_2225 : _GEN_1917; // @[executor.scala 473:84]
  wire [7:0] _GEN_2230 = mask_3[0] ? byte_480 : _GEN_1918; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2231 = mask_3[1] ? byte_481 : _GEN_1919; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2232 = mask_3[2] ? byte_482 : _GEN_1920; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2233 = mask_3[3] ? byte_483 : _GEN_1921; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2234 = _GEN_2850 == 8'h26 ? _GEN_2230 : _GEN_1918; // @[executor.scala 473:84]
  wire [7:0] _GEN_2235 = _GEN_2850 == 8'h26 ? _GEN_2231 : _GEN_1919; // @[executor.scala 473:84]
  wire [7:0] _GEN_2236 = _GEN_2850 == 8'h26 ? _GEN_2232 : _GEN_1920; // @[executor.scala 473:84]
  wire [7:0] _GEN_2237 = _GEN_2850 == 8'h26 ? _GEN_2233 : _GEN_1921; // @[executor.scala 473:84]
  wire [7:0] _GEN_2238 = mask_3[0] ? byte_480 : _GEN_1922; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2239 = mask_3[1] ? byte_481 : _GEN_1923; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2240 = mask_3[2] ? byte_482 : _GEN_1924; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2241 = mask_3[3] ? byte_483 : _GEN_1925; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2242 = _GEN_2850 == 8'h27 ? _GEN_2238 : _GEN_1922; // @[executor.scala 473:84]
  wire [7:0] _GEN_2243 = _GEN_2850 == 8'h27 ? _GEN_2239 : _GEN_1923; // @[executor.scala 473:84]
  wire [7:0] _GEN_2244 = _GEN_2850 == 8'h27 ? _GEN_2240 : _GEN_1924; // @[executor.scala 473:84]
  wire [7:0] _GEN_2245 = _GEN_2850 == 8'h27 ? _GEN_2241 : _GEN_1925; // @[executor.scala 473:84]
  wire [7:0] _GEN_2246 = opcode_3 != 4'h0 ? _GEN_1930 : _GEN_1766; // @[executor.scala 470:55]
  wire [7:0] _GEN_2247 = opcode_3 != 4'h0 ? _GEN_1931 : _GEN_1767; // @[executor.scala 470:55]
  wire [7:0] _GEN_2248 = opcode_3 != 4'h0 ? _GEN_1932 : _GEN_1768; // @[executor.scala 470:55]
  wire [7:0] _GEN_2249 = opcode_3 != 4'h0 ? _GEN_1933 : _GEN_1769; // @[executor.scala 470:55]
  wire [7:0] _GEN_2250 = opcode_3 != 4'h0 ? _GEN_1938 : _GEN_1770; // @[executor.scala 470:55]
  wire [7:0] _GEN_2251 = opcode_3 != 4'h0 ? _GEN_1939 : _GEN_1771; // @[executor.scala 470:55]
  wire [7:0] _GEN_2252 = opcode_3 != 4'h0 ? _GEN_1940 : _GEN_1772; // @[executor.scala 470:55]
  wire [7:0] _GEN_2253 = opcode_3 != 4'h0 ? _GEN_1941 : _GEN_1773; // @[executor.scala 470:55]
  wire [7:0] _GEN_2254 = opcode_3 != 4'h0 ? _GEN_1946 : _GEN_1774; // @[executor.scala 470:55]
  wire [7:0] _GEN_2255 = opcode_3 != 4'h0 ? _GEN_1947 : _GEN_1775; // @[executor.scala 470:55]
  wire [7:0] _GEN_2256 = opcode_3 != 4'h0 ? _GEN_1948 : _GEN_1776; // @[executor.scala 470:55]
  wire [7:0] _GEN_2257 = opcode_3 != 4'h0 ? _GEN_1949 : _GEN_1777; // @[executor.scala 470:55]
  wire [7:0] _GEN_2258 = opcode_3 != 4'h0 ? _GEN_1954 : _GEN_1778; // @[executor.scala 470:55]
  wire [7:0] _GEN_2259 = opcode_3 != 4'h0 ? _GEN_1955 : _GEN_1779; // @[executor.scala 470:55]
  wire [7:0] _GEN_2260 = opcode_3 != 4'h0 ? _GEN_1956 : _GEN_1780; // @[executor.scala 470:55]
  wire [7:0] _GEN_2261 = opcode_3 != 4'h0 ? _GEN_1957 : _GEN_1781; // @[executor.scala 470:55]
  wire [7:0] _GEN_2262 = opcode_3 != 4'h0 ? _GEN_1962 : _GEN_1782; // @[executor.scala 470:55]
  wire [7:0] _GEN_2263 = opcode_3 != 4'h0 ? _GEN_1963 : _GEN_1783; // @[executor.scala 470:55]
  wire [7:0] _GEN_2264 = opcode_3 != 4'h0 ? _GEN_1964 : _GEN_1784; // @[executor.scala 470:55]
  wire [7:0] _GEN_2265 = opcode_3 != 4'h0 ? _GEN_1965 : _GEN_1785; // @[executor.scala 470:55]
  wire [7:0] _GEN_2266 = opcode_3 != 4'h0 ? _GEN_1970 : _GEN_1786; // @[executor.scala 470:55]
  wire [7:0] _GEN_2267 = opcode_3 != 4'h0 ? _GEN_1971 : _GEN_1787; // @[executor.scala 470:55]
  wire [7:0] _GEN_2268 = opcode_3 != 4'h0 ? _GEN_1972 : _GEN_1788; // @[executor.scala 470:55]
  wire [7:0] _GEN_2269 = opcode_3 != 4'h0 ? _GEN_1973 : _GEN_1789; // @[executor.scala 470:55]
  wire [7:0] _GEN_2270 = opcode_3 != 4'h0 ? _GEN_1978 : _GEN_1790; // @[executor.scala 470:55]
  wire [7:0] _GEN_2271 = opcode_3 != 4'h0 ? _GEN_1979 : _GEN_1791; // @[executor.scala 470:55]
  wire [7:0] _GEN_2272 = opcode_3 != 4'h0 ? _GEN_1980 : _GEN_1792; // @[executor.scala 470:55]
  wire [7:0] _GEN_2273 = opcode_3 != 4'h0 ? _GEN_1981 : _GEN_1793; // @[executor.scala 470:55]
  wire [7:0] _GEN_2274 = opcode_3 != 4'h0 ? _GEN_1986 : _GEN_1794; // @[executor.scala 470:55]
  wire [7:0] _GEN_2275 = opcode_3 != 4'h0 ? _GEN_1987 : _GEN_1795; // @[executor.scala 470:55]
  wire [7:0] _GEN_2276 = opcode_3 != 4'h0 ? _GEN_1988 : _GEN_1796; // @[executor.scala 470:55]
  wire [7:0] _GEN_2277 = opcode_3 != 4'h0 ? _GEN_1989 : _GEN_1797; // @[executor.scala 470:55]
  wire [7:0] _GEN_2278 = opcode_3 != 4'h0 ? _GEN_1994 : _GEN_1798; // @[executor.scala 470:55]
  wire [7:0] _GEN_2279 = opcode_3 != 4'h0 ? _GEN_1995 : _GEN_1799; // @[executor.scala 470:55]
  wire [7:0] _GEN_2280 = opcode_3 != 4'h0 ? _GEN_1996 : _GEN_1800; // @[executor.scala 470:55]
  wire [7:0] _GEN_2281 = opcode_3 != 4'h0 ? _GEN_1997 : _GEN_1801; // @[executor.scala 470:55]
  wire [7:0] _GEN_2282 = opcode_3 != 4'h0 ? _GEN_2002 : _GEN_1802; // @[executor.scala 470:55]
  wire [7:0] _GEN_2283 = opcode_3 != 4'h0 ? _GEN_2003 : _GEN_1803; // @[executor.scala 470:55]
  wire [7:0] _GEN_2284 = opcode_3 != 4'h0 ? _GEN_2004 : _GEN_1804; // @[executor.scala 470:55]
  wire [7:0] _GEN_2285 = opcode_3 != 4'h0 ? _GEN_2005 : _GEN_1805; // @[executor.scala 470:55]
  wire [7:0] _GEN_2286 = opcode_3 != 4'h0 ? _GEN_2010 : _GEN_1806; // @[executor.scala 470:55]
  wire [7:0] _GEN_2287 = opcode_3 != 4'h0 ? _GEN_2011 : _GEN_1807; // @[executor.scala 470:55]
  wire [7:0] _GEN_2288 = opcode_3 != 4'h0 ? _GEN_2012 : _GEN_1808; // @[executor.scala 470:55]
  wire [7:0] _GEN_2289 = opcode_3 != 4'h0 ? _GEN_2013 : _GEN_1809; // @[executor.scala 470:55]
  wire [7:0] _GEN_2290 = opcode_3 != 4'h0 ? _GEN_2018 : _GEN_1810; // @[executor.scala 470:55]
  wire [7:0] _GEN_2291 = opcode_3 != 4'h0 ? _GEN_2019 : _GEN_1811; // @[executor.scala 470:55]
  wire [7:0] _GEN_2292 = opcode_3 != 4'h0 ? _GEN_2020 : _GEN_1812; // @[executor.scala 470:55]
  wire [7:0] _GEN_2293 = opcode_3 != 4'h0 ? _GEN_2021 : _GEN_1813; // @[executor.scala 470:55]
  wire [7:0] _GEN_2294 = opcode_3 != 4'h0 ? _GEN_2026 : _GEN_1814; // @[executor.scala 470:55]
  wire [7:0] _GEN_2295 = opcode_3 != 4'h0 ? _GEN_2027 : _GEN_1815; // @[executor.scala 470:55]
  wire [7:0] _GEN_2296 = opcode_3 != 4'h0 ? _GEN_2028 : _GEN_1816; // @[executor.scala 470:55]
  wire [7:0] _GEN_2297 = opcode_3 != 4'h0 ? _GEN_2029 : _GEN_1817; // @[executor.scala 470:55]
  wire [7:0] _GEN_2298 = opcode_3 != 4'h0 ? _GEN_2034 : _GEN_1818; // @[executor.scala 470:55]
  wire [7:0] _GEN_2299 = opcode_3 != 4'h0 ? _GEN_2035 : _GEN_1819; // @[executor.scala 470:55]
  wire [7:0] _GEN_2300 = opcode_3 != 4'h0 ? _GEN_2036 : _GEN_1820; // @[executor.scala 470:55]
  wire [7:0] _GEN_2301 = opcode_3 != 4'h0 ? _GEN_2037 : _GEN_1821; // @[executor.scala 470:55]
  wire [7:0] _GEN_2302 = opcode_3 != 4'h0 ? _GEN_2042 : _GEN_1822; // @[executor.scala 470:55]
  wire [7:0] _GEN_2303 = opcode_3 != 4'h0 ? _GEN_2043 : _GEN_1823; // @[executor.scala 470:55]
  wire [7:0] _GEN_2304 = opcode_3 != 4'h0 ? _GEN_2044 : _GEN_1824; // @[executor.scala 470:55]
  wire [7:0] _GEN_2305 = opcode_3 != 4'h0 ? _GEN_2045 : _GEN_1825; // @[executor.scala 470:55]
  wire [7:0] _GEN_2306 = opcode_3 != 4'h0 ? _GEN_2050 : _GEN_1826; // @[executor.scala 470:55]
  wire [7:0] _GEN_2307 = opcode_3 != 4'h0 ? _GEN_2051 : _GEN_1827; // @[executor.scala 470:55]
  wire [7:0] _GEN_2308 = opcode_3 != 4'h0 ? _GEN_2052 : _GEN_1828; // @[executor.scala 470:55]
  wire [7:0] _GEN_2309 = opcode_3 != 4'h0 ? _GEN_2053 : _GEN_1829; // @[executor.scala 470:55]
  wire [7:0] _GEN_2310 = opcode_3 != 4'h0 ? _GEN_2058 : _GEN_1830; // @[executor.scala 470:55]
  wire [7:0] _GEN_2311 = opcode_3 != 4'h0 ? _GEN_2059 : _GEN_1831; // @[executor.scala 470:55]
  wire [7:0] _GEN_2312 = opcode_3 != 4'h0 ? _GEN_2060 : _GEN_1832; // @[executor.scala 470:55]
  wire [7:0] _GEN_2313 = opcode_3 != 4'h0 ? _GEN_2061 : _GEN_1833; // @[executor.scala 470:55]
  wire [7:0] _GEN_2314 = opcode_3 != 4'h0 ? _GEN_2066 : _GEN_1834; // @[executor.scala 470:55]
  wire [7:0] _GEN_2315 = opcode_3 != 4'h0 ? _GEN_2067 : _GEN_1835; // @[executor.scala 470:55]
  wire [7:0] _GEN_2316 = opcode_3 != 4'h0 ? _GEN_2068 : _GEN_1836; // @[executor.scala 470:55]
  wire [7:0] _GEN_2317 = opcode_3 != 4'h0 ? _GEN_2069 : _GEN_1837; // @[executor.scala 470:55]
  wire [7:0] _GEN_2318 = opcode_3 != 4'h0 ? _GEN_2074 : _GEN_1838; // @[executor.scala 470:55]
  wire [7:0] _GEN_2319 = opcode_3 != 4'h0 ? _GEN_2075 : _GEN_1839; // @[executor.scala 470:55]
  wire [7:0] _GEN_2320 = opcode_3 != 4'h0 ? _GEN_2076 : _GEN_1840; // @[executor.scala 470:55]
  wire [7:0] _GEN_2321 = opcode_3 != 4'h0 ? _GEN_2077 : _GEN_1841; // @[executor.scala 470:55]
  wire [7:0] _GEN_2322 = opcode_3 != 4'h0 ? _GEN_2082 : _GEN_1842; // @[executor.scala 470:55]
  wire [7:0] _GEN_2323 = opcode_3 != 4'h0 ? _GEN_2083 : _GEN_1843; // @[executor.scala 470:55]
  wire [7:0] _GEN_2324 = opcode_3 != 4'h0 ? _GEN_2084 : _GEN_1844; // @[executor.scala 470:55]
  wire [7:0] _GEN_2325 = opcode_3 != 4'h0 ? _GEN_2085 : _GEN_1845; // @[executor.scala 470:55]
  wire [7:0] _GEN_2326 = opcode_3 != 4'h0 ? _GEN_2090 : _GEN_1846; // @[executor.scala 470:55]
  wire [7:0] _GEN_2327 = opcode_3 != 4'h0 ? _GEN_2091 : _GEN_1847; // @[executor.scala 470:55]
  wire [7:0] _GEN_2328 = opcode_3 != 4'h0 ? _GEN_2092 : _GEN_1848; // @[executor.scala 470:55]
  wire [7:0] _GEN_2329 = opcode_3 != 4'h0 ? _GEN_2093 : _GEN_1849; // @[executor.scala 470:55]
  wire [7:0] _GEN_2330 = opcode_3 != 4'h0 ? _GEN_2098 : _GEN_1850; // @[executor.scala 470:55]
  wire [7:0] _GEN_2331 = opcode_3 != 4'h0 ? _GEN_2099 : _GEN_1851; // @[executor.scala 470:55]
  wire [7:0] _GEN_2332 = opcode_3 != 4'h0 ? _GEN_2100 : _GEN_1852; // @[executor.scala 470:55]
  wire [7:0] _GEN_2333 = opcode_3 != 4'h0 ? _GEN_2101 : _GEN_1853; // @[executor.scala 470:55]
  wire [7:0] _GEN_2334 = opcode_3 != 4'h0 ? _GEN_2106 : _GEN_1854; // @[executor.scala 470:55]
  wire [7:0] _GEN_2335 = opcode_3 != 4'h0 ? _GEN_2107 : _GEN_1855; // @[executor.scala 470:55]
  wire [7:0] _GEN_2336 = opcode_3 != 4'h0 ? _GEN_2108 : _GEN_1856; // @[executor.scala 470:55]
  wire [7:0] _GEN_2337 = opcode_3 != 4'h0 ? _GEN_2109 : _GEN_1857; // @[executor.scala 470:55]
  wire [7:0] _GEN_2338 = opcode_3 != 4'h0 ? _GEN_2114 : _GEN_1858; // @[executor.scala 470:55]
  wire [7:0] _GEN_2339 = opcode_3 != 4'h0 ? _GEN_2115 : _GEN_1859; // @[executor.scala 470:55]
  wire [7:0] _GEN_2340 = opcode_3 != 4'h0 ? _GEN_2116 : _GEN_1860; // @[executor.scala 470:55]
  wire [7:0] _GEN_2341 = opcode_3 != 4'h0 ? _GEN_2117 : _GEN_1861; // @[executor.scala 470:55]
  wire [7:0] _GEN_2342 = opcode_3 != 4'h0 ? _GEN_2122 : _GEN_1862; // @[executor.scala 470:55]
  wire [7:0] _GEN_2343 = opcode_3 != 4'h0 ? _GEN_2123 : _GEN_1863; // @[executor.scala 470:55]
  wire [7:0] _GEN_2344 = opcode_3 != 4'h0 ? _GEN_2124 : _GEN_1864; // @[executor.scala 470:55]
  wire [7:0] _GEN_2345 = opcode_3 != 4'h0 ? _GEN_2125 : _GEN_1865; // @[executor.scala 470:55]
  wire [7:0] _GEN_2346 = opcode_3 != 4'h0 ? _GEN_2130 : _GEN_1866; // @[executor.scala 470:55]
  wire [7:0] _GEN_2347 = opcode_3 != 4'h0 ? _GEN_2131 : _GEN_1867; // @[executor.scala 470:55]
  wire [7:0] _GEN_2348 = opcode_3 != 4'h0 ? _GEN_2132 : _GEN_1868; // @[executor.scala 470:55]
  wire [7:0] _GEN_2349 = opcode_3 != 4'h0 ? _GEN_2133 : _GEN_1869; // @[executor.scala 470:55]
  wire [7:0] _GEN_2350 = opcode_3 != 4'h0 ? _GEN_2138 : _GEN_1870; // @[executor.scala 470:55]
  wire [7:0] _GEN_2351 = opcode_3 != 4'h0 ? _GEN_2139 : _GEN_1871; // @[executor.scala 470:55]
  wire [7:0] _GEN_2352 = opcode_3 != 4'h0 ? _GEN_2140 : _GEN_1872; // @[executor.scala 470:55]
  wire [7:0] _GEN_2353 = opcode_3 != 4'h0 ? _GEN_2141 : _GEN_1873; // @[executor.scala 470:55]
  wire [7:0] _GEN_2354 = opcode_3 != 4'h0 ? _GEN_2146 : _GEN_1874; // @[executor.scala 470:55]
  wire [7:0] _GEN_2355 = opcode_3 != 4'h0 ? _GEN_2147 : _GEN_1875; // @[executor.scala 470:55]
  wire [7:0] _GEN_2356 = opcode_3 != 4'h0 ? _GEN_2148 : _GEN_1876; // @[executor.scala 470:55]
  wire [7:0] _GEN_2357 = opcode_3 != 4'h0 ? _GEN_2149 : _GEN_1877; // @[executor.scala 470:55]
  wire [7:0] _GEN_2358 = opcode_3 != 4'h0 ? _GEN_2154 : _GEN_1878; // @[executor.scala 470:55]
  wire [7:0] _GEN_2359 = opcode_3 != 4'h0 ? _GEN_2155 : _GEN_1879; // @[executor.scala 470:55]
  wire [7:0] _GEN_2360 = opcode_3 != 4'h0 ? _GEN_2156 : _GEN_1880; // @[executor.scala 470:55]
  wire [7:0] _GEN_2361 = opcode_3 != 4'h0 ? _GEN_2157 : _GEN_1881; // @[executor.scala 470:55]
  wire [7:0] _GEN_2362 = opcode_3 != 4'h0 ? _GEN_2162 : _GEN_1882; // @[executor.scala 470:55]
  wire [7:0] _GEN_2363 = opcode_3 != 4'h0 ? _GEN_2163 : _GEN_1883; // @[executor.scala 470:55]
  wire [7:0] _GEN_2364 = opcode_3 != 4'h0 ? _GEN_2164 : _GEN_1884; // @[executor.scala 470:55]
  wire [7:0] _GEN_2365 = opcode_3 != 4'h0 ? _GEN_2165 : _GEN_1885; // @[executor.scala 470:55]
  wire [7:0] _GEN_2366 = opcode_3 != 4'h0 ? _GEN_2170 : _GEN_1886; // @[executor.scala 470:55]
  wire [7:0] _GEN_2367 = opcode_3 != 4'h0 ? _GEN_2171 : _GEN_1887; // @[executor.scala 470:55]
  wire [7:0] _GEN_2368 = opcode_3 != 4'h0 ? _GEN_2172 : _GEN_1888; // @[executor.scala 470:55]
  wire [7:0] _GEN_2369 = opcode_3 != 4'h0 ? _GEN_2173 : _GEN_1889; // @[executor.scala 470:55]
  wire [7:0] _GEN_2370 = opcode_3 != 4'h0 ? _GEN_2178 : _GEN_1890; // @[executor.scala 470:55]
  wire [7:0] _GEN_2371 = opcode_3 != 4'h0 ? _GEN_2179 : _GEN_1891; // @[executor.scala 470:55]
  wire [7:0] _GEN_2372 = opcode_3 != 4'h0 ? _GEN_2180 : _GEN_1892; // @[executor.scala 470:55]
  wire [7:0] _GEN_2373 = opcode_3 != 4'h0 ? _GEN_2181 : _GEN_1893; // @[executor.scala 470:55]
  wire [7:0] _GEN_2374 = opcode_3 != 4'h0 ? _GEN_2186 : _GEN_1894; // @[executor.scala 470:55]
  wire [7:0] _GEN_2375 = opcode_3 != 4'h0 ? _GEN_2187 : _GEN_1895; // @[executor.scala 470:55]
  wire [7:0] _GEN_2376 = opcode_3 != 4'h0 ? _GEN_2188 : _GEN_1896; // @[executor.scala 470:55]
  wire [7:0] _GEN_2377 = opcode_3 != 4'h0 ? _GEN_2189 : _GEN_1897; // @[executor.scala 470:55]
  wire [7:0] _GEN_2378 = opcode_3 != 4'h0 ? _GEN_2194 : _GEN_1898; // @[executor.scala 470:55]
  wire [7:0] _GEN_2379 = opcode_3 != 4'h0 ? _GEN_2195 : _GEN_1899; // @[executor.scala 470:55]
  wire [7:0] _GEN_2380 = opcode_3 != 4'h0 ? _GEN_2196 : _GEN_1900; // @[executor.scala 470:55]
  wire [7:0] _GEN_2381 = opcode_3 != 4'h0 ? _GEN_2197 : _GEN_1901; // @[executor.scala 470:55]
  wire [7:0] _GEN_2382 = opcode_3 != 4'h0 ? _GEN_2202 : _GEN_1902; // @[executor.scala 470:55]
  wire [7:0] _GEN_2383 = opcode_3 != 4'h0 ? _GEN_2203 : _GEN_1903; // @[executor.scala 470:55]
  wire [7:0] _GEN_2384 = opcode_3 != 4'h0 ? _GEN_2204 : _GEN_1904; // @[executor.scala 470:55]
  wire [7:0] _GEN_2385 = opcode_3 != 4'h0 ? _GEN_2205 : _GEN_1905; // @[executor.scala 470:55]
  wire [7:0] _GEN_2386 = opcode_3 != 4'h0 ? _GEN_2210 : _GEN_1906; // @[executor.scala 470:55]
  wire [7:0] _GEN_2387 = opcode_3 != 4'h0 ? _GEN_2211 : _GEN_1907; // @[executor.scala 470:55]
  wire [7:0] _GEN_2388 = opcode_3 != 4'h0 ? _GEN_2212 : _GEN_1908; // @[executor.scala 470:55]
  wire [7:0] _GEN_2389 = opcode_3 != 4'h0 ? _GEN_2213 : _GEN_1909; // @[executor.scala 470:55]
  wire [7:0] _GEN_2390 = opcode_3 != 4'h0 ? _GEN_2218 : _GEN_1910; // @[executor.scala 470:55]
  wire [7:0] _GEN_2391 = opcode_3 != 4'h0 ? _GEN_2219 : _GEN_1911; // @[executor.scala 470:55]
  wire [7:0] _GEN_2392 = opcode_3 != 4'h0 ? _GEN_2220 : _GEN_1912; // @[executor.scala 470:55]
  wire [7:0] _GEN_2393 = opcode_3 != 4'h0 ? _GEN_2221 : _GEN_1913; // @[executor.scala 470:55]
  wire [7:0] _GEN_2394 = opcode_3 != 4'h0 ? _GEN_2226 : _GEN_1914; // @[executor.scala 470:55]
  wire [7:0] _GEN_2395 = opcode_3 != 4'h0 ? _GEN_2227 : _GEN_1915; // @[executor.scala 470:55]
  wire [7:0] _GEN_2396 = opcode_3 != 4'h0 ? _GEN_2228 : _GEN_1916; // @[executor.scala 470:55]
  wire [7:0] _GEN_2397 = opcode_3 != 4'h0 ? _GEN_2229 : _GEN_1917; // @[executor.scala 470:55]
  wire [7:0] _GEN_2398 = opcode_3 != 4'h0 ? _GEN_2234 : _GEN_1918; // @[executor.scala 470:55]
  wire [7:0] _GEN_2399 = opcode_3 != 4'h0 ? _GEN_2235 : _GEN_1919; // @[executor.scala 470:55]
  wire [7:0] _GEN_2400 = opcode_3 != 4'h0 ? _GEN_2236 : _GEN_1920; // @[executor.scala 470:55]
  wire [7:0] _GEN_2401 = opcode_3 != 4'h0 ? _GEN_2237 : _GEN_1921; // @[executor.scala 470:55]
  wire [7:0] _GEN_2402 = opcode_3 != 4'h0 ? _GEN_2242 : _GEN_1922; // @[executor.scala 470:55]
  wire [7:0] _GEN_2403 = opcode_3 != 4'h0 ? _GEN_2243 : _GEN_1923; // @[executor.scala 470:55]
  wire [7:0] _GEN_2404 = opcode_3 != 4'h0 ? _GEN_2244 : _GEN_1924; // @[executor.scala 470:55]
  wire [7:0] _GEN_2405 = opcode_3 != 4'h0 ? _GEN_2245 : _GEN_1925; // @[executor.scala 470:55]
  wire [3:0] _GEN_2406 = opcode_3 == 4'hf ? parameter_2_3[13:10] : _GEN_1764; // @[executor.scala 466:52 executor.scala 467:55]
  wire  _GEN_2407 = opcode_3 == 4'hf ? parameter_2_3[0] : _GEN_1765; // @[executor.scala 466:52 executor.scala 468:55]
  wire [7:0] _GEN_2408 = opcode_3 == 4'hf ? _GEN_1766 : _GEN_2246; // @[executor.scala 466:52]
  wire [7:0] _GEN_2409 = opcode_3 == 4'hf ? _GEN_1767 : _GEN_2247; // @[executor.scala 466:52]
  wire [7:0] _GEN_2410 = opcode_3 == 4'hf ? _GEN_1768 : _GEN_2248; // @[executor.scala 466:52]
  wire [7:0] _GEN_2411 = opcode_3 == 4'hf ? _GEN_1769 : _GEN_2249; // @[executor.scala 466:52]
  wire [7:0] _GEN_2412 = opcode_3 == 4'hf ? _GEN_1770 : _GEN_2250; // @[executor.scala 466:52]
  wire [7:0] _GEN_2413 = opcode_3 == 4'hf ? _GEN_1771 : _GEN_2251; // @[executor.scala 466:52]
  wire [7:0] _GEN_2414 = opcode_3 == 4'hf ? _GEN_1772 : _GEN_2252; // @[executor.scala 466:52]
  wire [7:0] _GEN_2415 = opcode_3 == 4'hf ? _GEN_1773 : _GEN_2253; // @[executor.scala 466:52]
  wire [7:0] _GEN_2416 = opcode_3 == 4'hf ? _GEN_1774 : _GEN_2254; // @[executor.scala 466:52]
  wire [7:0] _GEN_2417 = opcode_3 == 4'hf ? _GEN_1775 : _GEN_2255; // @[executor.scala 466:52]
  wire [7:0] _GEN_2418 = opcode_3 == 4'hf ? _GEN_1776 : _GEN_2256; // @[executor.scala 466:52]
  wire [7:0] _GEN_2419 = opcode_3 == 4'hf ? _GEN_1777 : _GEN_2257; // @[executor.scala 466:52]
  wire [7:0] _GEN_2420 = opcode_3 == 4'hf ? _GEN_1778 : _GEN_2258; // @[executor.scala 466:52]
  wire [7:0] _GEN_2421 = opcode_3 == 4'hf ? _GEN_1779 : _GEN_2259; // @[executor.scala 466:52]
  wire [7:0] _GEN_2422 = opcode_3 == 4'hf ? _GEN_1780 : _GEN_2260; // @[executor.scala 466:52]
  wire [7:0] _GEN_2423 = opcode_3 == 4'hf ? _GEN_1781 : _GEN_2261; // @[executor.scala 466:52]
  wire [7:0] _GEN_2424 = opcode_3 == 4'hf ? _GEN_1782 : _GEN_2262; // @[executor.scala 466:52]
  wire [7:0] _GEN_2425 = opcode_3 == 4'hf ? _GEN_1783 : _GEN_2263; // @[executor.scala 466:52]
  wire [7:0] _GEN_2426 = opcode_3 == 4'hf ? _GEN_1784 : _GEN_2264; // @[executor.scala 466:52]
  wire [7:0] _GEN_2427 = opcode_3 == 4'hf ? _GEN_1785 : _GEN_2265; // @[executor.scala 466:52]
  wire [7:0] _GEN_2428 = opcode_3 == 4'hf ? _GEN_1786 : _GEN_2266; // @[executor.scala 466:52]
  wire [7:0] _GEN_2429 = opcode_3 == 4'hf ? _GEN_1787 : _GEN_2267; // @[executor.scala 466:52]
  wire [7:0] _GEN_2430 = opcode_3 == 4'hf ? _GEN_1788 : _GEN_2268; // @[executor.scala 466:52]
  wire [7:0] _GEN_2431 = opcode_3 == 4'hf ? _GEN_1789 : _GEN_2269; // @[executor.scala 466:52]
  wire [7:0] _GEN_2432 = opcode_3 == 4'hf ? _GEN_1790 : _GEN_2270; // @[executor.scala 466:52]
  wire [7:0] _GEN_2433 = opcode_3 == 4'hf ? _GEN_1791 : _GEN_2271; // @[executor.scala 466:52]
  wire [7:0] _GEN_2434 = opcode_3 == 4'hf ? _GEN_1792 : _GEN_2272; // @[executor.scala 466:52]
  wire [7:0] _GEN_2435 = opcode_3 == 4'hf ? _GEN_1793 : _GEN_2273; // @[executor.scala 466:52]
  wire [7:0] _GEN_2436 = opcode_3 == 4'hf ? _GEN_1794 : _GEN_2274; // @[executor.scala 466:52]
  wire [7:0] _GEN_2437 = opcode_3 == 4'hf ? _GEN_1795 : _GEN_2275; // @[executor.scala 466:52]
  wire [7:0] _GEN_2438 = opcode_3 == 4'hf ? _GEN_1796 : _GEN_2276; // @[executor.scala 466:52]
  wire [7:0] _GEN_2439 = opcode_3 == 4'hf ? _GEN_1797 : _GEN_2277; // @[executor.scala 466:52]
  wire [7:0] _GEN_2440 = opcode_3 == 4'hf ? _GEN_1798 : _GEN_2278; // @[executor.scala 466:52]
  wire [7:0] _GEN_2441 = opcode_3 == 4'hf ? _GEN_1799 : _GEN_2279; // @[executor.scala 466:52]
  wire [7:0] _GEN_2442 = opcode_3 == 4'hf ? _GEN_1800 : _GEN_2280; // @[executor.scala 466:52]
  wire [7:0] _GEN_2443 = opcode_3 == 4'hf ? _GEN_1801 : _GEN_2281; // @[executor.scala 466:52]
  wire [7:0] _GEN_2444 = opcode_3 == 4'hf ? _GEN_1802 : _GEN_2282; // @[executor.scala 466:52]
  wire [7:0] _GEN_2445 = opcode_3 == 4'hf ? _GEN_1803 : _GEN_2283; // @[executor.scala 466:52]
  wire [7:0] _GEN_2446 = opcode_3 == 4'hf ? _GEN_1804 : _GEN_2284; // @[executor.scala 466:52]
  wire [7:0] _GEN_2447 = opcode_3 == 4'hf ? _GEN_1805 : _GEN_2285; // @[executor.scala 466:52]
  wire [7:0] _GEN_2448 = opcode_3 == 4'hf ? _GEN_1806 : _GEN_2286; // @[executor.scala 466:52]
  wire [7:0] _GEN_2449 = opcode_3 == 4'hf ? _GEN_1807 : _GEN_2287; // @[executor.scala 466:52]
  wire [7:0] _GEN_2450 = opcode_3 == 4'hf ? _GEN_1808 : _GEN_2288; // @[executor.scala 466:52]
  wire [7:0] _GEN_2451 = opcode_3 == 4'hf ? _GEN_1809 : _GEN_2289; // @[executor.scala 466:52]
  wire [7:0] _GEN_2452 = opcode_3 == 4'hf ? _GEN_1810 : _GEN_2290; // @[executor.scala 466:52]
  wire [7:0] _GEN_2453 = opcode_3 == 4'hf ? _GEN_1811 : _GEN_2291; // @[executor.scala 466:52]
  wire [7:0] _GEN_2454 = opcode_3 == 4'hf ? _GEN_1812 : _GEN_2292; // @[executor.scala 466:52]
  wire [7:0] _GEN_2455 = opcode_3 == 4'hf ? _GEN_1813 : _GEN_2293; // @[executor.scala 466:52]
  wire [7:0] _GEN_2456 = opcode_3 == 4'hf ? _GEN_1814 : _GEN_2294; // @[executor.scala 466:52]
  wire [7:0] _GEN_2457 = opcode_3 == 4'hf ? _GEN_1815 : _GEN_2295; // @[executor.scala 466:52]
  wire [7:0] _GEN_2458 = opcode_3 == 4'hf ? _GEN_1816 : _GEN_2296; // @[executor.scala 466:52]
  wire [7:0] _GEN_2459 = opcode_3 == 4'hf ? _GEN_1817 : _GEN_2297; // @[executor.scala 466:52]
  wire [7:0] _GEN_2460 = opcode_3 == 4'hf ? _GEN_1818 : _GEN_2298; // @[executor.scala 466:52]
  wire [7:0] _GEN_2461 = opcode_3 == 4'hf ? _GEN_1819 : _GEN_2299; // @[executor.scala 466:52]
  wire [7:0] _GEN_2462 = opcode_3 == 4'hf ? _GEN_1820 : _GEN_2300; // @[executor.scala 466:52]
  wire [7:0] _GEN_2463 = opcode_3 == 4'hf ? _GEN_1821 : _GEN_2301; // @[executor.scala 466:52]
  wire [7:0] _GEN_2464 = opcode_3 == 4'hf ? _GEN_1822 : _GEN_2302; // @[executor.scala 466:52]
  wire [7:0] _GEN_2465 = opcode_3 == 4'hf ? _GEN_1823 : _GEN_2303; // @[executor.scala 466:52]
  wire [7:0] _GEN_2466 = opcode_3 == 4'hf ? _GEN_1824 : _GEN_2304; // @[executor.scala 466:52]
  wire [7:0] _GEN_2467 = opcode_3 == 4'hf ? _GEN_1825 : _GEN_2305; // @[executor.scala 466:52]
  wire [7:0] _GEN_2468 = opcode_3 == 4'hf ? _GEN_1826 : _GEN_2306; // @[executor.scala 466:52]
  wire [7:0] _GEN_2469 = opcode_3 == 4'hf ? _GEN_1827 : _GEN_2307; // @[executor.scala 466:52]
  wire [7:0] _GEN_2470 = opcode_3 == 4'hf ? _GEN_1828 : _GEN_2308; // @[executor.scala 466:52]
  wire [7:0] _GEN_2471 = opcode_3 == 4'hf ? _GEN_1829 : _GEN_2309; // @[executor.scala 466:52]
  wire [7:0] _GEN_2472 = opcode_3 == 4'hf ? _GEN_1830 : _GEN_2310; // @[executor.scala 466:52]
  wire [7:0] _GEN_2473 = opcode_3 == 4'hf ? _GEN_1831 : _GEN_2311; // @[executor.scala 466:52]
  wire [7:0] _GEN_2474 = opcode_3 == 4'hf ? _GEN_1832 : _GEN_2312; // @[executor.scala 466:52]
  wire [7:0] _GEN_2475 = opcode_3 == 4'hf ? _GEN_1833 : _GEN_2313; // @[executor.scala 466:52]
  wire [7:0] _GEN_2476 = opcode_3 == 4'hf ? _GEN_1834 : _GEN_2314; // @[executor.scala 466:52]
  wire [7:0] _GEN_2477 = opcode_3 == 4'hf ? _GEN_1835 : _GEN_2315; // @[executor.scala 466:52]
  wire [7:0] _GEN_2478 = opcode_3 == 4'hf ? _GEN_1836 : _GEN_2316; // @[executor.scala 466:52]
  wire [7:0] _GEN_2479 = opcode_3 == 4'hf ? _GEN_1837 : _GEN_2317; // @[executor.scala 466:52]
  wire [7:0] _GEN_2480 = opcode_3 == 4'hf ? _GEN_1838 : _GEN_2318; // @[executor.scala 466:52]
  wire [7:0] _GEN_2481 = opcode_3 == 4'hf ? _GEN_1839 : _GEN_2319; // @[executor.scala 466:52]
  wire [7:0] _GEN_2482 = opcode_3 == 4'hf ? _GEN_1840 : _GEN_2320; // @[executor.scala 466:52]
  wire [7:0] _GEN_2483 = opcode_3 == 4'hf ? _GEN_1841 : _GEN_2321; // @[executor.scala 466:52]
  wire [7:0] _GEN_2484 = opcode_3 == 4'hf ? _GEN_1842 : _GEN_2322; // @[executor.scala 466:52]
  wire [7:0] _GEN_2485 = opcode_3 == 4'hf ? _GEN_1843 : _GEN_2323; // @[executor.scala 466:52]
  wire [7:0] _GEN_2486 = opcode_3 == 4'hf ? _GEN_1844 : _GEN_2324; // @[executor.scala 466:52]
  wire [7:0] _GEN_2487 = opcode_3 == 4'hf ? _GEN_1845 : _GEN_2325; // @[executor.scala 466:52]
  wire [7:0] _GEN_2488 = opcode_3 == 4'hf ? _GEN_1846 : _GEN_2326; // @[executor.scala 466:52]
  wire [7:0] _GEN_2489 = opcode_3 == 4'hf ? _GEN_1847 : _GEN_2327; // @[executor.scala 466:52]
  wire [7:0] _GEN_2490 = opcode_3 == 4'hf ? _GEN_1848 : _GEN_2328; // @[executor.scala 466:52]
  wire [7:0] _GEN_2491 = opcode_3 == 4'hf ? _GEN_1849 : _GEN_2329; // @[executor.scala 466:52]
  wire [7:0] _GEN_2492 = opcode_3 == 4'hf ? _GEN_1850 : _GEN_2330; // @[executor.scala 466:52]
  wire [7:0] _GEN_2493 = opcode_3 == 4'hf ? _GEN_1851 : _GEN_2331; // @[executor.scala 466:52]
  wire [7:0] _GEN_2494 = opcode_3 == 4'hf ? _GEN_1852 : _GEN_2332; // @[executor.scala 466:52]
  wire [7:0] _GEN_2495 = opcode_3 == 4'hf ? _GEN_1853 : _GEN_2333; // @[executor.scala 466:52]
  wire [7:0] _GEN_2496 = opcode_3 == 4'hf ? _GEN_1854 : _GEN_2334; // @[executor.scala 466:52]
  wire [7:0] _GEN_2497 = opcode_3 == 4'hf ? _GEN_1855 : _GEN_2335; // @[executor.scala 466:52]
  wire [7:0] _GEN_2498 = opcode_3 == 4'hf ? _GEN_1856 : _GEN_2336; // @[executor.scala 466:52]
  wire [7:0] _GEN_2499 = opcode_3 == 4'hf ? _GEN_1857 : _GEN_2337; // @[executor.scala 466:52]
  wire [7:0] _GEN_2500 = opcode_3 == 4'hf ? _GEN_1858 : _GEN_2338; // @[executor.scala 466:52]
  wire [7:0] _GEN_2501 = opcode_3 == 4'hf ? _GEN_1859 : _GEN_2339; // @[executor.scala 466:52]
  wire [7:0] _GEN_2502 = opcode_3 == 4'hf ? _GEN_1860 : _GEN_2340; // @[executor.scala 466:52]
  wire [7:0] _GEN_2503 = opcode_3 == 4'hf ? _GEN_1861 : _GEN_2341; // @[executor.scala 466:52]
  wire [7:0] _GEN_2504 = opcode_3 == 4'hf ? _GEN_1862 : _GEN_2342; // @[executor.scala 466:52]
  wire [7:0] _GEN_2505 = opcode_3 == 4'hf ? _GEN_1863 : _GEN_2343; // @[executor.scala 466:52]
  wire [7:0] _GEN_2506 = opcode_3 == 4'hf ? _GEN_1864 : _GEN_2344; // @[executor.scala 466:52]
  wire [7:0] _GEN_2507 = opcode_3 == 4'hf ? _GEN_1865 : _GEN_2345; // @[executor.scala 466:52]
  wire [7:0] _GEN_2508 = opcode_3 == 4'hf ? _GEN_1866 : _GEN_2346; // @[executor.scala 466:52]
  wire [7:0] _GEN_2509 = opcode_3 == 4'hf ? _GEN_1867 : _GEN_2347; // @[executor.scala 466:52]
  wire [7:0] _GEN_2510 = opcode_3 == 4'hf ? _GEN_1868 : _GEN_2348; // @[executor.scala 466:52]
  wire [7:0] _GEN_2511 = opcode_3 == 4'hf ? _GEN_1869 : _GEN_2349; // @[executor.scala 466:52]
  wire [7:0] _GEN_2512 = opcode_3 == 4'hf ? _GEN_1870 : _GEN_2350; // @[executor.scala 466:52]
  wire [7:0] _GEN_2513 = opcode_3 == 4'hf ? _GEN_1871 : _GEN_2351; // @[executor.scala 466:52]
  wire [7:0] _GEN_2514 = opcode_3 == 4'hf ? _GEN_1872 : _GEN_2352; // @[executor.scala 466:52]
  wire [7:0] _GEN_2515 = opcode_3 == 4'hf ? _GEN_1873 : _GEN_2353; // @[executor.scala 466:52]
  wire [7:0] _GEN_2516 = opcode_3 == 4'hf ? _GEN_1874 : _GEN_2354; // @[executor.scala 466:52]
  wire [7:0] _GEN_2517 = opcode_3 == 4'hf ? _GEN_1875 : _GEN_2355; // @[executor.scala 466:52]
  wire [7:0] _GEN_2518 = opcode_3 == 4'hf ? _GEN_1876 : _GEN_2356; // @[executor.scala 466:52]
  wire [7:0] _GEN_2519 = opcode_3 == 4'hf ? _GEN_1877 : _GEN_2357; // @[executor.scala 466:52]
  wire [7:0] _GEN_2520 = opcode_3 == 4'hf ? _GEN_1878 : _GEN_2358; // @[executor.scala 466:52]
  wire [7:0] _GEN_2521 = opcode_3 == 4'hf ? _GEN_1879 : _GEN_2359; // @[executor.scala 466:52]
  wire [7:0] _GEN_2522 = opcode_3 == 4'hf ? _GEN_1880 : _GEN_2360; // @[executor.scala 466:52]
  wire [7:0] _GEN_2523 = opcode_3 == 4'hf ? _GEN_1881 : _GEN_2361; // @[executor.scala 466:52]
  wire [7:0] _GEN_2524 = opcode_3 == 4'hf ? _GEN_1882 : _GEN_2362; // @[executor.scala 466:52]
  wire [7:0] _GEN_2525 = opcode_3 == 4'hf ? _GEN_1883 : _GEN_2363; // @[executor.scala 466:52]
  wire [7:0] _GEN_2526 = opcode_3 == 4'hf ? _GEN_1884 : _GEN_2364; // @[executor.scala 466:52]
  wire [7:0] _GEN_2527 = opcode_3 == 4'hf ? _GEN_1885 : _GEN_2365; // @[executor.scala 466:52]
  wire [7:0] _GEN_2528 = opcode_3 == 4'hf ? _GEN_1886 : _GEN_2366; // @[executor.scala 466:52]
  wire [7:0] _GEN_2529 = opcode_3 == 4'hf ? _GEN_1887 : _GEN_2367; // @[executor.scala 466:52]
  wire [7:0] _GEN_2530 = opcode_3 == 4'hf ? _GEN_1888 : _GEN_2368; // @[executor.scala 466:52]
  wire [7:0] _GEN_2531 = opcode_3 == 4'hf ? _GEN_1889 : _GEN_2369; // @[executor.scala 466:52]
  wire [7:0] _GEN_2532 = opcode_3 == 4'hf ? _GEN_1890 : _GEN_2370; // @[executor.scala 466:52]
  wire [7:0] _GEN_2533 = opcode_3 == 4'hf ? _GEN_1891 : _GEN_2371; // @[executor.scala 466:52]
  wire [7:0] _GEN_2534 = opcode_3 == 4'hf ? _GEN_1892 : _GEN_2372; // @[executor.scala 466:52]
  wire [7:0] _GEN_2535 = opcode_3 == 4'hf ? _GEN_1893 : _GEN_2373; // @[executor.scala 466:52]
  wire [7:0] _GEN_2536 = opcode_3 == 4'hf ? _GEN_1894 : _GEN_2374; // @[executor.scala 466:52]
  wire [7:0] _GEN_2537 = opcode_3 == 4'hf ? _GEN_1895 : _GEN_2375; // @[executor.scala 466:52]
  wire [7:0] _GEN_2538 = opcode_3 == 4'hf ? _GEN_1896 : _GEN_2376; // @[executor.scala 466:52]
  wire [7:0] _GEN_2539 = opcode_3 == 4'hf ? _GEN_1897 : _GEN_2377; // @[executor.scala 466:52]
  wire [7:0] _GEN_2540 = opcode_3 == 4'hf ? _GEN_1898 : _GEN_2378; // @[executor.scala 466:52]
  wire [7:0] _GEN_2541 = opcode_3 == 4'hf ? _GEN_1899 : _GEN_2379; // @[executor.scala 466:52]
  wire [7:0] _GEN_2542 = opcode_3 == 4'hf ? _GEN_1900 : _GEN_2380; // @[executor.scala 466:52]
  wire [7:0] _GEN_2543 = opcode_3 == 4'hf ? _GEN_1901 : _GEN_2381; // @[executor.scala 466:52]
  wire [7:0] _GEN_2544 = opcode_3 == 4'hf ? _GEN_1902 : _GEN_2382; // @[executor.scala 466:52]
  wire [7:0] _GEN_2545 = opcode_3 == 4'hf ? _GEN_1903 : _GEN_2383; // @[executor.scala 466:52]
  wire [7:0] _GEN_2546 = opcode_3 == 4'hf ? _GEN_1904 : _GEN_2384; // @[executor.scala 466:52]
  wire [7:0] _GEN_2547 = opcode_3 == 4'hf ? _GEN_1905 : _GEN_2385; // @[executor.scala 466:52]
  wire [7:0] _GEN_2548 = opcode_3 == 4'hf ? _GEN_1906 : _GEN_2386; // @[executor.scala 466:52]
  wire [7:0] _GEN_2549 = opcode_3 == 4'hf ? _GEN_1907 : _GEN_2387; // @[executor.scala 466:52]
  wire [7:0] _GEN_2550 = opcode_3 == 4'hf ? _GEN_1908 : _GEN_2388; // @[executor.scala 466:52]
  wire [7:0] _GEN_2551 = opcode_3 == 4'hf ? _GEN_1909 : _GEN_2389; // @[executor.scala 466:52]
  wire [7:0] _GEN_2552 = opcode_3 == 4'hf ? _GEN_1910 : _GEN_2390; // @[executor.scala 466:52]
  wire [7:0] _GEN_2553 = opcode_3 == 4'hf ? _GEN_1911 : _GEN_2391; // @[executor.scala 466:52]
  wire [7:0] _GEN_2554 = opcode_3 == 4'hf ? _GEN_1912 : _GEN_2392; // @[executor.scala 466:52]
  wire [7:0] _GEN_2555 = opcode_3 == 4'hf ? _GEN_1913 : _GEN_2393; // @[executor.scala 466:52]
  wire [7:0] _GEN_2556 = opcode_3 == 4'hf ? _GEN_1914 : _GEN_2394; // @[executor.scala 466:52]
  wire [7:0] _GEN_2557 = opcode_3 == 4'hf ? _GEN_1915 : _GEN_2395; // @[executor.scala 466:52]
  wire [7:0] _GEN_2558 = opcode_3 == 4'hf ? _GEN_1916 : _GEN_2396; // @[executor.scala 466:52]
  wire [7:0] _GEN_2559 = opcode_3 == 4'hf ? _GEN_1917 : _GEN_2397; // @[executor.scala 466:52]
  wire [7:0] _GEN_2560 = opcode_3 == 4'hf ? _GEN_1918 : _GEN_2398; // @[executor.scala 466:52]
  wire [7:0] _GEN_2561 = opcode_3 == 4'hf ? _GEN_1919 : _GEN_2399; // @[executor.scala 466:52]
  wire [7:0] _GEN_2562 = opcode_3 == 4'hf ? _GEN_1920 : _GEN_2400; // @[executor.scala 466:52]
  wire [7:0] _GEN_2563 = opcode_3 == 4'hf ? _GEN_1921 : _GEN_2401; // @[executor.scala 466:52]
  wire [7:0] _GEN_2564 = opcode_3 == 4'hf ? _GEN_1922 : _GEN_2402; // @[executor.scala 466:52]
  wire [7:0] _GEN_2565 = opcode_3 == 4'hf ? _GEN_1923 : _GEN_2403; // @[executor.scala 466:52]
  wire [7:0] _GEN_2566 = opcode_3 == 4'hf ? _GEN_1924 : _GEN_2404; // @[executor.scala 466:52]
  wire [7:0] _GEN_2567 = opcode_3 == 4'hf ? _GEN_1925 : _GEN_2405; // @[executor.scala 466:52]
  assign io_pipe_phv_out_data_0 = phv_is_valid_processor ? _GEN_2411 : phv_data_0; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_1 = phv_is_valid_processor ? _GEN_2410 : phv_data_1; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_2 = phv_is_valid_processor ? _GEN_2409 : phv_data_2; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_3 = phv_is_valid_processor ? _GEN_2408 : phv_data_3; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_4 = phv_is_valid_processor ? _GEN_2415 : phv_data_4; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_5 = phv_is_valid_processor ? _GEN_2414 : phv_data_5; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_6 = phv_is_valid_processor ? _GEN_2413 : phv_data_6; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_7 = phv_is_valid_processor ? _GEN_2412 : phv_data_7; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_8 = phv_is_valid_processor ? _GEN_2419 : phv_data_8; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_9 = phv_is_valid_processor ? _GEN_2418 : phv_data_9; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_10 = phv_is_valid_processor ? _GEN_2417 : phv_data_10; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_11 = phv_is_valid_processor ? _GEN_2416 : phv_data_11; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_12 = phv_is_valid_processor ? _GEN_2423 : phv_data_12; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_13 = phv_is_valid_processor ? _GEN_2422 : phv_data_13; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_14 = phv_is_valid_processor ? _GEN_2421 : phv_data_14; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_15 = phv_is_valid_processor ? _GEN_2420 : phv_data_15; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_16 = phv_is_valid_processor ? _GEN_2427 : phv_data_16; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_17 = phv_is_valid_processor ? _GEN_2426 : phv_data_17; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_18 = phv_is_valid_processor ? _GEN_2425 : phv_data_18; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_19 = phv_is_valid_processor ? _GEN_2424 : phv_data_19; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_20 = phv_is_valid_processor ? _GEN_2431 : phv_data_20; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_21 = phv_is_valid_processor ? _GEN_2430 : phv_data_21; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_22 = phv_is_valid_processor ? _GEN_2429 : phv_data_22; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_23 = phv_is_valid_processor ? _GEN_2428 : phv_data_23; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_24 = phv_is_valid_processor ? _GEN_2435 : phv_data_24; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_25 = phv_is_valid_processor ? _GEN_2434 : phv_data_25; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_26 = phv_is_valid_processor ? _GEN_2433 : phv_data_26; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_27 = phv_is_valid_processor ? _GEN_2432 : phv_data_27; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_28 = phv_is_valid_processor ? _GEN_2439 : phv_data_28; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_29 = phv_is_valid_processor ? _GEN_2438 : phv_data_29; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_30 = phv_is_valid_processor ? _GEN_2437 : phv_data_30; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_31 = phv_is_valid_processor ? _GEN_2436 : phv_data_31; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_32 = phv_is_valid_processor ? _GEN_2443 : phv_data_32; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_33 = phv_is_valid_processor ? _GEN_2442 : phv_data_33; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_34 = phv_is_valid_processor ? _GEN_2441 : phv_data_34; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_35 = phv_is_valid_processor ? _GEN_2440 : phv_data_35; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_36 = phv_is_valid_processor ? _GEN_2447 : phv_data_36; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_37 = phv_is_valid_processor ? _GEN_2446 : phv_data_37; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_38 = phv_is_valid_processor ? _GEN_2445 : phv_data_38; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_39 = phv_is_valid_processor ? _GEN_2444 : phv_data_39; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_40 = phv_is_valid_processor ? _GEN_2451 : phv_data_40; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_41 = phv_is_valid_processor ? _GEN_2450 : phv_data_41; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_42 = phv_is_valid_processor ? _GEN_2449 : phv_data_42; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_43 = phv_is_valid_processor ? _GEN_2448 : phv_data_43; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_44 = phv_is_valid_processor ? _GEN_2455 : phv_data_44; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_45 = phv_is_valid_processor ? _GEN_2454 : phv_data_45; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_46 = phv_is_valid_processor ? _GEN_2453 : phv_data_46; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_47 = phv_is_valid_processor ? _GEN_2452 : phv_data_47; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_48 = phv_is_valid_processor ? _GEN_2459 : phv_data_48; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_49 = phv_is_valid_processor ? _GEN_2458 : phv_data_49; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_50 = phv_is_valid_processor ? _GEN_2457 : phv_data_50; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_51 = phv_is_valid_processor ? _GEN_2456 : phv_data_51; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_52 = phv_is_valid_processor ? _GEN_2463 : phv_data_52; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_53 = phv_is_valid_processor ? _GEN_2462 : phv_data_53; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_54 = phv_is_valid_processor ? _GEN_2461 : phv_data_54; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_55 = phv_is_valid_processor ? _GEN_2460 : phv_data_55; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_56 = phv_is_valid_processor ? _GEN_2467 : phv_data_56; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_57 = phv_is_valid_processor ? _GEN_2466 : phv_data_57; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_58 = phv_is_valid_processor ? _GEN_2465 : phv_data_58; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_59 = phv_is_valid_processor ? _GEN_2464 : phv_data_59; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_60 = phv_is_valid_processor ? _GEN_2471 : phv_data_60; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_61 = phv_is_valid_processor ? _GEN_2470 : phv_data_61; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_62 = phv_is_valid_processor ? _GEN_2469 : phv_data_62; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_63 = phv_is_valid_processor ? _GEN_2468 : phv_data_63; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_64 = phv_is_valid_processor ? _GEN_2475 : phv_data_64; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_65 = phv_is_valid_processor ? _GEN_2474 : phv_data_65; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_66 = phv_is_valid_processor ? _GEN_2473 : phv_data_66; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_67 = phv_is_valid_processor ? _GEN_2472 : phv_data_67; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_68 = phv_is_valid_processor ? _GEN_2479 : phv_data_68; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_69 = phv_is_valid_processor ? _GEN_2478 : phv_data_69; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_70 = phv_is_valid_processor ? _GEN_2477 : phv_data_70; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_71 = phv_is_valid_processor ? _GEN_2476 : phv_data_71; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_72 = phv_is_valid_processor ? _GEN_2483 : phv_data_72; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_73 = phv_is_valid_processor ? _GEN_2482 : phv_data_73; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_74 = phv_is_valid_processor ? _GEN_2481 : phv_data_74; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_75 = phv_is_valid_processor ? _GEN_2480 : phv_data_75; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_76 = phv_is_valid_processor ? _GEN_2487 : phv_data_76; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_77 = phv_is_valid_processor ? _GEN_2486 : phv_data_77; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_78 = phv_is_valid_processor ? _GEN_2485 : phv_data_78; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_79 = phv_is_valid_processor ? _GEN_2484 : phv_data_79; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_80 = phv_is_valid_processor ? _GEN_2491 : phv_data_80; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_81 = phv_is_valid_processor ? _GEN_2490 : phv_data_81; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_82 = phv_is_valid_processor ? _GEN_2489 : phv_data_82; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_83 = phv_is_valid_processor ? _GEN_2488 : phv_data_83; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_84 = phv_is_valid_processor ? _GEN_2495 : phv_data_84; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_85 = phv_is_valid_processor ? _GEN_2494 : phv_data_85; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_86 = phv_is_valid_processor ? _GEN_2493 : phv_data_86; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_87 = phv_is_valid_processor ? _GEN_2492 : phv_data_87; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_88 = phv_is_valid_processor ? _GEN_2499 : phv_data_88; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_89 = phv_is_valid_processor ? _GEN_2498 : phv_data_89; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_90 = phv_is_valid_processor ? _GEN_2497 : phv_data_90; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_91 = phv_is_valid_processor ? _GEN_2496 : phv_data_91; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_92 = phv_is_valid_processor ? _GEN_2503 : phv_data_92; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_93 = phv_is_valid_processor ? _GEN_2502 : phv_data_93; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_94 = phv_is_valid_processor ? _GEN_2501 : phv_data_94; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_95 = phv_is_valid_processor ? _GEN_2500 : phv_data_95; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_96 = phv_is_valid_processor ? _GEN_2507 : phv_data_96; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_97 = phv_is_valid_processor ? _GEN_2506 : phv_data_97; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_98 = phv_is_valid_processor ? _GEN_2505 : phv_data_98; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_99 = phv_is_valid_processor ? _GEN_2504 : phv_data_99; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_100 = phv_is_valid_processor ? _GEN_2511 : phv_data_100; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_101 = phv_is_valid_processor ? _GEN_2510 : phv_data_101; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_102 = phv_is_valid_processor ? _GEN_2509 : phv_data_102; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_103 = phv_is_valid_processor ? _GEN_2508 : phv_data_103; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_104 = phv_is_valid_processor ? _GEN_2515 : phv_data_104; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_105 = phv_is_valid_processor ? _GEN_2514 : phv_data_105; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_106 = phv_is_valid_processor ? _GEN_2513 : phv_data_106; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_107 = phv_is_valid_processor ? _GEN_2512 : phv_data_107; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_108 = phv_is_valid_processor ? _GEN_2519 : phv_data_108; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_109 = phv_is_valid_processor ? _GEN_2518 : phv_data_109; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_110 = phv_is_valid_processor ? _GEN_2517 : phv_data_110; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_111 = phv_is_valid_processor ? _GEN_2516 : phv_data_111; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_112 = phv_is_valid_processor ? _GEN_2523 : phv_data_112; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_113 = phv_is_valid_processor ? _GEN_2522 : phv_data_113; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_114 = phv_is_valid_processor ? _GEN_2521 : phv_data_114; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_115 = phv_is_valid_processor ? _GEN_2520 : phv_data_115; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_116 = phv_is_valid_processor ? _GEN_2527 : phv_data_116; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_117 = phv_is_valid_processor ? _GEN_2526 : phv_data_117; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_118 = phv_is_valid_processor ? _GEN_2525 : phv_data_118; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_119 = phv_is_valid_processor ? _GEN_2524 : phv_data_119; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_120 = phv_is_valid_processor ? _GEN_2531 : phv_data_120; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_121 = phv_is_valid_processor ? _GEN_2530 : phv_data_121; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_122 = phv_is_valid_processor ? _GEN_2529 : phv_data_122; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_123 = phv_is_valid_processor ? _GEN_2528 : phv_data_123; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_124 = phv_is_valid_processor ? _GEN_2535 : phv_data_124; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_125 = phv_is_valid_processor ? _GEN_2534 : phv_data_125; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_126 = phv_is_valid_processor ? _GEN_2533 : phv_data_126; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_127 = phv_is_valid_processor ? _GEN_2532 : phv_data_127; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_128 = phv_is_valid_processor ? _GEN_2539 : phv_data_128; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_129 = phv_is_valid_processor ? _GEN_2538 : phv_data_129; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_130 = phv_is_valid_processor ? _GEN_2537 : phv_data_130; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_131 = phv_is_valid_processor ? _GEN_2536 : phv_data_131; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_132 = phv_is_valid_processor ? _GEN_2543 : phv_data_132; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_133 = phv_is_valid_processor ? _GEN_2542 : phv_data_133; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_134 = phv_is_valid_processor ? _GEN_2541 : phv_data_134; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_135 = phv_is_valid_processor ? _GEN_2540 : phv_data_135; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_136 = phv_is_valid_processor ? _GEN_2547 : phv_data_136; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_137 = phv_is_valid_processor ? _GEN_2546 : phv_data_137; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_138 = phv_is_valid_processor ? _GEN_2545 : phv_data_138; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_139 = phv_is_valid_processor ? _GEN_2544 : phv_data_139; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_140 = phv_is_valid_processor ? _GEN_2551 : phv_data_140; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_141 = phv_is_valid_processor ? _GEN_2550 : phv_data_141; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_142 = phv_is_valid_processor ? _GEN_2549 : phv_data_142; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_143 = phv_is_valid_processor ? _GEN_2548 : phv_data_143; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_144 = phv_is_valid_processor ? _GEN_2555 : phv_data_144; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_145 = phv_is_valid_processor ? _GEN_2554 : phv_data_145; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_146 = phv_is_valid_processor ? _GEN_2553 : phv_data_146; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_147 = phv_is_valid_processor ? _GEN_2552 : phv_data_147; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_148 = phv_is_valid_processor ? _GEN_2559 : phv_data_148; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_149 = phv_is_valid_processor ? _GEN_2558 : phv_data_149; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_150 = phv_is_valid_processor ? _GEN_2557 : phv_data_150; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_151 = phv_is_valid_processor ? _GEN_2556 : phv_data_151; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_152 = phv_is_valid_processor ? _GEN_2563 : phv_data_152; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_153 = phv_is_valid_processor ? _GEN_2562 : phv_data_153; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_154 = phv_is_valid_processor ? _GEN_2561 : phv_data_154; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_155 = phv_is_valid_processor ? _GEN_2560 : phv_data_155; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_156 = phv_is_valid_processor ? _GEN_2567 : phv_data_156; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_157 = phv_is_valid_processor ? _GEN_2566 : phv_data_157; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_158 = phv_is_valid_processor ? _GEN_2565 : phv_data_158; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_159 = phv_is_valid_processor ? _GEN_2564 : phv_data_159; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_header_0 = phv_header_0; // @[executor.scala 450:25]
  assign io_pipe_phv_out_header_1 = phv_header_1; // @[executor.scala 450:25]
  assign io_pipe_phv_out_header_2 = phv_header_2; // @[executor.scala 450:25]
  assign io_pipe_phv_out_header_3 = phv_header_3; // @[executor.scala 450:25]
  assign io_pipe_phv_out_header_4 = phv_header_4; // @[executor.scala 450:25]
  assign io_pipe_phv_out_header_5 = phv_header_5; // @[executor.scala 450:25]
  assign io_pipe_phv_out_header_6 = phv_header_6; // @[executor.scala 450:25]
  assign io_pipe_phv_out_header_7 = phv_header_7; // @[executor.scala 450:25]
  assign io_pipe_phv_out_header_8 = phv_header_8; // @[executor.scala 450:25]
  assign io_pipe_phv_out_header_9 = phv_header_9; // @[executor.scala 450:25]
  assign io_pipe_phv_out_header_10 = phv_header_10; // @[executor.scala 450:25]
  assign io_pipe_phv_out_header_11 = phv_header_11; // @[executor.scala 450:25]
  assign io_pipe_phv_out_header_12 = phv_header_12; // @[executor.scala 450:25]
  assign io_pipe_phv_out_header_13 = phv_header_13; // @[executor.scala 450:25]
  assign io_pipe_phv_out_header_14 = phv_header_14; // @[executor.scala 450:25]
  assign io_pipe_phv_out_header_15 = phv_header_15; // @[executor.scala 450:25]
  assign io_pipe_phv_out_parse_current_state = phv_parse_current_state; // @[executor.scala 450:25]
  assign io_pipe_phv_out_parse_current_offset = phv_parse_current_offset; // @[executor.scala 450:25]
  assign io_pipe_phv_out_parse_transition_field = phv_parse_transition_field; // @[executor.scala 450:25]
  assign io_pipe_phv_out_next_processor_id = phv_is_valid_processor ? _GEN_2406 : phv_next_processor_id; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_next_config_id = phv_is_valid_processor ? _GEN_2407 : phv_next_config_id; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_valid = phv_valid; // @[executor.scala 450:25]
  always @(posedge clock) begin
    phv_data_0 <= io_pipe_phv_in_data_0; // @[executor.scala 449:13]
    phv_data_1 <= io_pipe_phv_in_data_1; // @[executor.scala 449:13]
    phv_data_2 <= io_pipe_phv_in_data_2; // @[executor.scala 449:13]
    phv_data_3 <= io_pipe_phv_in_data_3; // @[executor.scala 449:13]
    phv_data_4 <= io_pipe_phv_in_data_4; // @[executor.scala 449:13]
    phv_data_5 <= io_pipe_phv_in_data_5; // @[executor.scala 449:13]
    phv_data_6 <= io_pipe_phv_in_data_6; // @[executor.scala 449:13]
    phv_data_7 <= io_pipe_phv_in_data_7; // @[executor.scala 449:13]
    phv_data_8 <= io_pipe_phv_in_data_8; // @[executor.scala 449:13]
    phv_data_9 <= io_pipe_phv_in_data_9; // @[executor.scala 449:13]
    phv_data_10 <= io_pipe_phv_in_data_10; // @[executor.scala 449:13]
    phv_data_11 <= io_pipe_phv_in_data_11; // @[executor.scala 449:13]
    phv_data_12 <= io_pipe_phv_in_data_12; // @[executor.scala 449:13]
    phv_data_13 <= io_pipe_phv_in_data_13; // @[executor.scala 449:13]
    phv_data_14 <= io_pipe_phv_in_data_14; // @[executor.scala 449:13]
    phv_data_15 <= io_pipe_phv_in_data_15; // @[executor.scala 449:13]
    phv_data_16 <= io_pipe_phv_in_data_16; // @[executor.scala 449:13]
    phv_data_17 <= io_pipe_phv_in_data_17; // @[executor.scala 449:13]
    phv_data_18 <= io_pipe_phv_in_data_18; // @[executor.scala 449:13]
    phv_data_19 <= io_pipe_phv_in_data_19; // @[executor.scala 449:13]
    phv_data_20 <= io_pipe_phv_in_data_20; // @[executor.scala 449:13]
    phv_data_21 <= io_pipe_phv_in_data_21; // @[executor.scala 449:13]
    phv_data_22 <= io_pipe_phv_in_data_22; // @[executor.scala 449:13]
    phv_data_23 <= io_pipe_phv_in_data_23; // @[executor.scala 449:13]
    phv_data_24 <= io_pipe_phv_in_data_24; // @[executor.scala 449:13]
    phv_data_25 <= io_pipe_phv_in_data_25; // @[executor.scala 449:13]
    phv_data_26 <= io_pipe_phv_in_data_26; // @[executor.scala 449:13]
    phv_data_27 <= io_pipe_phv_in_data_27; // @[executor.scala 449:13]
    phv_data_28 <= io_pipe_phv_in_data_28; // @[executor.scala 449:13]
    phv_data_29 <= io_pipe_phv_in_data_29; // @[executor.scala 449:13]
    phv_data_30 <= io_pipe_phv_in_data_30; // @[executor.scala 449:13]
    phv_data_31 <= io_pipe_phv_in_data_31; // @[executor.scala 449:13]
    phv_data_32 <= io_pipe_phv_in_data_32; // @[executor.scala 449:13]
    phv_data_33 <= io_pipe_phv_in_data_33; // @[executor.scala 449:13]
    phv_data_34 <= io_pipe_phv_in_data_34; // @[executor.scala 449:13]
    phv_data_35 <= io_pipe_phv_in_data_35; // @[executor.scala 449:13]
    phv_data_36 <= io_pipe_phv_in_data_36; // @[executor.scala 449:13]
    phv_data_37 <= io_pipe_phv_in_data_37; // @[executor.scala 449:13]
    phv_data_38 <= io_pipe_phv_in_data_38; // @[executor.scala 449:13]
    phv_data_39 <= io_pipe_phv_in_data_39; // @[executor.scala 449:13]
    phv_data_40 <= io_pipe_phv_in_data_40; // @[executor.scala 449:13]
    phv_data_41 <= io_pipe_phv_in_data_41; // @[executor.scala 449:13]
    phv_data_42 <= io_pipe_phv_in_data_42; // @[executor.scala 449:13]
    phv_data_43 <= io_pipe_phv_in_data_43; // @[executor.scala 449:13]
    phv_data_44 <= io_pipe_phv_in_data_44; // @[executor.scala 449:13]
    phv_data_45 <= io_pipe_phv_in_data_45; // @[executor.scala 449:13]
    phv_data_46 <= io_pipe_phv_in_data_46; // @[executor.scala 449:13]
    phv_data_47 <= io_pipe_phv_in_data_47; // @[executor.scala 449:13]
    phv_data_48 <= io_pipe_phv_in_data_48; // @[executor.scala 449:13]
    phv_data_49 <= io_pipe_phv_in_data_49; // @[executor.scala 449:13]
    phv_data_50 <= io_pipe_phv_in_data_50; // @[executor.scala 449:13]
    phv_data_51 <= io_pipe_phv_in_data_51; // @[executor.scala 449:13]
    phv_data_52 <= io_pipe_phv_in_data_52; // @[executor.scala 449:13]
    phv_data_53 <= io_pipe_phv_in_data_53; // @[executor.scala 449:13]
    phv_data_54 <= io_pipe_phv_in_data_54; // @[executor.scala 449:13]
    phv_data_55 <= io_pipe_phv_in_data_55; // @[executor.scala 449:13]
    phv_data_56 <= io_pipe_phv_in_data_56; // @[executor.scala 449:13]
    phv_data_57 <= io_pipe_phv_in_data_57; // @[executor.scala 449:13]
    phv_data_58 <= io_pipe_phv_in_data_58; // @[executor.scala 449:13]
    phv_data_59 <= io_pipe_phv_in_data_59; // @[executor.scala 449:13]
    phv_data_60 <= io_pipe_phv_in_data_60; // @[executor.scala 449:13]
    phv_data_61 <= io_pipe_phv_in_data_61; // @[executor.scala 449:13]
    phv_data_62 <= io_pipe_phv_in_data_62; // @[executor.scala 449:13]
    phv_data_63 <= io_pipe_phv_in_data_63; // @[executor.scala 449:13]
    phv_data_64 <= io_pipe_phv_in_data_64; // @[executor.scala 449:13]
    phv_data_65 <= io_pipe_phv_in_data_65; // @[executor.scala 449:13]
    phv_data_66 <= io_pipe_phv_in_data_66; // @[executor.scala 449:13]
    phv_data_67 <= io_pipe_phv_in_data_67; // @[executor.scala 449:13]
    phv_data_68 <= io_pipe_phv_in_data_68; // @[executor.scala 449:13]
    phv_data_69 <= io_pipe_phv_in_data_69; // @[executor.scala 449:13]
    phv_data_70 <= io_pipe_phv_in_data_70; // @[executor.scala 449:13]
    phv_data_71 <= io_pipe_phv_in_data_71; // @[executor.scala 449:13]
    phv_data_72 <= io_pipe_phv_in_data_72; // @[executor.scala 449:13]
    phv_data_73 <= io_pipe_phv_in_data_73; // @[executor.scala 449:13]
    phv_data_74 <= io_pipe_phv_in_data_74; // @[executor.scala 449:13]
    phv_data_75 <= io_pipe_phv_in_data_75; // @[executor.scala 449:13]
    phv_data_76 <= io_pipe_phv_in_data_76; // @[executor.scala 449:13]
    phv_data_77 <= io_pipe_phv_in_data_77; // @[executor.scala 449:13]
    phv_data_78 <= io_pipe_phv_in_data_78; // @[executor.scala 449:13]
    phv_data_79 <= io_pipe_phv_in_data_79; // @[executor.scala 449:13]
    phv_data_80 <= io_pipe_phv_in_data_80; // @[executor.scala 449:13]
    phv_data_81 <= io_pipe_phv_in_data_81; // @[executor.scala 449:13]
    phv_data_82 <= io_pipe_phv_in_data_82; // @[executor.scala 449:13]
    phv_data_83 <= io_pipe_phv_in_data_83; // @[executor.scala 449:13]
    phv_data_84 <= io_pipe_phv_in_data_84; // @[executor.scala 449:13]
    phv_data_85 <= io_pipe_phv_in_data_85; // @[executor.scala 449:13]
    phv_data_86 <= io_pipe_phv_in_data_86; // @[executor.scala 449:13]
    phv_data_87 <= io_pipe_phv_in_data_87; // @[executor.scala 449:13]
    phv_data_88 <= io_pipe_phv_in_data_88; // @[executor.scala 449:13]
    phv_data_89 <= io_pipe_phv_in_data_89; // @[executor.scala 449:13]
    phv_data_90 <= io_pipe_phv_in_data_90; // @[executor.scala 449:13]
    phv_data_91 <= io_pipe_phv_in_data_91; // @[executor.scala 449:13]
    phv_data_92 <= io_pipe_phv_in_data_92; // @[executor.scala 449:13]
    phv_data_93 <= io_pipe_phv_in_data_93; // @[executor.scala 449:13]
    phv_data_94 <= io_pipe_phv_in_data_94; // @[executor.scala 449:13]
    phv_data_95 <= io_pipe_phv_in_data_95; // @[executor.scala 449:13]
    phv_data_96 <= io_pipe_phv_in_data_96; // @[executor.scala 449:13]
    phv_data_97 <= io_pipe_phv_in_data_97; // @[executor.scala 449:13]
    phv_data_98 <= io_pipe_phv_in_data_98; // @[executor.scala 449:13]
    phv_data_99 <= io_pipe_phv_in_data_99; // @[executor.scala 449:13]
    phv_data_100 <= io_pipe_phv_in_data_100; // @[executor.scala 449:13]
    phv_data_101 <= io_pipe_phv_in_data_101; // @[executor.scala 449:13]
    phv_data_102 <= io_pipe_phv_in_data_102; // @[executor.scala 449:13]
    phv_data_103 <= io_pipe_phv_in_data_103; // @[executor.scala 449:13]
    phv_data_104 <= io_pipe_phv_in_data_104; // @[executor.scala 449:13]
    phv_data_105 <= io_pipe_phv_in_data_105; // @[executor.scala 449:13]
    phv_data_106 <= io_pipe_phv_in_data_106; // @[executor.scala 449:13]
    phv_data_107 <= io_pipe_phv_in_data_107; // @[executor.scala 449:13]
    phv_data_108 <= io_pipe_phv_in_data_108; // @[executor.scala 449:13]
    phv_data_109 <= io_pipe_phv_in_data_109; // @[executor.scala 449:13]
    phv_data_110 <= io_pipe_phv_in_data_110; // @[executor.scala 449:13]
    phv_data_111 <= io_pipe_phv_in_data_111; // @[executor.scala 449:13]
    phv_data_112 <= io_pipe_phv_in_data_112; // @[executor.scala 449:13]
    phv_data_113 <= io_pipe_phv_in_data_113; // @[executor.scala 449:13]
    phv_data_114 <= io_pipe_phv_in_data_114; // @[executor.scala 449:13]
    phv_data_115 <= io_pipe_phv_in_data_115; // @[executor.scala 449:13]
    phv_data_116 <= io_pipe_phv_in_data_116; // @[executor.scala 449:13]
    phv_data_117 <= io_pipe_phv_in_data_117; // @[executor.scala 449:13]
    phv_data_118 <= io_pipe_phv_in_data_118; // @[executor.scala 449:13]
    phv_data_119 <= io_pipe_phv_in_data_119; // @[executor.scala 449:13]
    phv_data_120 <= io_pipe_phv_in_data_120; // @[executor.scala 449:13]
    phv_data_121 <= io_pipe_phv_in_data_121; // @[executor.scala 449:13]
    phv_data_122 <= io_pipe_phv_in_data_122; // @[executor.scala 449:13]
    phv_data_123 <= io_pipe_phv_in_data_123; // @[executor.scala 449:13]
    phv_data_124 <= io_pipe_phv_in_data_124; // @[executor.scala 449:13]
    phv_data_125 <= io_pipe_phv_in_data_125; // @[executor.scala 449:13]
    phv_data_126 <= io_pipe_phv_in_data_126; // @[executor.scala 449:13]
    phv_data_127 <= io_pipe_phv_in_data_127; // @[executor.scala 449:13]
    phv_data_128 <= io_pipe_phv_in_data_128; // @[executor.scala 449:13]
    phv_data_129 <= io_pipe_phv_in_data_129; // @[executor.scala 449:13]
    phv_data_130 <= io_pipe_phv_in_data_130; // @[executor.scala 449:13]
    phv_data_131 <= io_pipe_phv_in_data_131; // @[executor.scala 449:13]
    phv_data_132 <= io_pipe_phv_in_data_132; // @[executor.scala 449:13]
    phv_data_133 <= io_pipe_phv_in_data_133; // @[executor.scala 449:13]
    phv_data_134 <= io_pipe_phv_in_data_134; // @[executor.scala 449:13]
    phv_data_135 <= io_pipe_phv_in_data_135; // @[executor.scala 449:13]
    phv_data_136 <= io_pipe_phv_in_data_136; // @[executor.scala 449:13]
    phv_data_137 <= io_pipe_phv_in_data_137; // @[executor.scala 449:13]
    phv_data_138 <= io_pipe_phv_in_data_138; // @[executor.scala 449:13]
    phv_data_139 <= io_pipe_phv_in_data_139; // @[executor.scala 449:13]
    phv_data_140 <= io_pipe_phv_in_data_140; // @[executor.scala 449:13]
    phv_data_141 <= io_pipe_phv_in_data_141; // @[executor.scala 449:13]
    phv_data_142 <= io_pipe_phv_in_data_142; // @[executor.scala 449:13]
    phv_data_143 <= io_pipe_phv_in_data_143; // @[executor.scala 449:13]
    phv_data_144 <= io_pipe_phv_in_data_144; // @[executor.scala 449:13]
    phv_data_145 <= io_pipe_phv_in_data_145; // @[executor.scala 449:13]
    phv_data_146 <= io_pipe_phv_in_data_146; // @[executor.scala 449:13]
    phv_data_147 <= io_pipe_phv_in_data_147; // @[executor.scala 449:13]
    phv_data_148 <= io_pipe_phv_in_data_148; // @[executor.scala 449:13]
    phv_data_149 <= io_pipe_phv_in_data_149; // @[executor.scala 449:13]
    phv_data_150 <= io_pipe_phv_in_data_150; // @[executor.scala 449:13]
    phv_data_151 <= io_pipe_phv_in_data_151; // @[executor.scala 449:13]
    phv_data_152 <= io_pipe_phv_in_data_152; // @[executor.scala 449:13]
    phv_data_153 <= io_pipe_phv_in_data_153; // @[executor.scala 449:13]
    phv_data_154 <= io_pipe_phv_in_data_154; // @[executor.scala 449:13]
    phv_data_155 <= io_pipe_phv_in_data_155; // @[executor.scala 449:13]
    phv_data_156 <= io_pipe_phv_in_data_156; // @[executor.scala 449:13]
    phv_data_157 <= io_pipe_phv_in_data_157; // @[executor.scala 449:13]
    phv_data_158 <= io_pipe_phv_in_data_158; // @[executor.scala 449:13]
    phv_data_159 <= io_pipe_phv_in_data_159; // @[executor.scala 449:13]
    phv_header_0 <= io_pipe_phv_in_header_0; // @[executor.scala 449:13]
    phv_header_1 <= io_pipe_phv_in_header_1; // @[executor.scala 449:13]
    phv_header_2 <= io_pipe_phv_in_header_2; // @[executor.scala 449:13]
    phv_header_3 <= io_pipe_phv_in_header_3; // @[executor.scala 449:13]
    phv_header_4 <= io_pipe_phv_in_header_4; // @[executor.scala 449:13]
    phv_header_5 <= io_pipe_phv_in_header_5; // @[executor.scala 449:13]
    phv_header_6 <= io_pipe_phv_in_header_6; // @[executor.scala 449:13]
    phv_header_7 <= io_pipe_phv_in_header_7; // @[executor.scala 449:13]
    phv_header_8 <= io_pipe_phv_in_header_8; // @[executor.scala 449:13]
    phv_header_9 <= io_pipe_phv_in_header_9; // @[executor.scala 449:13]
    phv_header_10 <= io_pipe_phv_in_header_10; // @[executor.scala 449:13]
    phv_header_11 <= io_pipe_phv_in_header_11; // @[executor.scala 449:13]
    phv_header_12 <= io_pipe_phv_in_header_12; // @[executor.scala 449:13]
    phv_header_13 <= io_pipe_phv_in_header_13; // @[executor.scala 449:13]
    phv_header_14 <= io_pipe_phv_in_header_14; // @[executor.scala 449:13]
    phv_header_15 <= io_pipe_phv_in_header_15; // @[executor.scala 449:13]
    phv_parse_current_state <= io_pipe_phv_in_parse_current_state; // @[executor.scala 449:13]
    phv_parse_current_offset <= io_pipe_phv_in_parse_current_offset; // @[executor.scala 449:13]
    phv_parse_transition_field <= io_pipe_phv_in_parse_transition_field; // @[executor.scala 449:13]
    phv_next_processor_id <= io_pipe_phv_in_next_processor_id; // @[executor.scala 449:13]
    phv_next_config_id <= io_pipe_phv_in_next_config_id; // @[executor.scala 449:13]
    phv_is_valid_processor <= io_pipe_phv_in_is_valid_processor; // @[executor.scala 449:13]
    phv_valid <= io_pipe_phv_in_valid; // @[executor.scala 449:13]
    vliw_0 <= io_vliw_in_0; // @[executor.scala 453:14]
    vliw_1 <= io_vliw_in_1; // @[executor.scala 453:14]
    vliw_2 <= io_vliw_in_2; // @[executor.scala 453:14]
    vliw_3 <= io_vliw_in_3; // @[executor.scala 453:14]
    field_0 <= io_field_in_0; // @[executor.scala 455:15]
    field_1 <= io_field_in_1; // @[executor.scala 455:15]
    field_2 <= io_field_in_2; // @[executor.scala 455:15]
    field_3 <= io_field_in_3; // @[executor.scala 455:15]
    mask_0 <= io_mask_in_0; // @[executor.scala 457:14]
    mask_1 <= io_mask_in_1; // @[executor.scala 457:14]
    mask_2 <= io_mask_in_2; // @[executor.scala 457:14]
    mask_3 <= io_mask_in_3; // @[executor.scala 457:14]
    dst_offset_0 <= io_dst_offset_in_0; // @[executor.scala 459:20]
    dst_offset_1 <= io_dst_offset_in_1; // @[executor.scala 459:20]
    dst_offset_2 <= io_dst_offset_in_2; // @[executor.scala 459:20]
    dst_offset_3 <= io_dst_offset_in_3; // @[executor.scala 459:20]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  phv_data_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  phv_data_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  phv_data_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  phv_data_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  phv_data_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  phv_data_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  phv_data_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  phv_data_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  phv_data_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  phv_data_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  phv_data_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  phv_data_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  phv_data_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  phv_data_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  phv_data_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  phv_data_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  phv_data_16 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  phv_data_17 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  phv_data_18 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  phv_data_19 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  phv_data_20 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  phv_data_21 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  phv_data_22 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  phv_data_23 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  phv_data_24 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  phv_data_25 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  phv_data_26 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  phv_data_27 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  phv_data_28 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  phv_data_29 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  phv_data_30 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  phv_data_31 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  phv_data_32 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  phv_data_33 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  phv_data_34 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  phv_data_35 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  phv_data_36 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  phv_data_37 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  phv_data_38 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  phv_data_39 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  phv_data_40 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  phv_data_41 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  phv_data_42 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  phv_data_43 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  phv_data_44 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  phv_data_45 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  phv_data_46 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  phv_data_47 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  phv_data_48 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  phv_data_49 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  phv_data_50 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  phv_data_51 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  phv_data_52 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  phv_data_53 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  phv_data_54 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  phv_data_55 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  phv_data_56 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  phv_data_57 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  phv_data_58 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  phv_data_59 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  phv_data_60 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  phv_data_61 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  phv_data_62 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  phv_data_63 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  phv_data_64 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  phv_data_65 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  phv_data_66 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  phv_data_67 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  phv_data_68 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  phv_data_69 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  phv_data_70 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  phv_data_71 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  phv_data_72 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  phv_data_73 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  phv_data_74 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  phv_data_75 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  phv_data_76 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  phv_data_77 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  phv_data_78 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  phv_data_79 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  phv_data_80 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  phv_data_81 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  phv_data_82 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  phv_data_83 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  phv_data_84 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  phv_data_85 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  phv_data_86 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  phv_data_87 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  phv_data_88 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  phv_data_89 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  phv_data_90 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  phv_data_91 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  phv_data_92 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  phv_data_93 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  phv_data_94 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  phv_data_95 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  phv_data_96 = _RAND_96[7:0];
  _RAND_97 = {1{`RANDOM}};
  phv_data_97 = _RAND_97[7:0];
  _RAND_98 = {1{`RANDOM}};
  phv_data_98 = _RAND_98[7:0];
  _RAND_99 = {1{`RANDOM}};
  phv_data_99 = _RAND_99[7:0];
  _RAND_100 = {1{`RANDOM}};
  phv_data_100 = _RAND_100[7:0];
  _RAND_101 = {1{`RANDOM}};
  phv_data_101 = _RAND_101[7:0];
  _RAND_102 = {1{`RANDOM}};
  phv_data_102 = _RAND_102[7:0];
  _RAND_103 = {1{`RANDOM}};
  phv_data_103 = _RAND_103[7:0];
  _RAND_104 = {1{`RANDOM}};
  phv_data_104 = _RAND_104[7:0];
  _RAND_105 = {1{`RANDOM}};
  phv_data_105 = _RAND_105[7:0];
  _RAND_106 = {1{`RANDOM}};
  phv_data_106 = _RAND_106[7:0];
  _RAND_107 = {1{`RANDOM}};
  phv_data_107 = _RAND_107[7:0];
  _RAND_108 = {1{`RANDOM}};
  phv_data_108 = _RAND_108[7:0];
  _RAND_109 = {1{`RANDOM}};
  phv_data_109 = _RAND_109[7:0];
  _RAND_110 = {1{`RANDOM}};
  phv_data_110 = _RAND_110[7:0];
  _RAND_111 = {1{`RANDOM}};
  phv_data_111 = _RAND_111[7:0];
  _RAND_112 = {1{`RANDOM}};
  phv_data_112 = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  phv_data_113 = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  phv_data_114 = _RAND_114[7:0];
  _RAND_115 = {1{`RANDOM}};
  phv_data_115 = _RAND_115[7:0];
  _RAND_116 = {1{`RANDOM}};
  phv_data_116 = _RAND_116[7:0];
  _RAND_117 = {1{`RANDOM}};
  phv_data_117 = _RAND_117[7:0];
  _RAND_118 = {1{`RANDOM}};
  phv_data_118 = _RAND_118[7:0];
  _RAND_119 = {1{`RANDOM}};
  phv_data_119 = _RAND_119[7:0];
  _RAND_120 = {1{`RANDOM}};
  phv_data_120 = _RAND_120[7:0];
  _RAND_121 = {1{`RANDOM}};
  phv_data_121 = _RAND_121[7:0];
  _RAND_122 = {1{`RANDOM}};
  phv_data_122 = _RAND_122[7:0];
  _RAND_123 = {1{`RANDOM}};
  phv_data_123 = _RAND_123[7:0];
  _RAND_124 = {1{`RANDOM}};
  phv_data_124 = _RAND_124[7:0];
  _RAND_125 = {1{`RANDOM}};
  phv_data_125 = _RAND_125[7:0];
  _RAND_126 = {1{`RANDOM}};
  phv_data_126 = _RAND_126[7:0];
  _RAND_127 = {1{`RANDOM}};
  phv_data_127 = _RAND_127[7:0];
  _RAND_128 = {1{`RANDOM}};
  phv_data_128 = _RAND_128[7:0];
  _RAND_129 = {1{`RANDOM}};
  phv_data_129 = _RAND_129[7:0];
  _RAND_130 = {1{`RANDOM}};
  phv_data_130 = _RAND_130[7:0];
  _RAND_131 = {1{`RANDOM}};
  phv_data_131 = _RAND_131[7:0];
  _RAND_132 = {1{`RANDOM}};
  phv_data_132 = _RAND_132[7:0];
  _RAND_133 = {1{`RANDOM}};
  phv_data_133 = _RAND_133[7:0];
  _RAND_134 = {1{`RANDOM}};
  phv_data_134 = _RAND_134[7:0];
  _RAND_135 = {1{`RANDOM}};
  phv_data_135 = _RAND_135[7:0];
  _RAND_136 = {1{`RANDOM}};
  phv_data_136 = _RAND_136[7:0];
  _RAND_137 = {1{`RANDOM}};
  phv_data_137 = _RAND_137[7:0];
  _RAND_138 = {1{`RANDOM}};
  phv_data_138 = _RAND_138[7:0];
  _RAND_139 = {1{`RANDOM}};
  phv_data_139 = _RAND_139[7:0];
  _RAND_140 = {1{`RANDOM}};
  phv_data_140 = _RAND_140[7:0];
  _RAND_141 = {1{`RANDOM}};
  phv_data_141 = _RAND_141[7:0];
  _RAND_142 = {1{`RANDOM}};
  phv_data_142 = _RAND_142[7:0];
  _RAND_143 = {1{`RANDOM}};
  phv_data_143 = _RAND_143[7:0];
  _RAND_144 = {1{`RANDOM}};
  phv_data_144 = _RAND_144[7:0];
  _RAND_145 = {1{`RANDOM}};
  phv_data_145 = _RAND_145[7:0];
  _RAND_146 = {1{`RANDOM}};
  phv_data_146 = _RAND_146[7:0];
  _RAND_147 = {1{`RANDOM}};
  phv_data_147 = _RAND_147[7:0];
  _RAND_148 = {1{`RANDOM}};
  phv_data_148 = _RAND_148[7:0];
  _RAND_149 = {1{`RANDOM}};
  phv_data_149 = _RAND_149[7:0];
  _RAND_150 = {1{`RANDOM}};
  phv_data_150 = _RAND_150[7:0];
  _RAND_151 = {1{`RANDOM}};
  phv_data_151 = _RAND_151[7:0];
  _RAND_152 = {1{`RANDOM}};
  phv_data_152 = _RAND_152[7:0];
  _RAND_153 = {1{`RANDOM}};
  phv_data_153 = _RAND_153[7:0];
  _RAND_154 = {1{`RANDOM}};
  phv_data_154 = _RAND_154[7:0];
  _RAND_155 = {1{`RANDOM}};
  phv_data_155 = _RAND_155[7:0];
  _RAND_156 = {1{`RANDOM}};
  phv_data_156 = _RAND_156[7:0];
  _RAND_157 = {1{`RANDOM}};
  phv_data_157 = _RAND_157[7:0];
  _RAND_158 = {1{`RANDOM}};
  phv_data_158 = _RAND_158[7:0];
  _RAND_159 = {1{`RANDOM}};
  phv_data_159 = _RAND_159[7:0];
  _RAND_160 = {1{`RANDOM}};
  phv_header_0 = _RAND_160[15:0];
  _RAND_161 = {1{`RANDOM}};
  phv_header_1 = _RAND_161[15:0];
  _RAND_162 = {1{`RANDOM}};
  phv_header_2 = _RAND_162[15:0];
  _RAND_163 = {1{`RANDOM}};
  phv_header_3 = _RAND_163[15:0];
  _RAND_164 = {1{`RANDOM}};
  phv_header_4 = _RAND_164[15:0];
  _RAND_165 = {1{`RANDOM}};
  phv_header_5 = _RAND_165[15:0];
  _RAND_166 = {1{`RANDOM}};
  phv_header_6 = _RAND_166[15:0];
  _RAND_167 = {1{`RANDOM}};
  phv_header_7 = _RAND_167[15:0];
  _RAND_168 = {1{`RANDOM}};
  phv_header_8 = _RAND_168[15:0];
  _RAND_169 = {1{`RANDOM}};
  phv_header_9 = _RAND_169[15:0];
  _RAND_170 = {1{`RANDOM}};
  phv_header_10 = _RAND_170[15:0];
  _RAND_171 = {1{`RANDOM}};
  phv_header_11 = _RAND_171[15:0];
  _RAND_172 = {1{`RANDOM}};
  phv_header_12 = _RAND_172[15:0];
  _RAND_173 = {1{`RANDOM}};
  phv_header_13 = _RAND_173[15:0];
  _RAND_174 = {1{`RANDOM}};
  phv_header_14 = _RAND_174[15:0];
  _RAND_175 = {1{`RANDOM}};
  phv_header_15 = _RAND_175[15:0];
  _RAND_176 = {1{`RANDOM}};
  phv_parse_current_state = _RAND_176[7:0];
  _RAND_177 = {1{`RANDOM}};
  phv_parse_current_offset = _RAND_177[7:0];
  _RAND_178 = {1{`RANDOM}};
  phv_parse_transition_field = _RAND_178[15:0];
  _RAND_179 = {1{`RANDOM}};
  phv_next_processor_id = _RAND_179[3:0];
  _RAND_180 = {1{`RANDOM}};
  phv_next_config_id = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  phv_is_valid_processor = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  phv_valid = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  vliw_0 = _RAND_183[31:0];
  _RAND_184 = {1{`RANDOM}};
  vliw_1 = _RAND_184[31:0];
  _RAND_185 = {1{`RANDOM}};
  vliw_2 = _RAND_185[31:0];
  _RAND_186 = {1{`RANDOM}};
  vliw_3 = _RAND_186[31:0];
  _RAND_187 = {1{`RANDOM}};
  field_0 = _RAND_187[31:0];
  _RAND_188 = {1{`RANDOM}};
  field_1 = _RAND_188[31:0];
  _RAND_189 = {1{`RANDOM}};
  field_2 = _RAND_189[31:0];
  _RAND_190 = {1{`RANDOM}};
  field_3 = _RAND_190[31:0];
  _RAND_191 = {1{`RANDOM}};
  mask_0 = _RAND_191[3:0];
  _RAND_192 = {1{`RANDOM}};
  mask_1 = _RAND_192[3:0];
  _RAND_193 = {1{`RANDOM}};
  mask_2 = _RAND_193[3:0];
  _RAND_194 = {1{`RANDOM}};
  mask_3 = _RAND_194[3:0];
  _RAND_195 = {1{`RANDOM}};
  dst_offset_0 = _RAND_195[5:0];
  _RAND_196 = {1{`RANDOM}};
  dst_offset_1 = _RAND_196[5:0];
  _RAND_197 = {1{`RANDOM}};
  dst_offset_2 = _RAND_197[5:0];
  _RAND_198 = {1{`RANDOM}};
  dst_offset_3 = _RAND_198[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
