module InPort(
  input        clock,
  input        reset,
  output [7:0] io_phv_out_data_0,
  output [7:0] io_phv_out_data_1,
  output [7:0] io_phv_out_data_2,
  output [7:0] io_phv_out_data_3,
  output [7:0] io_phv_out_data_4,
  output [7:0] io_phv_out_data_5,
  output [7:0] io_phv_out_data_6,
  output [7:0] io_phv_out_data_7,
  output [7:0] io_phv_out_data_8,
  output [7:0] io_phv_out_data_9,
  output [7:0] io_phv_out_data_10,
  output [7:0] io_phv_out_data_11,
  output [7:0] io_phv_out_data_12,
  output [7:0] io_phv_out_data_13,
  output [7:0] io_phv_out_data_14,
  output [7:0] io_phv_out_data_15,
  output [7:0] io_phv_out_data_16,
  output [7:0] io_phv_out_data_17,
  output [7:0] io_phv_out_data_18,
  output [7:0] io_phv_out_data_19,
  output [7:0] io_phv_out_data_20,
  output [7:0] io_phv_out_data_21,
  output [7:0] io_phv_out_data_22,
  output [7:0] io_phv_out_data_23,
  output [7:0] io_phv_out_data_24,
  output [7:0] io_phv_out_data_25,
  output [7:0] io_phv_out_data_26,
  output [7:0] io_phv_out_data_27,
  output [7:0] io_phv_out_data_28,
  output [7:0] io_phv_out_data_29,
  output [7:0] io_phv_out_data_30,
  output [7:0] io_phv_out_data_31,
  output [7:0] io_phv_out_data_32,
  output [7:0] io_phv_out_data_33,
  output [7:0] io_phv_out_data_34,
  output [7:0] io_phv_out_data_35,
  output [7:0] io_phv_out_data_36,
  output [7:0] io_phv_out_data_37,
  output [7:0] io_phv_out_data_38,
  output [7:0] io_phv_out_data_39,
  output [7:0] io_phv_out_data_40,
  output [7:0] io_phv_out_data_41,
  output [7:0] io_phv_out_data_42,
  output [7:0] io_phv_out_data_43,
  output [7:0] io_phv_out_data_44,
  output [7:0] io_phv_out_data_45,
  output [7:0] io_phv_out_data_46,
  output [7:0] io_phv_out_data_47,
  output [7:0] io_phv_out_data_48,
  output [7:0] io_phv_out_data_49,
  output [7:0] io_phv_out_data_50,
  output [7:0] io_phv_out_data_51,
  output [7:0] io_phv_out_data_52,
  output [7:0] io_phv_out_data_53,
  output [7:0] io_phv_out_data_54,
  output [7:0] io_phv_out_data_55,
  output [7:0] io_phv_out_data_56,
  output [7:0] io_phv_out_data_57,
  output [7:0] io_phv_out_data_58,
  output [7:0] io_phv_out_data_59,
  output [7:0] io_phv_out_data_60,
  output [7:0] io_phv_out_data_61,
  output [7:0] io_phv_out_data_62,
  output [7:0] io_phv_out_data_63,
  output [7:0] io_phv_out_data_64,
  output [7:0] io_phv_out_data_65,
  output [7:0] io_phv_out_data_66,
  output [7:0] io_phv_out_data_67,
  output [7:0] io_phv_out_data_68,
  output [7:0] io_phv_out_data_69,
  output [7:0] io_phv_out_data_70,
  output [7:0] io_phv_out_data_71,
  output [7:0] io_phv_out_data_72,
  output [7:0] io_phv_out_data_73,
  output [7:0] io_phv_out_data_74,
  output [7:0] io_phv_out_data_75,
  output [7:0] io_phv_out_data_76,
  output [7:0] io_phv_out_data_77,
  output [7:0] io_phv_out_data_78,
  output [7:0] io_phv_out_data_79,
  output [7:0] io_phv_out_data_80,
  output [7:0] io_phv_out_data_81,
  output [7:0] io_phv_out_data_82,
  output [7:0] io_phv_out_data_83,
  output [7:0] io_phv_out_data_84,
  output [7:0] io_phv_out_data_85,
  output [7:0] io_phv_out_data_86,
  output [7:0] io_phv_out_data_87,
  output [7:0] io_phv_out_data_88,
  output [7:0] io_phv_out_data_89,
  output [7:0] io_phv_out_data_90,
  output [7:0] io_phv_out_data_91,
  output [7:0] io_phv_out_data_92,
  output [7:0] io_phv_out_data_93,
  output [7:0] io_phv_out_data_94,
  output [7:0] io_phv_out_data_95,
  output [7:0] io_phv_out_data_96,
  output [7:0] io_phv_out_data_97,
  output [7:0] io_phv_out_data_98,
  output [7:0] io_phv_out_data_99,
  output [7:0] io_phv_out_data_100,
  output [7:0] io_phv_out_data_101,
  output [7:0] io_phv_out_data_102,
  output [7:0] io_phv_out_data_103,
  output [7:0] io_phv_out_data_104,
  output [7:0] io_phv_out_data_105,
  output [7:0] io_phv_out_data_106,
  output [7:0] io_phv_out_data_107,
  output [7:0] io_phv_out_data_108,
  output [7:0] io_phv_out_data_109,
  output [7:0] io_phv_out_data_110,
  output [7:0] io_phv_out_data_111,
  output [7:0] io_phv_out_data_112,
  output [7:0] io_phv_out_data_113,
  output [7:0] io_phv_out_data_114,
  output [7:0] io_phv_out_data_115,
  output [7:0] io_phv_out_data_116,
  output [7:0] io_phv_out_data_117,
  output [7:0] io_phv_out_data_118,
  output [7:0] io_phv_out_data_119,
  output [7:0] io_phv_out_data_120,
  output [7:0] io_phv_out_data_121,
  output [7:0] io_phv_out_data_122,
  output [7:0] io_phv_out_data_123,
  output [7:0] io_phv_out_data_124,
  output [7:0] io_phv_out_data_125,
  output [7:0] io_phv_out_data_126,
  output [7:0] io_phv_out_data_127
);
  wire  rand_exe_prng_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_1_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_1_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_1_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_1_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_1_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_1_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_1_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_1_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_1_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_1_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_1_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_1_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_1_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_1_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_1_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_1_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_1_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_1_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_2_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_2_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_2_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_2_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_2_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_2_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_2_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_2_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_2_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_2_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_2_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_2_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_2_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_2_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_2_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_2_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_2_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_2_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_3_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_3_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_3_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_3_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_3_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_3_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_3_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_3_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_3_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_3_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_3_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_3_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_3_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_3_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_3_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_3_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_3_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_3_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_4_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_4_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_4_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_4_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_4_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_4_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_4_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_4_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_4_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_4_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_4_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_4_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_4_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_4_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_4_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_4_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_4_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_4_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_5_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_5_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_5_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_5_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_5_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_5_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_5_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_5_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_5_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_5_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_5_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_5_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_5_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_5_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_5_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_5_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_5_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_5_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_6_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_6_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_6_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_6_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_6_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_6_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_6_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_6_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_6_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_6_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_6_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_6_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_6_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_6_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_6_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_6_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_6_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_6_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_7_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_7_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_7_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_7_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_7_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_7_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_7_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_7_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_7_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_7_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_7_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_7_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_7_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_7_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_7_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_7_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_7_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_7_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_8_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_8_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_8_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_8_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_8_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_8_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_8_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_8_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_8_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_8_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_8_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_8_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_8_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_8_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_8_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_8_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_8_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_8_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_9_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_9_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_9_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_9_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_9_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_9_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_9_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_9_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_9_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_9_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_9_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_9_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_9_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_9_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_9_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_9_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_9_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_9_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_10_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_10_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_10_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_10_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_10_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_10_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_10_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_10_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_10_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_10_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_10_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_10_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_10_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_10_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_10_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_10_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_10_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_10_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_11_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_11_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_11_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_11_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_11_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_11_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_11_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_11_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_11_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_11_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_11_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_11_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_11_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_11_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_11_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_11_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_11_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_11_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_12_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_12_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_12_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_12_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_12_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_12_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_12_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_12_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_12_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_12_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_12_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_12_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_12_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_12_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_12_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_12_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_12_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_12_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_13_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_13_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_13_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_13_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_13_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_13_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_13_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_13_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_13_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_13_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_13_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_13_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_13_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_13_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_13_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_13_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_13_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_13_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_14_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_14_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_14_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_14_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_14_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_14_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_14_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_14_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_14_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_14_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_14_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_14_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_14_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_14_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_14_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_14_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_14_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_14_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_15_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_15_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_15_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_15_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_15_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_15_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_15_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_15_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_15_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_15_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_15_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_15_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_15_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_15_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_15_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_15_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_15_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_15_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_16_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_16_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_16_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_16_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_16_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_16_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_16_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_16_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_16_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_16_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_16_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_16_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_16_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_16_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_16_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_16_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_16_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_16_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_17_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_17_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_17_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_17_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_17_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_17_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_17_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_17_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_17_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_17_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_17_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_17_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_17_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_17_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_17_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_17_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_17_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_17_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_18_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_18_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_18_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_18_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_18_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_18_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_18_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_18_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_18_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_18_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_18_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_18_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_18_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_18_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_18_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_18_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_18_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_18_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_19_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_19_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_19_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_19_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_19_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_19_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_19_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_19_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_19_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_19_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_19_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_19_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_19_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_19_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_19_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_19_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_19_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_19_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_20_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_20_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_20_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_20_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_20_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_20_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_20_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_20_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_20_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_20_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_20_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_20_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_20_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_20_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_20_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_20_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_20_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_20_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_21_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_21_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_21_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_21_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_21_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_21_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_21_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_21_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_21_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_21_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_21_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_21_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_21_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_21_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_21_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_21_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_21_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_21_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_22_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_22_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_22_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_22_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_22_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_22_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_22_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_22_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_22_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_22_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_22_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_22_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_22_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_22_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_22_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_22_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_22_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_22_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_23_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_23_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_23_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_23_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_23_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_23_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_23_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_23_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_23_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_23_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_23_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_23_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_23_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_23_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_23_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_23_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_23_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_23_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_24_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_24_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_24_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_24_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_24_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_24_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_24_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_24_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_24_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_24_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_24_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_24_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_24_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_24_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_24_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_24_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_24_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_24_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_25_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_25_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_25_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_25_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_25_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_25_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_25_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_25_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_25_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_25_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_25_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_25_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_25_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_25_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_25_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_25_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_25_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_25_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_26_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_26_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_26_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_26_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_26_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_26_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_26_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_26_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_26_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_26_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_26_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_26_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_26_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_26_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_26_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_26_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_26_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_26_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_27_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_27_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_27_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_27_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_27_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_27_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_27_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_27_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_27_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_27_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_27_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_27_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_27_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_27_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_27_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_27_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_27_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_27_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_28_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_28_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_28_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_28_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_28_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_28_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_28_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_28_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_28_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_28_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_28_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_28_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_28_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_28_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_28_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_28_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_28_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_28_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_29_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_29_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_29_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_29_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_29_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_29_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_29_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_29_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_29_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_29_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_29_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_29_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_29_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_29_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_29_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_29_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_29_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_29_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_30_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_30_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_30_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_30_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_30_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_30_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_30_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_30_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_30_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_30_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_30_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_30_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_30_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_30_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_30_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_30_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_30_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_30_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_31_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_31_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_31_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_31_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_31_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_31_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_31_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_31_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_31_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_31_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_31_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_31_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_31_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_31_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_31_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_31_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_31_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_31_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_32_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_32_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_32_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_32_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_32_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_32_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_32_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_32_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_32_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_32_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_32_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_32_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_32_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_32_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_32_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_32_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_32_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_32_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_33_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_33_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_33_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_33_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_33_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_33_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_33_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_33_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_33_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_33_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_33_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_33_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_33_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_33_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_33_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_33_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_33_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_33_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_34_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_34_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_34_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_34_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_34_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_34_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_34_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_34_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_34_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_34_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_34_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_34_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_34_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_34_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_34_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_34_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_34_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_34_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_35_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_35_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_35_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_35_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_35_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_35_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_35_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_35_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_35_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_35_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_35_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_35_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_35_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_35_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_35_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_35_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_35_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_35_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_36_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_36_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_36_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_36_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_36_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_36_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_36_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_36_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_36_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_36_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_36_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_36_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_36_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_36_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_36_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_36_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_36_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_36_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_37_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_37_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_37_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_37_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_37_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_37_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_37_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_37_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_37_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_37_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_37_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_37_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_37_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_37_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_37_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_37_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_37_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_37_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_38_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_38_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_38_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_38_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_38_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_38_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_38_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_38_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_38_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_38_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_38_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_38_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_38_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_38_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_38_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_38_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_38_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_38_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_39_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_39_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_39_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_39_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_39_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_39_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_39_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_39_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_39_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_39_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_39_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_39_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_39_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_39_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_39_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_39_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_39_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_39_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_40_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_40_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_40_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_40_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_40_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_40_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_40_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_40_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_40_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_40_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_40_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_40_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_40_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_40_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_40_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_40_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_40_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_40_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_41_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_41_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_41_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_41_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_41_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_41_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_41_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_41_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_41_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_41_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_41_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_41_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_41_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_41_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_41_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_41_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_41_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_41_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_42_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_42_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_42_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_42_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_42_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_42_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_42_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_42_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_42_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_42_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_42_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_42_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_42_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_42_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_42_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_42_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_42_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_42_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_43_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_43_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_43_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_43_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_43_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_43_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_43_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_43_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_43_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_43_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_43_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_43_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_43_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_43_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_43_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_43_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_43_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_43_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_44_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_44_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_44_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_44_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_44_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_44_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_44_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_44_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_44_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_44_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_44_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_44_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_44_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_44_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_44_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_44_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_44_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_44_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_45_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_45_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_45_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_45_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_45_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_45_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_45_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_45_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_45_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_45_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_45_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_45_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_45_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_45_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_45_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_45_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_45_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_45_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_46_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_46_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_46_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_46_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_46_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_46_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_46_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_46_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_46_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_46_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_46_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_46_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_46_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_46_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_46_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_46_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_46_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_46_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_47_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_47_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_47_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_47_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_47_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_47_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_47_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_47_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_47_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_47_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_47_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_47_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_47_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_47_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_47_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_47_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_47_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_47_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_48_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_48_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_48_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_48_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_48_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_48_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_48_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_48_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_48_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_48_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_48_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_48_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_48_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_48_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_48_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_48_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_48_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_48_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_49_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_49_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_49_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_49_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_49_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_49_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_49_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_49_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_49_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_49_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_49_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_49_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_49_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_49_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_49_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_49_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_49_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_49_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_50_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_50_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_50_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_50_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_50_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_50_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_50_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_50_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_50_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_50_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_50_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_50_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_50_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_50_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_50_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_50_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_50_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_50_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_51_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_51_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_51_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_51_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_51_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_51_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_51_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_51_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_51_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_51_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_51_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_51_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_51_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_51_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_51_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_51_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_51_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_51_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_52_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_52_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_52_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_52_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_52_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_52_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_52_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_52_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_52_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_52_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_52_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_52_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_52_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_52_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_52_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_52_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_52_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_52_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_53_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_53_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_53_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_53_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_53_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_53_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_53_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_53_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_53_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_53_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_53_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_53_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_53_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_53_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_53_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_53_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_53_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_53_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_54_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_54_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_54_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_54_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_54_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_54_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_54_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_54_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_54_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_54_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_54_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_54_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_54_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_54_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_54_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_54_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_54_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_54_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_55_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_55_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_55_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_55_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_55_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_55_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_55_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_55_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_55_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_55_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_55_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_55_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_55_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_55_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_55_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_55_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_55_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_55_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_56_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_56_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_56_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_56_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_56_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_56_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_56_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_56_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_56_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_56_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_56_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_56_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_56_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_56_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_56_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_56_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_56_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_56_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_57_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_57_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_57_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_57_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_57_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_57_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_57_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_57_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_57_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_57_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_57_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_57_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_57_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_57_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_57_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_57_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_57_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_57_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_58_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_58_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_58_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_58_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_58_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_58_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_58_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_58_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_58_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_58_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_58_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_58_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_58_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_58_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_58_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_58_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_58_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_58_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_59_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_59_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_59_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_59_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_59_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_59_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_59_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_59_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_59_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_59_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_59_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_59_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_59_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_59_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_59_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_59_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_59_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_59_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_60_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_60_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_60_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_60_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_60_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_60_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_60_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_60_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_60_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_60_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_60_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_60_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_60_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_60_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_60_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_60_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_60_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_60_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_61_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_61_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_61_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_61_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_61_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_61_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_61_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_61_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_61_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_61_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_61_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_61_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_61_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_61_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_61_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_61_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_61_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_61_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_62_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_62_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_62_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_62_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_62_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_62_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_62_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_62_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_62_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_62_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_62_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_62_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_62_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_62_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_62_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_62_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_62_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_62_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_63_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_63_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_63_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_63_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_63_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_63_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_63_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_63_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_63_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_63_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_63_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_63_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_63_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_63_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_63_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_63_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_63_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_63_io_out_15; // @[PRNG.scala 82:22]
  wire [7:0] rand_exe_lo = {rand_exe_prng_io_out_7,rand_exe_prng_io_out_6,rand_exe_prng_io_out_5,rand_exe_prng_io_out_4,
    rand_exe_prng_io_out_3,rand_exe_prng_io_out_2,rand_exe_prng_io_out_1,rand_exe_prng_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_0 = {rand_exe_prng_io_out_15,rand_exe_prng_io_out_14,rand_exe_prng_io_out_13,rand_exe_prng_io_out_12,
    rand_exe_prng_io_out_11,rand_exe_prng_io_out_10,rand_exe_prng_io_out_9,rand_exe_prng_io_out_8,rand_exe_lo}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_1 = {rand_exe_prng_1_io_out_7,rand_exe_prng_1_io_out_6,rand_exe_prng_1_io_out_5,
    rand_exe_prng_1_io_out_4,rand_exe_prng_1_io_out_3,rand_exe_prng_1_io_out_2,rand_exe_prng_1_io_out_1,
    rand_exe_prng_1_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_1 = {rand_exe_prng_1_io_out_15,rand_exe_prng_1_io_out_14,rand_exe_prng_1_io_out_13,
    rand_exe_prng_1_io_out_12,rand_exe_prng_1_io_out_11,rand_exe_prng_1_io_out_10,rand_exe_prng_1_io_out_9,
    rand_exe_prng_1_io_out_8,rand_exe_lo_1}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_2 = {rand_exe_prng_2_io_out_7,rand_exe_prng_2_io_out_6,rand_exe_prng_2_io_out_5,
    rand_exe_prng_2_io_out_4,rand_exe_prng_2_io_out_3,rand_exe_prng_2_io_out_2,rand_exe_prng_2_io_out_1,
    rand_exe_prng_2_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_2 = {rand_exe_prng_2_io_out_15,rand_exe_prng_2_io_out_14,rand_exe_prng_2_io_out_13,
    rand_exe_prng_2_io_out_12,rand_exe_prng_2_io_out_11,rand_exe_prng_2_io_out_10,rand_exe_prng_2_io_out_9,
    rand_exe_prng_2_io_out_8,rand_exe_lo_2}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_3 = {rand_exe_prng_3_io_out_7,rand_exe_prng_3_io_out_6,rand_exe_prng_3_io_out_5,
    rand_exe_prng_3_io_out_4,rand_exe_prng_3_io_out_3,rand_exe_prng_3_io_out_2,rand_exe_prng_3_io_out_1,
    rand_exe_prng_3_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_3 = {rand_exe_prng_3_io_out_15,rand_exe_prng_3_io_out_14,rand_exe_prng_3_io_out_13,
    rand_exe_prng_3_io_out_12,rand_exe_prng_3_io_out_11,rand_exe_prng_3_io_out_10,rand_exe_prng_3_io_out_9,
    rand_exe_prng_3_io_out_8,rand_exe_lo_3}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_4 = {rand_exe_prng_4_io_out_7,rand_exe_prng_4_io_out_6,rand_exe_prng_4_io_out_5,
    rand_exe_prng_4_io_out_4,rand_exe_prng_4_io_out_3,rand_exe_prng_4_io_out_2,rand_exe_prng_4_io_out_1,
    rand_exe_prng_4_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_4 = {rand_exe_prng_4_io_out_15,rand_exe_prng_4_io_out_14,rand_exe_prng_4_io_out_13,
    rand_exe_prng_4_io_out_12,rand_exe_prng_4_io_out_11,rand_exe_prng_4_io_out_10,rand_exe_prng_4_io_out_9,
    rand_exe_prng_4_io_out_8,rand_exe_lo_4}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_5 = {rand_exe_prng_5_io_out_7,rand_exe_prng_5_io_out_6,rand_exe_prng_5_io_out_5,
    rand_exe_prng_5_io_out_4,rand_exe_prng_5_io_out_3,rand_exe_prng_5_io_out_2,rand_exe_prng_5_io_out_1,
    rand_exe_prng_5_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_5 = {rand_exe_prng_5_io_out_15,rand_exe_prng_5_io_out_14,rand_exe_prng_5_io_out_13,
    rand_exe_prng_5_io_out_12,rand_exe_prng_5_io_out_11,rand_exe_prng_5_io_out_10,rand_exe_prng_5_io_out_9,
    rand_exe_prng_5_io_out_8,rand_exe_lo_5}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_6 = {rand_exe_prng_6_io_out_7,rand_exe_prng_6_io_out_6,rand_exe_prng_6_io_out_5,
    rand_exe_prng_6_io_out_4,rand_exe_prng_6_io_out_3,rand_exe_prng_6_io_out_2,rand_exe_prng_6_io_out_1,
    rand_exe_prng_6_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_6 = {rand_exe_prng_6_io_out_15,rand_exe_prng_6_io_out_14,rand_exe_prng_6_io_out_13,
    rand_exe_prng_6_io_out_12,rand_exe_prng_6_io_out_11,rand_exe_prng_6_io_out_10,rand_exe_prng_6_io_out_9,
    rand_exe_prng_6_io_out_8,rand_exe_lo_6}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_7 = {rand_exe_prng_7_io_out_7,rand_exe_prng_7_io_out_6,rand_exe_prng_7_io_out_5,
    rand_exe_prng_7_io_out_4,rand_exe_prng_7_io_out_3,rand_exe_prng_7_io_out_2,rand_exe_prng_7_io_out_1,
    rand_exe_prng_7_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_7 = {rand_exe_prng_7_io_out_15,rand_exe_prng_7_io_out_14,rand_exe_prng_7_io_out_13,
    rand_exe_prng_7_io_out_12,rand_exe_prng_7_io_out_11,rand_exe_prng_7_io_out_10,rand_exe_prng_7_io_out_9,
    rand_exe_prng_7_io_out_8,rand_exe_lo_7}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_8 = {rand_exe_prng_8_io_out_7,rand_exe_prng_8_io_out_6,rand_exe_prng_8_io_out_5,
    rand_exe_prng_8_io_out_4,rand_exe_prng_8_io_out_3,rand_exe_prng_8_io_out_2,rand_exe_prng_8_io_out_1,
    rand_exe_prng_8_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_8 = {rand_exe_prng_8_io_out_15,rand_exe_prng_8_io_out_14,rand_exe_prng_8_io_out_13,
    rand_exe_prng_8_io_out_12,rand_exe_prng_8_io_out_11,rand_exe_prng_8_io_out_10,rand_exe_prng_8_io_out_9,
    rand_exe_prng_8_io_out_8,rand_exe_lo_8}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_9 = {rand_exe_prng_9_io_out_7,rand_exe_prng_9_io_out_6,rand_exe_prng_9_io_out_5,
    rand_exe_prng_9_io_out_4,rand_exe_prng_9_io_out_3,rand_exe_prng_9_io_out_2,rand_exe_prng_9_io_out_1,
    rand_exe_prng_9_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_9 = {rand_exe_prng_9_io_out_15,rand_exe_prng_9_io_out_14,rand_exe_prng_9_io_out_13,
    rand_exe_prng_9_io_out_12,rand_exe_prng_9_io_out_11,rand_exe_prng_9_io_out_10,rand_exe_prng_9_io_out_9,
    rand_exe_prng_9_io_out_8,rand_exe_lo_9}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_10 = {rand_exe_prng_10_io_out_7,rand_exe_prng_10_io_out_6,rand_exe_prng_10_io_out_5,
    rand_exe_prng_10_io_out_4,rand_exe_prng_10_io_out_3,rand_exe_prng_10_io_out_2,rand_exe_prng_10_io_out_1,
    rand_exe_prng_10_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_10 = {rand_exe_prng_10_io_out_15,rand_exe_prng_10_io_out_14,rand_exe_prng_10_io_out_13,
    rand_exe_prng_10_io_out_12,rand_exe_prng_10_io_out_11,rand_exe_prng_10_io_out_10,rand_exe_prng_10_io_out_9,
    rand_exe_prng_10_io_out_8,rand_exe_lo_10}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_11 = {rand_exe_prng_11_io_out_7,rand_exe_prng_11_io_out_6,rand_exe_prng_11_io_out_5,
    rand_exe_prng_11_io_out_4,rand_exe_prng_11_io_out_3,rand_exe_prng_11_io_out_2,rand_exe_prng_11_io_out_1,
    rand_exe_prng_11_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_11 = {rand_exe_prng_11_io_out_15,rand_exe_prng_11_io_out_14,rand_exe_prng_11_io_out_13,
    rand_exe_prng_11_io_out_12,rand_exe_prng_11_io_out_11,rand_exe_prng_11_io_out_10,rand_exe_prng_11_io_out_9,
    rand_exe_prng_11_io_out_8,rand_exe_lo_11}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_12 = {rand_exe_prng_12_io_out_7,rand_exe_prng_12_io_out_6,rand_exe_prng_12_io_out_5,
    rand_exe_prng_12_io_out_4,rand_exe_prng_12_io_out_3,rand_exe_prng_12_io_out_2,rand_exe_prng_12_io_out_1,
    rand_exe_prng_12_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_12 = {rand_exe_prng_12_io_out_15,rand_exe_prng_12_io_out_14,rand_exe_prng_12_io_out_13,
    rand_exe_prng_12_io_out_12,rand_exe_prng_12_io_out_11,rand_exe_prng_12_io_out_10,rand_exe_prng_12_io_out_9,
    rand_exe_prng_12_io_out_8,rand_exe_lo_12}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_13 = {rand_exe_prng_13_io_out_7,rand_exe_prng_13_io_out_6,rand_exe_prng_13_io_out_5,
    rand_exe_prng_13_io_out_4,rand_exe_prng_13_io_out_3,rand_exe_prng_13_io_out_2,rand_exe_prng_13_io_out_1,
    rand_exe_prng_13_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_13 = {rand_exe_prng_13_io_out_15,rand_exe_prng_13_io_out_14,rand_exe_prng_13_io_out_13,
    rand_exe_prng_13_io_out_12,rand_exe_prng_13_io_out_11,rand_exe_prng_13_io_out_10,rand_exe_prng_13_io_out_9,
    rand_exe_prng_13_io_out_8,rand_exe_lo_13}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_14 = {rand_exe_prng_14_io_out_7,rand_exe_prng_14_io_out_6,rand_exe_prng_14_io_out_5,
    rand_exe_prng_14_io_out_4,rand_exe_prng_14_io_out_3,rand_exe_prng_14_io_out_2,rand_exe_prng_14_io_out_1,
    rand_exe_prng_14_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_14 = {rand_exe_prng_14_io_out_15,rand_exe_prng_14_io_out_14,rand_exe_prng_14_io_out_13,
    rand_exe_prng_14_io_out_12,rand_exe_prng_14_io_out_11,rand_exe_prng_14_io_out_10,rand_exe_prng_14_io_out_9,
    rand_exe_prng_14_io_out_8,rand_exe_lo_14}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_15 = {rand_exe_prng_15_io_out_7,rand_exe_prng_15_io_out_6,rand_exe_prng_15_io_out_5,
    rand_exe_prng_15_io_out_4,rand_exe_prng_15_io_out_3,rand_exe_prng_15_io_out_2,rand_exe_prng_15_io_out_1,
    rand_exe_prng_15_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_15 = {rand_exe_prng_15_io_out_15,rand_exe_prng_15_io_out_14,rand_exe_prng_15_io_out_13,
    rand_exe_prng_15_io_out_12,rand_exe_prng_15_io_out_11,rand_exe_prng_15_io_out_10,rand_exe_prng_15_io_out_9,
    rand_exe_prng_15_io_out_8,rand_exe_lo_15}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_16 = {rand_exe_prng_16_io_out_7,rand_exe_prng_16_io_out_6,rand_exe_prng_16_io_out_5,
    rand_exe_prng_16_io_out_4,rand_exe_prng_16_io_out_3,rand_exe_prng_16_io_out_2,rand_exe_prng_16_io_out_1,
    rand_exe_prng_16_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_16 = {rand_exe_prng_16_io_out_15,rand_exe_prng_16_io_out_14,rand_exe_prng_16_io_out_13,
    rand_exe_prng_16_io_out_12,rand_exe_prng_16_io_out_11,rand_exe_prng_16_io_out_10,rand_exe_prng_16_io_out_9,
    rand_exe_prng_16_io_out_8,rand_exe_lo_16}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_17 = {rand_exe_prng_17_io_out_7,rand_exe_prng_17_io_out_6,rand_exe_prng_17_io_out_5,
    rand_exe_prng_17_io_out_4,rand_exe_prng_17_io_out_3,rand_exe_prng_17_io_out_2,rand_exe_prng_17_io_out_1,
    rand_exe_prng_17_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_17 = {rand_exe_prng_17_io_out_15,rand_exe_prng_17_io_out_14,rand_exe_prng_17_io_out_13,
    rand_exe_prng_17_io_out_12,rand_exe_prng_17_io_out_11,rand_exe_prng_17_io_out_10,rand_exe_prng_17_io_out_9,
    rand_exe_prng_17_io_out_8,rand_exe_lo_17}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_18 = {rand_exe_prng_18_io_out_7,rand_exe_prng_18_io_out_6,rand_exe_prng_18_io_out_5,
    rand_exe_prng_18_io_out_4,rand_exe_prng_18_io_out_3,rand_exe_prng_18_io_out_2,rand_exe_prng_18_io_out_1,
    rand_exe_prng_18_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_18 = {rand_exe_prng_18_io_out_15,rand_exe_prng_18_io_out_14,rand_exe_prng_18_io_out_13,
    rand_exe_prng_18_io_out_12,rand_exe_prng_18_io_out_11,rand_exe_prng_18_io_out_10,rand_exe_prng_18_io_out_9,
    rand_exe_prng_18_io_out_8,rand_exe_lo_18}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_19 = {rand_exe_prng_19_io_out_7,rand_exe_prng_19_io_out_6,rand_exe_prng_19_io_out_5,
    rand_exe_prng_19_io_out_4,rand_exe_prng_19_io_out_3,rand_exe_prng_19_io_out_2,rand_exe_prng_19_io_out_1,
    rand_exe_prng_19_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_19 = {rand_exe_prng_19_io_out_15,rand_exe_prng_19_io_out_14,rand_exe_prng_19_io_out_13,
    rand_exe_prng_19_io_out_12,rand_exe_prng_19_io_out_11,rand_exe_prng_19_io_out_10,rand_exe_prng_19_io_out_9,
    rand_exe_prng_19_io_out_8,rand_exe_lo_19}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_20 = {rand_exe_prng_20_io_out_7,rand_exe_prng_20_io_out_6,rand_exe_prng_20_io_out_5,
    rand_exe_prng_20_io_out_4,rand_exe_prng_20_io_out_3,rand_exe_prng_20_io_out_2,rand_exe_prng_20_io_out_1,
    rand_exe_prng_20_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_20 = {rand_exe_prng_20_io_out_15,rand_exe_prng_20_io_out_14,rand_exe_prng_20_io_out_13,
    rand_exe_prng_20_io_out_12,rand_exe_prng_20_io_out_11,rand_exe_prng_20_io_out_10,rand_exe_prng_20_io_out_9,
    rand_exe_prng_20_io_out_8,rand_exe_lo_20}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_21 = {rand_exe_prng_21_io_out_7,rand_exe_prng_21_io_out_6,rand_exe_prng_21_io_out_5,
    rand_exe_prng_21_io_out_4,rand_exe_prng_21_io_out_3,rand_exe_prng_21_io_out_2,rand_exe_prng_21_io_out_1,
    rand_exe_prng_21_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_21 = {rand_exe_prng_21_io_out_15,rand_exe_prng_21_io_out_14,rand_exe_prng_21_io_out_13,
    rand_exe_prng_21_io_out_12,rand_exe_prng_21_io_out_11,rand_exe_prng_21_io_out_10,rand_exe_prng_21_io_out_9,
    rand_exe_prng_21_io_out_8,rand_exe_lo_21}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_22 = {rand_exe_prng_22_io_out_7,rand_exe_prng_22_io_out_6,rand_exe_prng_22_io_out_5,
    rand_exe_prng_22_io_out_4,rand_exe_prng_22_io_out_3,rand_exe_prng_22_io_out_2,rand_exe_prng_22_io_out_1,
    rand_exe_prng_22_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_22 = {rand_exe_prng_22_io_out_15,rand_exe_prng_22_io_out_14,rand_exe_prng_22_io_out_13,
    rand_exe_prng_22_io_out_12,rand_exe_prng_22_io_out_11,rand_exe_prng_22_io_out_10,rand_exe_prng_22_io_out_9,
    rand_exe_prng_22_io_out_8,rand_exe_lo_22}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_23 = {rand_exe_prng_23_io_out_7,rand_exe_prng_23_io_out_6,rand_exe_prng_23_io_out_5,
    rand_exe_prng_23_io_out_4,rand_exe_prng_23_io_out_3,rand_exe_prng_23_io_out_2,rand_exe_prng_23_io_out_1,
    rand_exe_prng_23_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_23 = {rand_exe_prng_23_io_out_15,rand_exe_prng_23_io_out_14,rand_exe_prng_23_io_out_13,
    rand_exe_prng_23_io_out_12,rand_exe_prng_23_io_out_11,rand_exe_prng_23_io_out_10,rand_exe_prng_23_io_out_9,
    rand_exe_prng_23_io_out_8,rand_exe_lo_23}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_24 = {rand_exe_prng_24_io_out_7,rand_exe_prng_24_io_out_6,rand_exe_prng_24_io_out_5,
    rand_exe_prng_24_io_out_4,rand_exe_prng_24_io_out_3,rand_exe_prng_24_io_out_2,rand_exe_prng_24_io_out_1,
    rand_exe_prng_24_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_24 = {rand_exe_prng_24_io_out_15,rand_exe_prng_24_io_out_14,rand_exe_prng_24_io_out_13,
    rand_exe_prng_24_io_out_12,rand_exe_prng_24_io_out_11,rand_exe_prng_24_io_out_10,rand_exe_prng_24_io_out_9,
    rand_exe_prng_24_io_out_8,rand_exe_lo_24}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_25 = {rand_exe_prng_25_io_out_7,rand_exe_prng_25_io_out_6,rand_exe_prng_25_io_out_5,
    rand_exe_prng_25_io_out_4,rand_exe_prng_25_io_out_3,rand_exe_prng_25_io_out_2,rand_exe_prng_25_io_out_1,
    rand_exe_prng_25_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_25 = {rand_exe_prng_25_io_out_15,rand_exe_prng_25_io_out_14,rand_exe_prng_25_io_out_13,
    rand_exe_prng_25_io_out_12,rand_exe_prng_25_io_out_11,rand_exe_prng_25_io_out_10,rand_exe_prng_25_io_out_9,
    rand_exe_prng_25_io_out_8,rand_exe_lo_25}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_26 = {rand_exe_prng_26_io_out_7,rand_exe_prng_26_io_out_6,rand_exe_prng_26_io_out_5,
    rand_exe_prng_26_io_out_4,rand_exe_prng_26_io_out_3,rand_exe_prng_26_io_out_2,rand_exe_prng_26_io_out_1,
    rand_exe_prng_26_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_26 = {rand_exe_prng_26_io_out_15,rand_exe_prng_26_io_out_14,rand_exe_prng_26_io_out_13,
    rand_exe_prng_26_io_out_12,rand_exe_prng_26_io_out_11,rand_exe_prng_26_io_out_10,rand_exe_prng_26_io_out_9,
    rand_exe_prng_26_io_out_8,rand_exe_lo_26}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_27 = {rand_exe_prng_27_io_out_7,rand_exe_prng_27_io_out_6,rand_exe_prng_27_io_out_5,
    rand_exe_prng_27_io_out_4,rand_exe_prng_27_io_out_3,rand_exe_prng_27_io_out_2,rand_exe_prng_27_io_out_1,
    rand_exe_prng_27_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_27 = {rand_exe_prng_27_io_out_15,rand_exe_prng_27_io_out_14,rand_exe_prng_27_io_out_13,
    rand_exe_prng_27_io_out_12,rand_exe_prng_27_io_out_11,rand_exe_prng_27_io_out_10,rand_exe_prng_27_io_out_9,
    rand_exe_prng_27_io_out_8,rand_exe_lo_27}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_28 = {rand_exe_prng_28_io_out_7,rand_exe_prng_28_io_out_6,rand_exe_prng_28_io_out_5,
    rand_exe_prng_28_io_out_4,rand_exe_prng_28_io_out_3,rand_exe_prng_28_io_out_2,rand_exe_prng_28_io_out_1,
    rand_exe_prng_28_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_28 = {rand_exe_prng_28_io_out_15,rand_exe_prng_28_io_out_14,rand_exe_prng_28_io_out_13,
    rand_exe_prng_28_io_out_12,rand_exe_prng_28_io_out_11,rand_exe_prng_28_io_out_10,rand_exe_prng_28_io_out_9,
    rand_exe_prng_28_io_out_8,rand_exe_lo_28}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_29 = {rand_exe_prng_29_io_out_7,rand_exe_prng_29_io_out_6,rand_exe_prng_29_io_out_5,
    rand_exe_prng_29_io_out_4,rand_exe_prng_29_io_out_3,rand_exe_prng_29_io_out_2,rand_exe_prng_29_io_out_1,
    rand_exe_prng_29_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_29 = {rand_exe_prng_29_io_out_15,rand_exe_prng_29_io_out_14,rand_exe_prng_29_io_out_13,
    rand_exe_prng_29_io_out_12,rand_exe_prng_29_io_out_11,rand_exe_prng_29_io_out_10,rand_exe_prng_29_io_out_9,
    rand_exe_prng_29_io_out_8,rand_exe_lo_29}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_30 = {rand_exe_prng_30_io_out_7,rand_exe_prng_30_io_out_6,rand_exe_prng_30_io_out_5,
    rand_exe_prng_30_io_out_4,rand_exe_prng_30_io_out_3,rand_exe_prng_30_io_out_2,rand_exe_prng_30_io_out_1,
    rand_exe_prng_30_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_30 = {rand_exe_prng_30_io_out_15,rand_exe_prng_30_io_out_14,rand_exe_prng_30_io_out_13,
    rand_exe_prng_30_io_out_12,rand_exe_prng_30_io_out_11,rand_exe_prng_30_io_out_10,rand_exe_prng_30_io_out_9,
    rand_exe_prng_30_io_out_8,rand_exe_lo_30}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_31 = {rand_exe_prng_31_io_out_7,rand_exe_prng_31_io_out_6,rand_exe_prng_31_io_out_5,
    rand_exe_prng_31_io_out_4,rand_exe_prng_31_io_out_3,rand_exe_prng_31_io_out_2,rand_exe_prng_31_io_out_1,
    rand_exe_prng_31_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_31 = {rand_exe_prng_31_io_out_15,rand_exe_prng_31_io_out_14,rand_exe_prng_31_io_out_13,
    rand_exe_prng_31_io_out_12,rand_exe_prng_31_io_out_11,rand_exe_prng_31_io_out_10,rand_exe_prng_31_io_out_9,
    rand_exe_prng_31_io_out_8,rand_exe_lo_31}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_32 = {rand_exe_prng_32_io_out_7,rand_exe_prng_32_io_out_6,rand_exe_prng_32_io_out_5,
    rand_exe_prng_32_io_out_4,rand_exe_prng_32_io_out_3,rand_exe_prng_32_io_out_2,rand_exe_prng_32_io_out_1,
    rand_exe_prng_32_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_32 = {rand_exe_prng_32_io_out_15,rand_exe_prng_32_io_out_14,rand_exe_prng_32_io_out_13,
    rand_exe_prng_32_io_out_12,rand_exe_prng_32_io_out_11,rand_exe_prng_32_io_out_10,rand_exe_prng_32_io_out_9,
    rand_exe_prng_32_io_out_8,rand_exe_lo_32}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_33 = {rand_exe_prng_33_io_out_7,rand_exe_prng_33_io_out_6,rand_exe_prng_33_io_out_5,
    rand_exe_prng_33_io_out_4,rand_exe_prng_33_io_out_3,rand_exe_prng_33_io_out_2,rand_exe_prng_33_io_out_1,
    rand_exe_prng_33_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_33 = {rand_exe_prng_33_io_out_15,rand_exe_prng_33_io_out_14,rand_exe_prng_33_io_out_13,
    rand_exe_prng_33_io_out_12,rand_exe_prng_33_io_out_11,rand_exe_prng_33_io_out_10,rand_exe_prng_33_io_out_9,
    rand_exe_prng_33_io_out_8,rand_exe_lo_33}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_34 = {rand_exe_prng_34_io_out_7,rand_exe_prng_34_io_out_6,rand_exe_prng_34_io_out_5,
    rand_exe_prng_34_io_out_4,rand_exe_prng_34_io_out_3,rand_exe_prng_34_io_out_2,rand_exe_prng_34_io_out_1,
    rand_exe_prng_34_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_34 = {rand_exe_prng_34_io_out_15,rand_exe_prng_34_io_out_14,rand_exe_prng_34_io_out_13,
    rand_exe_prng_34_io_out_12,rand_exe_prng_34_io_out_11,rand_exe_prng_34_io_out_10,rand_exe_prng_34_io_out_9,
    rand_exe_prng_34_io_out_8,rand_exe_lo_34}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_35 = {rand_exe_prng_35_io_out_7,rand_exe_prng_35_io_out_6,rand_exe_prng_35_io_out_5,
    rand_exe_prng_35_io_out_4,rand_exe_prng_35_io_out_3,rand_exe_prng_35_io_out_2,rand_exe_prng_35_io_out_1,
    rand_exe_prng_35_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_35 = {rand_exe_prng_35_io_out_15,rand_exe_prng_35_io_out_14,rand_exe_prng_35_io_out_13,
    rand_exe_prng_35_io_out_12,rand_exe_prng_35_io_out_11,rand_exe_prng_35_io_out_10,rand_exe_prng_35_io_out_9,
    rand_exe_prng_35_io_out_8,rand_exe_lo_35}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_36 = {rand_exe_prng_36_io_out_7,rand_exe_prng_36_io_out_6,rand_exe_prng_36_io_out_5,
    rand_exe_prng_36_io_out_4,rand_exe_prng_36_io_out_3,rand_exe_prng_36_io_out_2,rand_exe_prng_36_io_out_1,
    rand_exe_prng_36_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_36 = {rand_exe_prng_36_io_out_15,rand_exe_prng_36_io_out_14,rand_exe_prng_36_io_out_13,
    rand_exe_prng_36_io_out_12,rand_exe_prng_36_io_out_11,rand_exe_prng_36_io_out_10,rand_exe_prng_36_io_out_9,
    rand_exe_prng_36_io_out_8,rand_exe_lo_36}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_37 = {rand_exe_prng_37_io_out_7,rand_exe_prng_37_io_out_6,rand_exe_prng_37_io_out_5,
    rand_exe_prng_37_io_out_4,rand_exe_prng_37_io_out_3,rand_exe_prng_37_io_out_2,rand_exe_prng_37_io_out_1,
    rand_exe_prng_37_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_37 = {rand_exe_prng_37_io_out_15,rand_exe_prng_37_io_out_14,rand_exe_prng_37_io_out_13,
    rand_exe_prng_37_io_out_12,rand_exe_prng_37_io_out_11,rand_exe_prng_37_io_out_10,rand_exe_prng_37_io_out_9,
    rand_exe_prng_37_io_out_8,rand_exe_lo_37}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_38 = {rand_exe_prng_38_io_out_7,rand_exe_prng_38_io_out_6,rand_exe_prng_38_io_out_5,
    rand_exe_prng_38_io_out_4,rand_exe_prng_38_io_out_3,rand_exe_prng_38_io_out_2,rand_exe_prng_38_io_out_1,
    rand_exe_prng_38_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_38 = {rand_exe_prng_38_io_out_15,rand_exe_prng_38_io_out_14,rand_exe_prng_38_io_out_13,
    rand_exe_prng_38_io_out_12,rand_exe_prng_38_io_out_11,rand_exe_prng_38_io_out_10,rand_exe_prng_38_io_out_9,
    rand_exe_prng_38_io_out_8,rand_exe_lo_38}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_39 = {rand_exe_prng_39_io_out_7,rand_exe_prng_39_io_out_6,rand_exe_prng_39_io_out_5,
    rand_exe_prng_39_io_out_4,rand_exe_prng_39_io_out_3,rand_exe_prng_39_io_out_2,rand_exe_prng_39_io_out_1,
    rand_exe_prng_39_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_39 = {rand_exe_prng_39_io_out_15,rand_exe_prng_39_io_out_14,rand_exe_prng_39_io_out_13,
    rand_exe_prng_39_io_out_12,rand_exe_prng_39_io_out_11,rand_exe_prng_39_io_out_10,rand_exe_prng_39_io_out_9,
    rand_exe_prng_39_io_out_8,rand_exe_lo_39}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_40 = {rand_exe_prng_40_io_out_7,rand_exe_prng_40_io_out_6,rand_exe_prng_40_io_out_5,
    rand_exe_prng_40_io_out_4,rand_exe_prng_40_io_out_3,rand_exe_prng_40_io_out_2,rand_exe_prng_40_io_out_1,
    rand_exe_prng_40_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_40 = {rand_exe_prng_40_io_out_15,rand_exe_prng_40_io_out_14,rand_exe_prng_40_io_out_13,
    rand_exe_prng_40_io_out_12,rand_exe_prng_40_io_out_11,rand_exe_prng_40_io_out_10,rand_exe_prng_40_io_out_9,
    rand_exe_prng_40_io_out_8,rand_exe_lo_40}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_41 = {rand_exe_prng_41_io_out_7,rand_exe_prng_41_io_out_6,rand_exe_prng_41_io_out_5,
    rand_exe_prng_41_io_out_4,rand_exe_prng_41_io_out_3,rand_exe_prng_41_io_out_2,rand_exe_prng_41_io_out_1,
    rand_exe_prng_41_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_41 = {rand_exe_prng_41_io_out_15,rand_exe_prng_41_io_out_14,rand_exe_prng_41_io_out_13,
    rand_exe_prng_41_io_out_12,rand_exe_prng_41_io_out_11,rand_exe_prng_41_io_out_10,rand_exe_prng_41_io_out_9,
    rand_exe_prng_41_io_out_8,rand_exe_lo_41}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_42 = {rand_exe_prng_42_io_out_7,rand_exe_prng_42_io_out_6,rand_exe_prng_42_io_out_5,
    rand_exe_prng_42_io_out_4,rand_exe_prng_42_io_out_3,rand_exe_prng_42_io_out_2,rand_exe_prng_42_io_out_1,
    rand_exe_prng_42_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_42 = {rand_exe_prng_42_io_out_15,rand_exe_prng_42_io_out_14,rand_exe_prng_42_io_out_13,
    rand_exe_prng_42_io_out_12,rand_exe_prng_42_io_out_11,rand_exe_prng_42_io_out_10,rand_exe_prng_42_io_out_9,
    rand_exe_prng_42_io_out_8,rand_exe_lo_42}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_43 = {rand_exe_prng_43_io_out_7,rand_exe_prng_43_io_out_6,rand_exe_prng_43_io_out_5,
    rand_exe_prng_43_io_out_4,rand_exe_prng_43_io_out_3,rand_exe_prng_43_io_out_2,rand_exe_prng_43_io_out_1,
    rand_exe_prng_43_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_43 = {rand_exe_prng_43_io_out_15,rand_exe_prng_43_io_out_14,rand_exe_prng_43_io_out_13,
    rand_exe_prng_43_io_out_12,rand_exe_prng_43_io_out_11,rand_exe_prng_43_io_out_10,rand_exe_prng_43_io_out_9,
    rand_exe_prng_43_io_out_8,rand_exe_lo_43}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_44 = {rand_exe_prng_44_io_out_7,rand_exe_prng_44_io_out_6,rand_exe_prng_44_io_out_5,
    rand_exe_prng_44_io_out_4,rand_exe_prng_44_io_out_3,rand_exe_prng_44_io_out_2,rand_exe_prng_44_io_out_1,
    rand_exe_prng_44_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_44 = {rand_exe_prng_44_io_out_15,rand_exe_prng_44_io_out_14,rand_exe_prng_44_io_out_13,
    rand_exe_prng_44_io_out_12,rand_exe_prng_44_io_out_11,rand_exe_prng_44_io_out_10,rand_exe_prng_44_io_out_9,
    rand_exe_prng_44_io_out_8,rand_exe_lo_44}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_45 = {rand_exe_prng_45_io_out_7,rand_exe_prng_45_io_out_6,rand_exe_prng_45_io_out_5,
    rand_exe_prng_45_io_out_4,rand_exe_prng_45_io_out_3,rand_exe_prng_45_io_out_2,rand_exe_prng_45_io_out_1,
    rand_exe_prng_45_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_45 = {rand_exe_prng_45_io_out_15,rand_exe_prng_45_io_out_14,rand_exe_prng_45_io_out_13,
    rand_exe_prng_45_io_out_12,rand_exe_prng_45_io_out_11,rand_exe_prng_45_io_out_10,rand_exe_prng_45_io_out_9,
    rand_exe_prng_45_io_out_8,rand_exe_lo_45}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_46 = {rand_exe_prng_46_io_out_7,rand_exe_prng_46_io_out_6,rand_exe_prng_46_io_out_5,
    rand_exe_prng_46_io_out_4,rand_exe_prng_46_io_out_3,rand_exe_prng_46_io_out_2,rand_exe_prng_46_io_out_1,
    rand_exe_prng_46_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_46 = {rand_exe_prng_46_io_out_15,rand_exe_prng_46_io_out_14,rand_exe_prng_46_io_out_13,
    rand_exe_prng_46_io_out_12,rand_exe_prng_46_io_out_11,rand_exe_prng_46_io_out_10,rand_exe_prng_46_io_out_9,
    rand_exe_prng_46_io_out_8,rand_exe_lo_46}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_47 = {rand_exe_prng_47_io_out_7,rand_exe_prng_47_io_out_6,rand_exe_prng_47_io_out_5,
    rand_exe_prng_47_io_out_4,rand_exe_prng_47_io_out_3,rand_exe_prng_47_io_out_2,rand_exe_prng_47_io_out_1,
    rand_exe_prng_47_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_47 = {rand_exe_prng_47_io_out_15,rand_exe_prng_47_io_out_14,rand_exe_prng_47_io_out_13,
    rand_exe_prng_47_io_out_12,rand_exe_prng_47_io_out_11,rand_exe_prng_47_io_out_10,rand_exe_prng_47_io_out_9,
    rand_exe_prng_47_io_out_8,rand_exe_lo_47}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_48 = {rand_exe_prng_48_io_out_7,rand_exe_prng_48_io_out_6,rand_exe_prng_48_io_out_5,
    rand_exe_prng_48_io_out_4,rand_exe_prng_48_io_out_3,rand_exe_prng_48_io_out_2,rand_exe_prng_48_io_out_1,
    rand_exe_prng_48_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_48 = {rand_exe_prng_48_io_out_15,rand_exe_prng_48_io_out_14,rand_exe_prng_48_io_out_13,
    rand_exe_prng_48_io_out_12,rand_exe_prng_48_io_out_11,rand_exe_prng_48_io_out_10,rand_exe_prng_48_io_out_9,
    rand_exe_prng_48_io_out_8,rand_exe_lo_48}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_49 = {rand_exe_prng_49_io_out_7,rand_exe_prng_49_io_out_6,rand_exe_prng_49_io_out_5,
    rand_exe_prng_49_io_out_4,rand_exe_prng_49_io_out_3,rand_exe_prng_49_io_out_2,rand_exe_prng_49_io_out_1,
    rand_exe_prng_49_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_49 = {rand_exe_prng_49_io_out_15,rand_exe_prng_49_io_out_14,rand_exe_prng_49_io_out_13,
    rand_exe_prng_49_io_out_12,rand_exe_prng_49_io_out_11,rand_exe_prng_49_io_out_10,rand_exe_prng_49_io_out_9,
    rand_exe_prng_49_io_out_8,rand_exe_lo_49}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_50 = {rand_exe_prng_50_io_out_7,rand_exe_prng_50_io_out_6,rand_exe_prng_50_io_out_5,
    rand_exe_prng_50_io_out_4,rand_exe_prng_50_io_out_3,rand_exe_prng_50_io_out_2,rand_exe_prng_50_io_out_1,
    rand_exe_prng_50_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_50 = {rand_exe_prng_50_io_out_15,rand_exe_prng_50_io_out_14,rand_exe_prng_50_io_out_13,
    rand_exe_prng_50_io_out_12,rand_exe_prng_50_io_out_11,rand_exe_prng_50_io_out_10,rand_exe_prng_50_io_out_9,
    rand_exe_prng_50_io_out_8,rand_exe_lo_50}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_51 = {rand_exe_prng_51_io_out_7,rand_exe_prng_51_io_out_6,rand_exe_prng_51_io_out_5,
    rand_exe_prng_51_io_out_4,rand_exe_prng_51_io_out_3,rand_exe_prng_51_io_out_2,rand_exe_prng_51_io_out_1,
    rand_exe_prng_51_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_51 = {rand_exe_prng_51_io_out_15,rand_exe_prng_51_io_out_14,rand_exe_prng_51_io_out_13,
    rand_exe_prng_51_io_out_12,rand_exe_prng_51_io_out_11,rand_exe_prng_51_io_out_10,rand_exe_prng_51_io_out_9,
    rand_exe_prng_51_io_out_8,rand_exe_lo_51}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_52 = {rand_exe_prng_52_io_out_7,rand_exe_prng_52_io_out_6,rand_exe_prng_52_io_out_5,
    rand_exe_prng_52_io_out_4,rand_exe_prng_52_io_out_3,rand_exe_prng_52_io_out_2,rand_exe_prng_52_io_out_1,
    rand_exe_prng_52_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_52 = {rand_exe_prng_52_io_out_15,rand_exe_prng_52_io_out_14,rand_exe_prng_52_io_out_13,
    rand_exe_prng_52_io_out_12,rand_exe_prng_52_io_out_11,rand_exe_prng_52_io_out_10,rand_exe_prng_52_io_out_9,
    rand_exe_prng_52_io_out_8,rand_exe_lo_52}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_53 = {rand_exe_prng_53_io_out_7,rand_exe_prng_53_io_out_6,rand_exe_prng_53_io_out_5,
    rand_exe_prng_53_io_out_4,rand_exe_prng_53_io_out_3,rand_exe_prng_53_io_out_2,rand_exe_prng_53_io_out_1,
    rand_exe_prng_53_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_53 = {rand_exe_prng_53_io_out_15,rand_exe_prng_53_io_out_14,rand_exe_prng_53_io_out_13,
    rand_exe_prng_53_io_out_12,rand_exe_prng_53_io_out_11,rand_exe_prng_53_io_out_10,rand_exe_prng_53_io_out_9,
    rand_exe_prng_53_io_out_8,rand_exe_lo_53}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_54 = {rand_exe_prng_54_io_out_7,rand_exe_prng_54_io_out_6,rand_exe_prng_54_io_out_5,
    rand_exe_prng_54_io_out_4,rand_exe_prng_54_io_out_3,rand_exe_prng_54_io_out_2,rand_exe_prng_54_io_out_1,
    rand_exe_prng_54_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_54 = {rand_exe_prng_54_io_out_15,rand_exe_prng_54_io_out_14,rand_exe_prng_54_io_out_13,
    rand_exe_prng_54_io_out_12,rand_exe_prng_54_io_out_11,rand_exe_prng_54_io_out_10,rand_exe_prng_54_io_out_9,
    rand_exe_prng_54_io_out_8,rand_exe_lo_54}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_55 = {rand_exe_prng_55_io_out_7,rand_exe_prng_55_io_out_6,rand_exe_prng_55_io_out_5,
    rand_exe_prng_55_io_out_4,rand_exe_prng_55_io_out_3,rand_exe_prng_55_io_out_2,rand_exe_prng_55_io_out_1,
    rand_exe_prng_55_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_55 = {rand_exe_prng_55_io_out_15,rand_exe_prng_55_io_out_14,rand_exe_prng_55_io_out_13,
    rand_exe_prng_55_io_out_12,rand_exe_prng_55_io_out_11,rand_exe_prng_55_io_out_10,rand_exe_prng_55_io_out_9,
    rand_exe_prng_55_io_out_8,rand_exe_lo_55}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_56 = {rand_exe_prng_56_io_out_7,rand_exe_prng_56_io_out_6,rand_exe_prng_56_io_out_5,
    rand_exe_prng_56_io_out_4,rand_exe_prng_56_io_out_3,rand_exe_prng_56_io_out_2,rand_exe_prng_56_io_out_1,
    rand_exe_prng_56_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_56 = {rand_exe_prng_56_io_out_15,rand_exe_prng_56_io_out_14,rand_exe_prng_56_io_out_13,
    rand_exe_prng_56_io_out_12,rand_exe_prng_56_io_out_11,rand_exe_prng_56_io_out_10,rand_exe_prng_56_io_out_9,
    rand_exe_prng_56_io_out_8,rand_exe_lo_56}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_57 = {rand_exe_prng_57_io_out_7,rand_exe_prng_57_io_out_6,rand_exe_prng_57_io_out_5,
    rand_exe_prng_57_io_out_4,rand_exe_prng_57_io_out_3,rand_exe_prng_57_io_out_2,rand_exe_prng_57_io_out_1,
    rand_exe_prng_57_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_57 = {rand_exe_prng_57_io_out_15,rand_exe_prng_57_io_out_14,rand_exe_prng_57_io_out_13,
    rand_exe_prng_57_io_out_12,rand_exe_prng_57_io_out_11,rand_exe_prng_57_io_out_10,rand_exe_prng_57_io_out_9,
    rand_exe_prng_57_io_out_8,rand_exe_lo_57}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_58 = {rand_exe_prng_58_io_out_7,rand_exe_prng_58_io_out_6,rand_exe_prng_58_io_out_5,
    rand_exe_prng_58_io_out_4,rand_exe_prng_58_io_out_3,rand_exe_prng_58_io_out_2,rand_exe_prng_58_io_out_1,
    rand_exe_prng_58_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_58 = {rand_exe_prng_58_io_out_15,rand_exe_prng_58_io_out_14,rand_exe_prng_58_io_out_13,
    rand_exe_prng_58_io_out_12,rand_exe_prng_58_io_out_11,rand_exe_prng_58_io_out_10,rand_exe_prng_58_io_out_9,
    rand_exe_prng_58_io_out_8,rand_exe_lo_58}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_59 = {rand_exe_prng_59_io_out_7,rand_exe_prng_59_io_out_6,rand_exe_prng_59_io_out_5,
    rand_exe_prng_59_io_out_4,rand_exe_prng_59_io_out_3,rand_exe_prng_59_io_out_2,rand_exe_prng_59_io_out_1,
    rand_exe_prng_59_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_59 = {rand_exe_prng_59_io_out_15,rand_exe_prng_59_io_out_14,rand_exe_prng_59_io_out_13,
    rand_exe_prng_59_io_out_12,rand_exe_prng_59_io_out_11,rand_exe_prng_59_io_out_10,rand_exe_prng_59_io_out_9,
    rand_exe_prng_59_io_out_8,rand_exe_lo_59}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_60 = {rand_exe_prng_60_io_out_7,rand_exe_prng_60_io_out_6,rand_exe_prng_60_io_out_5,
    rand_exe_prng_60_io_out_4,rand_exe_prng_60_io_out_3,rand_exe_prng_60_io_out_2,rand_exe_prng_60_io_out_1,
    rand_exe_prng_60_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_60 = {rand_exe_prng_60_io_out_15,rand_exe_prng_60_io_out_14,rand_exe_prng_60_io_out_13,
    rand_exe_prng_60_io_out_12,rand_exe_prng_60_io_out_11,rand_exe_prng_60_io_out_10,rand_exe_prng_60_io_out_9,
    rand_exe_prng_60_io_out_8,rand_exe_lo_60}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_61 = {rand_exe_prng_61_io_out_7,rand_exe_prng_61_io_out_6,rand_exe_prng_61_io_out_5,
    rand_exe_prng_61_io_out_4,rand_exe_prng_61_io_out_3,rand_exe_prng_61_io_out_2,rand_exe_prng_61_io_out_1,
    rand_exe_prng_61_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_61 = {rand_exe_prng_61_io_out_15,rand_exe_prng_61_io_out_14,rand_exe_prng_61_io_out_13,
    rand_exe_prng_61_io_out_12,rand_exe_prng_61_io_out_11,rand_exe_prng_61_io_out_10,rand_exe_prng_61_io_out_9,
    rand_exe_prng_61_io_out_8,rand_exe_lo_61}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_62 = {rand_exe_prng_62_io_out_7,rand_exe_prng_62_io_out_6,rand_exe_prng_62_io_out_5,
    rand_exe_prng_62_io_out_4,rand_exe_prng_62_io_out_3,rand_exe_prng_62_io_out_2,rand_exe_prng_62_io_out_1,
    rand_exe_prng_62_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_62 = {rand_exe_prng_62_io_out_15,rand_exe_prng_62_io_out_14,rand_exe_prng_62_io_out_13,
    rand_exe_prng_62_io_out_12,rand_exe_prng_62_io_out_11,rand_exe_prng_62_io_out_10,rand_exe_prng_62_io_out_9,
    rand_exe_prng_62_io_out_8,rand_exe_lo_62}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_63 = {rand_exe_prng_63_io_out_7,rand_exe_prng_63_io_out_6,rand_exe_prng_63_io_out_5,
    rand_exe_prng_63_io_out_4,rand_exe_prng_63_io_out_3,rand_exe_prng_63_io_out_2,rand_exe_prng_63_io_out_1,
    rand_exe_prng_63_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_63 = {rand_exe_prng_63_io_out_15,rand_exe_prng_63_io_out_14,rand_exe_prng_63_io_out_13,
    rand_exe_prng_63_io_out_12,rand_exe_prng_63_io_out_11,rand_exe_prng_63_io_out_10,rand_exe_prng_63_io_out_9,
    rand_exe_prng_63_io_out_8,rand_exe_lo_63}; // @[PRNG.scala 86:17]
  MaxPeriodFibonacciLFSR rand_exe_prng ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_clock),
    .reset(rand_exe_prng_reset),
    .io_out_0(rand_exe_prng_io_out_0),
    .io_out_1(rand_exe_prng_io_out_1),
    .io_out_2(rand_exe_prng_io_out_2),
    .io_out_3(rand_exe_prng_io_out_3),
    .io_out_4(rand_exe_prng_io_out_4),
    .io_out_5(rand_exe_prng_io_out_5),
    .io_out_6(rand_exe_prng_io_out_6),
    .io_out_7(rand_exe_prng_io_out_7),
    .io_out_8(rand_exe_prng_io_out_8),
    .io_out_9(rand_exe_prng_io_out_9),
    .io_out_10(rand_exe_prng_io_out_10),
    .io_out_11(rand_exe_prng_io_out_11),
    .io_out_12(rand_exe_prng_io_out_12),
    .io_out_13(rand_exe_prng_io_out_13),
    .io_out_14(rand_exe_prng_io_out_14),
    .io_out_15(rand_exe_prng_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_1 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_1_clock),
    .reset(rand_exe_prng_1_reset),
    .io_out_0(rand_exe_prng_1_io_out_0),
    .io_out_1(rand_exe_prng_1_io_out_1),
    .io_out_2(rand_exe_prng_1_io_out_2),
    .io_out_3(rand_exe_prng_1_io_out_3),
    .io_out_4(rand_exe_prng_1_io_out_4),
    .io_out_5(rand_exe_prng_1_io_out_5),
    .io_out_6(rand_exe_prng_1_io_out_6),
    .io_out_7(rand_exe_prng_1_io_out_7),
    .io_out_8(rand_exe_prng_1_io_out_8),
    .io_out_9(rand_exe_prng_1_io_out_9),
    .io_out_10(rand_exe_prng_1_io_out_10),
    .io_out_11(rand_exe_prng_1_io_out_11),
    .io_out_12(rand_exe_prng_1_io_out_12),
    .io_out_13(rand_exe_prng_1_io_out_13),
    .io_out_14(rand_exe_prng_1_io_out_14),
    .io_out_15(rand_exe_prng_1_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_2 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_2_clock),
    .reset(rand_exe_prng_2_reset),
    .io_out_0(rand_exe_prng_2_io_out_0),
    .io_out_1(rand_exe_prng_2_io_out_1),
    .io_out_2(rand_exe_prng_2_io_out_2),
    .io_out_3(rand_exe_prng_2_io_out_3),
    .io_out_4(rand_exe_prng_2_io_out_4),
    .io_out_5(rand_exe_prng_2_io_out_5),
    .io_out_6(rand_exe_prng_2_io_out_6),
    .io_out_7(rand_exe_prng_2_io_out_7),
    .io_out_8(rand_exe_prng_2_io_out_8),
    .io_out_9(rand_exe_prng_2_io_out_9),
    .io_out_10(rand_exe_prng_2_io_out_10),
    .io_out_11(rand_exe_prng_2_io_out_11),
    .io_out_12(rand_exe_prng_2_io_out_12),
    .io_out_13(rand_exe_prng_2_io_out_13),
    .io_out_14(rand_exe_prng_2_io_out_14),
    .io_out_15(rand_exe_prng_2_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_3 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_3_clock),
    .reset(rand_exe_prng_3_reset),
    .io_out_0(rand_exe_prng_3_io_out_0),
    .io_out_1(rand_exe_prng_3_io_out_1),
    .io_out_2(rand_exe_prng_3_io_out_2),
    .io_out_3(rand_exe_prng_3_io_out_3),
    .io_out_4(rand_exe_prng_3_io_out_4),
    .io_out_5(rand_exe_prng_3_io_out_5),
    .io_out_6(rand_exe_prng_3_io_out_6),
    .io_out_7(rand_exe_prng_3_io_out_7),
    .io_out_8(rand_exe_prng_3_io_out_8),
    .io_out_9(rand_exe_prng_3_io_out_9),
    .io_out_10(rand_exe_prng_3_io_out_10),
    .io_out_11(rand_exe_prng_3_io_out_11),
    .io_out_12(rand_exe_prng_3_io_out_12),
    .io_out_13(rand_exe_prng_3_io_out_13),
    .io_out_14(rand_exe_prng_3_io_out_14),
    .io_out_15(rand_exe_prng_3_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_4 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_4_clock),
    .reset(rand_exe_prng_4_reset),
    .io_out_0(rand_exe_prng_4_io_out_0),
    .io_out_1(rand_exe_prng_4_io_out_1),
    .io_out_2(rand_exe_prng_4_io_out_2),
    .io_out_3(rand_exe_prng_4_io_out_3),
    .io_out_4(rand_exe_prng_4_io_out_4),
    .io_out_5(rand_exe_prng_4_io_out_5),
    .io_out_6(rand_exe_prng_4_io_out_6),
    .io_out_7(rand_exe_prng_4_io_out_7),
    .io_out_8(rand_exe_prng_4_io_out_8),
    .io_out_9(rand_exe_prng_4_io_out_9),
    .io_out_10(rand_exe_prng_4_io_out_10),
    .io_out_11(rand_exe_prng_4_io_out_11),
    .io_out_12(rand_exe_prng_4_io_out_12),
    .io_out_13(rand_exe_prng_4_io_out_13),
    .io_out_14(rand_exe_prng_4_io_out_14),
    .io_out_15(rand_exe_prng_4_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_5 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_5_clock),
    .reset(rand_exe_prng_5_reset),
    .io_out_0(rand_exe_prng_5_io_out_0),
    .io_out_1(rand_exe_prng_5_io_out_1),
    .io_out_2(rand_exe_prng_5_io_out_2),
    .io_out_3(rand_exe_prng_5_io_out_3),
    .io_out_4(rand_exe_prng_5_io_out_4),
    .io_out_5(rand_exe_prng_5_io_out_5),
    .io_out_6(rand_exe_prng_5_io_out_6),
    .io_out_7(rand_exe_prng_5_io_out_7),
    .io_out_8(rand_exe_prng_5_io_out_8),
    .io_out_9(rand_exe_prng_5_io_out_9),
    .io_out_10(rand_exe_prng_5_io_out_10),
    .io_out_11(rand_exe_prng_5_io_out_11),
    .io_out_12(rand_exe_prng_5_io_out_12),
    .io_out_13(rand_exe_prng_5_io_out_13),
    .io_out_14(rand_exe_prng_5_io_out_14),
    .io_out_15(rand_exe_prng_5_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_6 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_6_clock),
    .reset(rand_exe_prng_6_reset),
    .io_out_0(rand_exe_prng_6_io_out_0),
    .io_out_1(rand_exe_prng_6_io_out_1),
    .io_out_2(rand_exe_prng_6_io_out_2),
    .io_out_3(rand_exe_prng_6_io_out_3),
    .io_out_4(rand_exe_prng_6_io_out_4),
    .io_out_5(rand_exe_prng_6_io_out_5),
    .io_out_6(rand_exe_prng_6_io_out_6),
    .io_out_7(rand_exe_prng_6_io_out_7),
    .io_out_8(rand_exe_prng_6_io_out_8),
    .io_out_9(rand_exe_prng_6_io_out_9),
    .io_out_10(rand_exe_prng_6_io_out_10),
    .io_out_11(rand_exe_prng_6_io_out_11),
    .io_out_12(rand_exe_prng_6_io_out_12),
    .io_out_13(rand_exe_prng_6_io_out_13),
    .io_out_14(rand_exe_prng_6_io_out_14),
    .io_out_15(rand_exe_prng_6_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_7 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_7_clock),
    .reset(rand_exe_prng_7_reset),
    .io_out_0(rand_exe_prng_7_io_out_0),
    .io_out_1(rand_exe_prng_7_io_out_1),
    .io_out_2(rand_exe_prng_7_io_out_2),
    .io_out_3(rand_exe_prng_7_io_out_3),
    .io_out_4(rand_exe_prng_7_io_out_4),
    .io_out_5(rand_exe_prng_7_io_out_5),
    .io_out_6(rand_exe_prng_7_io_out_6),
    .io_out_7(rand_exe_prng_7_io_out_7),
    .io_out_8(rand_exe_prng_7_io_out_8),
    .io_out_9(rand_exe_prng_7_io_out_9),
    .io_out_10(rand_exe_prng_7_io_out_10),
    .io_out_11(rand_exe_prng_7_io_out_11),
    .io_out_12(rand_exe_prng_7_io_out_12),
    .io_out_13(rand_exe_prng_7_io_out_13),
    .io_out_14(rand_exe_prng_7_io_out_14),
    .io_out_15(rand_exe_prng_7_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_8 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_8_clock),
    .reset(rand_exe_prng_8_reset),
    .io_out_0(rand_exe_prng_8_io_out_0),
    .io_out_1(rand_exe_prng_8_io_out_1),
    .io_out_2(rand_exe_prng_8_io_out_2),
    .io_out_3(rand_exe_prng_8_io_out_3),
    .io_out_4(rand_exe_prng_8_io_out_4),
    .io_out_5(rand_exe_prng_8_io_out_5),
    .io_out_6(rand_exe_prng_8_io_out_6),
    .io_out_7(rand_exe_prng_8_io_out_7),
    .io_out_8(rand_exe_prng_8_io_out_8),
    .io_out_9(rand_exe_prng_8_io_out_9),
    .io_out_10(rand_exe_prng_8_io_out_10),
    .io_out_11(rand_exe_prng_8_io_out_11),
    .io_out_12(rand_exe_prng_8_io_out_12),
    .io_out_13(rand_exe_prng_8_io_out_13),
    .io_out_14(rand_exe_prng_8_io_out_14),
    .io_out_15(rand_exe_prng_8_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_9 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_9_clock),
    .reset(rand_exe_prng_9_reset),
    .io_out_0(rand_exe_prng_9_io_out_0),
    .io_out_1(rand_exe_prng_9_io_out_1),
    .io_out_2(rand_exe_prng_9_io_out_2),
    .io_out_3(rand_exe_prng_9_io_out_3),
    .io_out_4(rand_exe_prng_9_io_out_4),
    .io_out_5(rand_exe_prng_9_io_out_5),
    .io_out_6(rand_exe_prng_9_io_out_6),
    .io_out_7(rand_exe_prng_9_io_out_7),
    .io_out_8(rand_exe_prng_9_io_out_8),
    .io_out_9(rand_exe_prng_9_io_out_9),
    .io_out_10(rand_exe_prng_9_io_out_10),
    .io_out_11(rand_exe_prng_9_io_out_11),
    .io_out_12(rand_exe_prng_9_io_out_12),
    .io_out_13(rand_exe_prng_9_io_out_13),
    .io_out_14(rand_exe_prng_9_io_out_14),
    .io_out_15(rand_exe_prng_9_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_10 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_10_clock),
    .reset(rand_exe_prng_10_reset),
    .io_out_0(rand_exe_prng_10_io_out_0),
    .io_out_1(rand_exe_prng_10_io_out_1),
    .io_out_2(rand_exe_prng_10_io_out_2),
    .io_out_3(rand_exe_prng_10_io_out_3),
    .io_out_4(rand_exe_prng_10_io_out_4),
    .io_out_5(rand_exe_prng_10_io_out_5),
    .io_out_6(rand_exe_prng_10_io_out_6),
    .io_out_7(rand_exe_prng_10_io_out_7),
    .io_out_8(rand_exe_prng_10_io_out_8),
    .io_out_9(rand_exe_prng_10_io_out_9),
    .io_out_10(rand_exe_prng_10_io_out_10),
    .io_out_11(rand_exe_prng_10_io_out_11),
    .io_out_12(rand_exe_prng_10_io_out_12),
    .io_out_13(rand_exe_prng_10_io_out_13),
    .io_out_14(rand_exe_prng_10_io_out_14),
    .io_out_15(rand_exe_prng_10_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_11 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_11_clock),
    .reset(rand_exe_prng_11_reset),
    .io_out_0(rand_exe_prng_11_io_out_0),
    .io_out_1(rand_exe_prng_11_io_out_1),
    .io_out_2(rand_exe_prng_11_io_out_2),
    .io_out_3(rand_exe_prng_11_io_out_3),
    .io_out_4(rand_exe_prng_11_io_out_4),
    .io_out_5(rand_exe_prng_11_io_out_5),
    .io_out_6(rand_exe_prng_11_io_out_6),
    .io_out_7(rand_exe_prng_11_io_out_7),
    .io_out_8(rand_exe_prng_11_io_out_8),
    .io_out_9(rand_exe_prng_11_io_out_9),
    .io_out_10(rand_exe_prng_11_io_out_10),
    .io_out_11(rand_exe_prng_11_io_out_11),
    .io_out_12(rand_exe_prng_11_io_out_12),
    .io_out_13(rand_exe_prng_11_io_out_13),
    .io_out_14(rand_exe_prng_11_io_out_14),
    .io_out_15(rand_exe_prng_11_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_12 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_12_clock),
    .reset(rand_exe_prng_12_reset),
    .io_out_0(rand_exe_prng_12_io_out_0),
    .io_out_1(rand_exe_prng_12_io_out_1),
    .io_out_2(rand_exe_prng_12_io_out_2),
    .io_out_3(rand_exe_prng_12_io_out_3),
    .io_out_4(rand_exe_prng_12_io_out_4),
    .io_out_5(rand_exe_prng_12_io_out_5),
    .io_out_6(rand_exe_prng_12_io_out_6),
    .io_out_7(rand_exe_prng_12_io_out_7),
    .io_out_8(rand_exe_prng_12_io_out_8),
    .io_out_9(rand_exe_prng_12_io_out_9),
    .io_out_10(rand_exe_prng_12_io_out_10),
    .io_out_11(rand_exe_prng_12_io_out_11),
    .io_out_12(rand_exe_prng_12_io_out_12),
    .io_out_13(rand_exe_prng_12_io_out_13),
    .io_out_14(rand_exe_prng_12_io_out_14),
    .io_out_15(rand_exe_prng_12_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_13 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_13_clock),
    .reset(rand_exe_prng_13_reset),
    .io_out_0(rand_exe_prng_13_io_out_0),
    .io_out_1(rand_exe_prng_13_io_out_1),
    .io_out_2(rand_exe_prng_13_io_out_2),
    .io_out_3(rand_exe_prng_13_io_out_3),
    .io_out_4(rand_exe_prng_13_io_out_4),
    .io_out_5(rand_exe_prng_13_io_out_5),
    .io_out_6(rand_exe_prng_13_io_out_6),
    .io_out_7(rand_exe_prng_13_io_out_7),
    .io_out_8(rand_exe_prng_13_io_out_8),
    .io_out_9(rand_exe_prng_13_io_out_9),
    .io_out_10(rand_exe_prng_13_io_out_10),
    .io_out_11(rand_exe_prng_13_io_out_11),
    .io_out_12(rand_exe_prng_13_io_out_12),
    .io_out_13(rand_exe_prng_13_io_out_13),
    .io_out_14(rand_exe_prng_13_io_out_14),
    .io_out_15(rand_exe_prng_13_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_14 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_14_clock),
    .reset(rand_exe_prng_14_reset),
    .io_out_0(rand_exe_prng_14_io_out_0),
    .io_out_1(rand_exe_prng_14_io_out_1),
    .io_out_2(rand_exe_prng_14_io_out_2),
    .io_out_3(rand_exe_prng_14_io_out_3),
    .io_out_4(rand_exe_prng_14_io_out_4),
    .io_out_5(rand_exe_prng_14_io_out_5),
    .io_out_6(rand_exe_prng_14_io_out_6),
    .io_out_7(rand_exe_prng_14_io_out_7),
    .io_out_8(rand_exe_prng_14_io_out_8),
    .io_out_9(rand_exe_prng_14_io_out_9),
    .io_out_10(rand_exe_prng_14_io_out_10),
    .io_out_11(rand_exe_prng_14_io_out_11),
    .io_out_12(rand_exe_prng_14_io_out_12),
    .io_out_13(rand_exe_prng_14_io_out_13),
    .io_out_14(rand_exe_prng_14_io_out_14),
    .io_out_15(rand_exe_prng_14_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_15 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_15_clock),
    .reset(rand_exe_prng_15_reset),
    .io_out_0(rand_exe_prng_15_io_out_0),
    .io_out_1(rand_exe_prng_15_io_out_1),
    .io_out_2(rand_exe_prng_15_io_out_2),
    .io_out_3(rand_exe_prng_15_io_out_3),
    .io_out_4(rand_exe_prng_15_io_out_4),
    .io_out_5(rand_exe_prng_15_io_out_5),
    .io_out_6(rand_exe_prng_15_io_out_6),
    .io_out_7(rand_exe_prng_15_io_out_7),
    .io_out_8(rand_exe_prng_15_io_out_8),
    .io_out_9(rand_exe_prng_15_io_out_9),
    .io_out_10(rand_exe_prng_15_io_out_10),
    .io_out_11(rand_exe_prng_15_io_out_11),
    .io_out_12(rand_exe_prng_15_io_out_12),
    .io_out_13(rand_exe_prng_15_io_out_13),
    .io_out_14(rand_exe_prng_15_io_out_14),
    .io_out_15(rand_exe_prng_15_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_16 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_16_clock),
    .reset(rand_exe_prng_16_reset),
    .io_out_0(rand_exe_prng_16_io_out_0),
    .io_out_1(rand_exe_prng_16_io_out_1),
    .io_out_2(rand_exe_prng_16_io_out_2),
    .io_out_3(rand_exe_prng_16_io_out_3),
    .io_out_4(rand_exe_prng_16_io_out_4),
    .io_out_5(rand_exe_prng_16_io_out_5),
    .io_out_6(rand_exe_prng_16_io_out_6),
    .io_out_7(rand_exe_prng_16_io_out_7),
    .io_out_8(rand_exe_prng_16_io_out_8),
    .io_out_9(rand_exe_prng_16_io_out_9),
    .io_out_10(rand_exe_prng_16_io_out_10),
    .io_out_11(rand_exe_prng_16_io_out_11),
    .io_out_12(rand_exe_prng_16_io_out_12),
    .io_out_13(rand_exe_prng_16_io_out_13),
    .io_out_14(rand_exe_prng_16_io_out_14),
    .io_out_15(rand_exe_prng_16_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_17 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_17_clock),
    .reset(rand_exe_prng_17_reset),
    .io_out_0(rand_exe_prng_17_io_out_0),
    .io_out_1(rand_exe_prng_17_io_out_1),
    .io_out_2(rand_exe_prng_17_io_out_2),
    .io_out_3(rand_exe_prng_17_io_out_3),
    .io_out_4(rand_exe_prng_17_io_out_4),
    .io_out_5(rand_exe_prng_17_io_out_5),
    .io_out_6(rand_exe_prng_17_io_out_6),
    .io_out_7(rand_exe_prng_17_io_out_7),
    .io_out_8(rand_exe_prng_17_io_out_8),
    .io_out_9(rand_exe_prng_17_io_out_9),
    .io_out_10(rand_exe_prng_17_io_out_10),
    .io_out_11(rand_exe_prng_17_io_out_11),
    .io_out_12(rand_exe_prng_17_io_out_12),
    .io_out_13(rand_exe_prng_17_io_out_13),
    .io_out_14(rand_exe_prng_17_io_out_14),
    .io_out_15(rand_exe_prng_17_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_18 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_18_clock),
    .reset(rand_exe_prng_18_reset),
    .io_out_0(rand_exe_prng_18_io_out_0),
    .io_out_1(rand_exe_prng_18_io_out_1),
    .io_out_2(rand_exe_prng_18_io_out_2),
    .io_out_3(rand_exe_prng_18_io_out_3),
    .io_out_4(rand_exe_prng_18_io_out_4),
    .io_out_5(rand_exe_prng_18_io_out_5),
    .io_out_6(rand_exe_prng_18_io_out_6),
    .io_out_7(rand_exe_prng_18_io_out_7),
    .io_out_8(rand_exe_prng_18_io_out_8),
    .io_out_9(rand_exe_prng_18_io_out_9),
    .io_out_10(rand_exe_prng_18_io_out_10),
    .io_out_11(rand_exe_prng_18_io_out_11),
    .io_out_12(rand_exe_prng_18_io_out_12),
    .io_out_13(rand_exe_prng_18_io_out_13),
    .io_out_14(rand_exe_prng_18_io_out_14),
    .io_out_15(rand_exe_prng_18_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_19 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_19_clock),
    .reset(rand_exe_prng_19_reset),
    .io_out_0(rand_exe_prng_19_io_out_0),
    .io_out_1(rand_exe_prng_19_io_out_1),
    .io_out_2(rand_exe_prng_19_io_out_2),
    .io_out_3(rand_exe_prng_19_io_out_3),
    .io_out_4(rand_exe_prng_19_io_out_4),
    .io_out_5(rand_exe_prng_19_io_out_5),
    .io_out_6(rand_exe_prng_19_io_out_6),
    .io_out_7(rand_exe_prng_19_io_out_7),
    .io_out_8(rand_exe_prng_19_io_out_8),
    .io_out_9(rand_exe_prng_19_io_out_9),
    .io_out_10(rand_exe_prng_19_io_out_10),
    .io_out_11(rand_exe_prng_19_io_out_11),
    .io_out_12(rand_exe_prng_19_io_out_12),
    .io_out_13(rand_exe_prng_19_io_out_13),
    .io_out_14(rand_exe_prng_19_io_out_14),
    .io_out_15(rand_exe_prng_19_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_20 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_20_clock),
    .reset(rand_exe_prng_20_reset),
    .io_out_0(rand_exe_prng_20_io_out_0),
    .io_out_1(rand_exe_prng_20_io_out_1),
    .io_out_2(rand_exe_prng_20_io_out_2),
    .io_out_3(rand_exe_prng_20_io_out_3),
    .io_out_4(rand_exe_prng_20_io_out_4),
    .io_out_5(rand_exe_prng_20_io_out_5),
    .io_out_6(rand_exe_prng_20_io_out_6),
    .io_out_7(rand_exe_prng_20_io_out_7),
    .io_out_8(rand_exe_prng_20_io_out_8),
    .io_out_9(rand_exe_prng_20_io_out_9),
    .io_out_10(rand_exe_prng_20_io_out_10),
    .io_out_11(rand_exe_prng_20_io_out_11),
    .io_out_12(rand_exe_prng_20_io_out_12),
    .io_out_13(rand_exe_prng_20_io_out_13),
    .io_out_14(rand_exe_prng_20_io_out_14),
    .io_out_15(rand_exe_prng_20_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_21 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_21_clock),
    .reset(rand_exe_prng_21_reset),
    .io_out_0(rand_exe_prng_21_io_out_0),
    .io_out_1(rand_exe_prng_21_io_out_1),
    .io_out_2(rand_exe_prng_21_io_out_2),
    .io_out_3(rand_exe_prng_21_io_out_3),
    .io_out_4(rand_exe_prng_21_io_out_4),
    .io_out_5(rand_exe_prng_21_io_out_5),
    .io_out_6(rand_exe_prng_21_io_out_6),
    .io_out_7(rand_exe_prng_21_io_out_7),
    .io_out_8(rand_exe_prng_21_io_out_8),
    .io_out_9(rand_exe_prng_21_io_out_9),
    .io_out_10(rand_exe_prng_21_io_out_10),
    .io_out_11(rand_exe_prng_21_io_out_11),
    .io_out_12(rand_exe_prng_21_io_out_12),
    .io_out_13(rand_exe_prng_21_io_out_13),
    .io_out_14(rand_exe_prng_21_io_out_14),
    .io_out_15(rand_exe_prng_21_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_22 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_22_clock),
    .reset(rand_exe_prng_22_reset),
    .io_out_0(rand_exe_prng_22_io_out_0),
    .io_out_1(rand_exe_prng_22_io_out_1),
    .io_out_2(rand_exe_prng_22_io_out_2),
    .io_out_3(rand_exe_prng_22_io_out_3),
    .io_out_4(rand_exe_prng_22_io_out_4),
    .io_out_5(rand_exe_prng_22_io_out_5),
    .io_out_6(rand_exe_prng_22_io_out_6),
    .io_out_7(rand_exe_prng_22_io_out_7),
    .io_out_8(rand_exe_prng_22_io_out_8),
    .io_out_9(rand_exe_prng_22_io_out_9),
    .io_out_10(rand_exe_prng_22_io_out_10),
    .io_out_11(rand_exe_prng_22_io_out_11),
    .io_out_12(rand_exe_prng_22_io_out_12),
    .io_out_13(rand_exe_prng_22_io_out_13),
    .io_out_14(rand_exe_prng_22_io_out_14),
    .io_out_15(rand_exe_prng_22_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_23 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_23_clock),
    .reset(rand_exe_prng_23_reset),
    .io_out_0(rand_exe_prng_23_io_out_0),
    .io_out_1(rand_exe_prng_23_io_out_1),
    .io_out_2(rand_exe_prng_23_io_out_2),
    .io_out_3(rand_exe_prng_23_io_out_3),
    .io_out_4(rand_exe_prng_23_io_out_4),
    .io_out_5(rand_exe_prng_23_io_out_5),
    .io_out_6(rand_exe_prng_23_io_out_6),
    .io_out_7(rand_exe_prng_23_io_out_7),
    .io_out_8(rand_exe_prng_23_io_out_8),
    .io_out_9(rand_exe_prng_23_io_out_9),
    .io_out_10(rand_exe_prng_23_io_out_10),
    .io_out_11(rand_exe_prng_23_io_out_11),
    .io_out_12(rand_exe_prng_23_io_out_12),
    .io_out_13(rand_exe_prng_23_io_out_13),
    .io_out_14(rand_exe_prng_23_io_out_14),
    .io_out_15(rand_exe_prng_23_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_24 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_24_clock),
    .reset(rand_exe_prng_24_reset),
    .io_out_0(rand_exe_prng_24_io_out_0),
    .io_out_1(rand_exe_prng_24_io_out_1),
    .io_out_2(rand_exe_prng_24_io_out_2),
    .io_out_3(rand_exe_prng_24_io_out_3),
    .io_out_4(rand_exe_prng_24_io_out_4),
    .io_out_5(rand_exe_prng_24_io_out_5),
    .io_out_6(rand_exe_prng_24_io_out_6),
    .io_out_7(rand_exe_prng_24_io_out_7),
    .io_out_8(rand_exe_prng_24_io_out_8),
    .io_out_9(rand_exe_prng_24_io_out_9),
    .io_out_10(rand_exe_prng_24_io_out_10),
    .io_out_11(rand_exe_prng_24_io_out_11),
    .io_out_12(rand_exe_prng_24_io_out_12),
    .io_out_13(rand_exe_prng_24_io_out_13),
    .io_out_14(rand_exe_prng_24_io_out_14),
    .io_out_15(rand_exe_prng_24_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_25 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_25_clock),
    .reset(rand_exe_prng_25_reset),
    .io_out_0(rand_exe_prng_25_io_out_0),
    .io_out_1(rand_exe_prng_25_io_out_1),
    .io_out_2(rand_exe_prng_25_io_out_2),
    .io_out_3(rand_exe_prng_25_io_out_3),
    .io_out_4(rand_exe_prng_25_io_out_4),
    .io_out_5(rand_exe_prng_25_io_out_5),
    .io_out_6(rand_exe_prng_25_io_out_6),
    .io_out_7(rand_exe_prng_25_io_out_7),
    .io_out_8(rand_exe_prng_25_io_out_8),
    .io_out_9(rand_exe_prng_25_io_out_9),
    .io_out_10(rand_exe_prng_25_io_out_10),
    .io_out_11(rand_exe_prng_25_io_out_11),
    .io_out_12(rand_exe_prng_25_io_out_12),
    .io_out_13(rand_exe_prng_25_io_out_13),
    .io_out_14(rand_exe_prng_25_io_out_14),
    .io_out_15(rand_exe_prng_25_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_26 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_26_clock),
    .reset(rand_exe_prng_26_reset),
    .io_out_0(rand_exe_prng_26_io_out_0),
    .io_out_1(rand_exe_prng_26_io_out_1),
    .io_out_2(rand_exe_prng_26_io_out_2),
    .io_out_3(rand_exe_prng_26_io_out_3),
    .io_out_4(rand_exe_prng_26_io_out_4),
    .io_out_5(rand_exe_prng_26_io_out_5),
    .io_out_6(rand_exe_prng_26_io_out_6),
    .io_out_7(rand_exe_prng_26_io_out_7),
    .io_out_8(rand_exe_prng_26_io_out_8),
    .io_out_9(rand_exe_prng_26_io_out_9),
    .io_out_10(rand_exe_prng_26_io_out_10),
    .io_out_11(rand_exe_prng_26_io_out_11),
    .io_out_12(rand_exe_prng_26_io_out_12),
    .io_out_13(rand_exe_prng_26_io_out_13),
    .io_out_14(rand_exe_prng_26_io_out_14),
    .io_out_15(rand_exe_prng_26_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_27 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_27_clock),
    .reset(rand_exe_prng_27_reset),
    .io_out_0(rand_exe_prng_27_io_out_0),
    .io_out_1(rand_exe_prng_27_io_out_1),
    .io_out_2(rand_exe_prng_27_io_out_2),
    .io_out_3(rand_exe_prng_27_io_out_3),
    .io_out_4(rand_exe_prng_27_io_out_4),
    .io_out_5(rand_exe_prng_27_io_out_5),
    .io_out_6(rand_exe_prng_27_io_out_6),
    .io_out_7(rand_exe_prng_27_io_out_7),
    .io_out_8(rand_exe_prng_27_io_out_8),
    .io_out_9(rand_exe_prng_27_io_out_9),
    .io_out_10(rand_exe_prng_27_io_out_10),
    .io_out_11(rand_exe_prng_27_io_out_11),
    .io_out_12(rand_exe_prng_27_io_out_12),
    .io_out_13(rand_exe_prng_27_io_out_13),
    .io_out_14(rand_exe_prng_27_io_out_14),
    .io_out_15(rand_exe_prng_27_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_28 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_28_clock),
    .reset(rand_exe_prng_28_reset),
    .io_out_0(rand_exe_prng_28_io_out_0),
    .io_out_1(rand_exe_prng_28_io_out_1),
    .io_out_2(rand_exe_prng_28_io_out_2),
    .io_out_3(rand_exe_prng_28_io_out_3),
    .io_out_4(rand_exe_prng_28_io_out_4),
    .io_out_5(rand_exe_prng_28_io_out_5),
    .io_out_6(rand_exe_prng_28_io_out_6),
    .io_out_7(rand_exe_prng_28_io_out_7),
    .io_out_8(rand_exe_prng_28_io_out_8),
    .io_out_9(rand_exe_prng_28_io_out_9),
    .io_out_10(rand_exe_prng_28_io_out_10),
    .io_out_11(rand_exe_prng_28_io_out_11),
    .io_out_12(rand_exe_prng_28_io_out_12),
    .io_out_13(rand_exe_prng_28_io_out_13),
    .io_out_14(rand_exe_prng_28_io_out_14),
    .io_out_15(rand_exe_prng_28_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_29 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_29_clock),
    .reset(rand_exe_prng_29_reset),
    .io_out_0(rand_exe_prng_29_io_out_0),
    .io_out_1(rand_exe_prng_29_io_out_1),
    .io_out_2(rand_exe_prng_29_io_out_2),
    .io_out_3(rand_exe_prng_29_io_out_3),
    .io_out_4(rand_exe_prng_29_io_out_4),
    .io_out_5(rand_exe_prng_29_io_out_5),
    .io_out_6(rand_exe_prng_29_io_out_6),
    .io_out_7(rand_exe_prng_29_io_out_7),
    .io_out_8(rand_exe_prng_29_io_out_8),
    .io_out_9(rand_exe_prng_29_io_out_9),
    .io_out_10(rand_exe_prng_29_io_out_10),
    .io_out_11(rand_exe_prng_29_io_out_11),
    .io_out_12(rand_exe_prng_29_io_out_12),
    .io_out_13(rand_exe_prng_29_io_out_13),
    .io_out_14(rand_exe_prng_29_io_out_14),
    .io_out_15(rand_exe_prng_29_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_30 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_30_clock),
    .reset(rand_exe_prng_30_reset),
    .io_out_0(rand_exe_prng_30_io_out_0),
    .io_out_1(rand_exe_prng_30_io_out_1),
    .io_out_2(rand_exe_prng_30_io_out_2),
    .io_out_3(rand_exe_prng_30_io_out_3),
    .io_out_4(rand_exe_prng_30_io_out_4),
    .io_out_5(rand_exe_prng_30_io_out_5),
    .io_out_6(rand_exe_prng_30_io_out_6),
    .io_out_7(rand_exe_prng_30_io_out_7),
    .io_out_8(rand_exe_prng_30_io_out_8),
    .io_out_9(rand_exe_prng_30_io_out_9),
    .io_out_10(rand_exe_prng_30_io_out_10),
    .io_out_11(rand_exe_prng_30_io_out_11),
    .io_out_12(rand_exe_prng_30_io_out_12),
    .io_out_13(rand_exe_prng_30_io_out_13),
    .io_out_14(rand_exe_prng_30_io_out_14),
    .io_out_15(rand_exe_prng_30_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_31 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_31_clock),
    .reset(rand_exe_prng_31_reset),
    .io_out_0(rand_exe_prng_31_io_out_0),
    .io_out_1(rand_exe_prng_31_io_out_1),
    .io_out_2(rand_exe_prng_31_io_out_2),
    .io_out_3(rand_exe_prng_31_io_out_3),
    .io_out_4(rand_exe_prng_31_io_out_4),
    .io_out_5(rand_exe_prng_31_io_out_5),
    .io_out_6(rand_exe_prng_31_io_out_6),
    .io_out_7(rand_exe_prng_31_io_out_7),
    .io_out_8(rand_exe_prng_31_io_out_8),
    .io_out_9(rand_exe_prng_31_io_out_9),
    .io_out_10(rand_exe_prng_31_io_out_10),
    .io_out_11(rand_exe_prng_31_io_out_11),
    .io_out_12(rand_exe_prng_31_io_out_12),
    .io_out_13(rand_exe_prng_31_io_out_13),
    .io_out_14(rand_exe_prng_31_io_out_14),
    .io_out_15(rand_exe_prng_31_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_32 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_32_clock),
    .reset(rand_exe_prng_32_reset),
    .io_out_0(rand_exe_prng_32_io_out_0),
    .io_out_1(rand_exe_prng_32_io_out_1),
    .io_out_2(rand_exe_prng_32_io_out_2),
    .io_out_3(rand_exe_prng_32_io_out_3),
    .io_out_4(rand_exe_prng_32_io_out_4),
    .io_out_5(rand_exe_prng_32_io_out_5),
    .io_out_6(rand_exe_prng_32_io_out_6),
    .io_out_7(rand_exe_prng_32_io_out_7),
    .io_out_8(rand_exe_prng_32_io_out_8),
    .io_out_9(rand_exe_prng_32_io_out_9),
    .io_out_10(rand_exe_prng_32_io_out_10),
    .io_out_11(rand_exe_prng_32_io_out_11),
    .io_out_12(rand_exe_prng_32_io_out_12),
    .io_out_13(rand_exe_prng_32_io_out_13),
    .io_out_14(rand_exe_prng_32_io_out_14),
    .io_out_15(rand_exe_prng_32_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_33 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_33_clock),
    .reset(rand_exe_prng_33_reset),
    .io_out_0(rand_exe_prng_33_io_out_0),
    .io_out_1(rand_exe_prng_33_io_out_1),
    .io_out_2(rand_exe_prng_33_io_out_2),
    .io_out_3(rand_exe_prng_33_io_out_3),
    .io_out_4(rand_exe_prng_33_io_out_4),
    .io_out_5(rand_exe_prng_33_io_out_5),
    .io_out_6(rand_exe_prng_33_io_out_6),
    .io_out_7(rand_exe_prng_33_io_out_7),
    .io_out_8(rand_exe_prng_33_io_out_8),
    .io_out_9(rand_exe_prng_33_io_out_9),
    .io_out_10(rand_exe_prng_33_io_out_10),
    .io_out_11(rand_exe_prng_33_io_out_11),
    .io_out_12(rand_exe_prng_33_io_out_12),
    .io_out_13(rand_exe_prng_33_io_out_13),
    .io_out_14(rand_exe_prng_33_io_out_14),
    .io_out_15(rand_exe_prng_33_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_34 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_34_clock),
    .reset(rand_exe_prng_34_reset),
    .io_out_0(rand_exe_prng_34_io_out_0),
    .io_out_1(rand_exe_prng_34_io_out_1),
    .io_out_2(rand_exe_prng_34_io_out_2),
    .io_out_3(rand_exe_prng_34_io_out_3),
    .io_out_4(rand_exe_prng_34_io_out_4),
    .io_out_5(rand_exe_prng_34_io_out_5),
    .io_out_6(rand_exe_prng_34_io_out_6),
    .io_out_7(rand_exe_prng_34_io_out_7),
    .io_out_8(rand_exe_prng_34_io_out_8),
    .io_out_9(rand_exe_prng_34_io_out_9),
    .io_out_10(rand_exe_prng_34_io_out_10),
    .io_out_11(rand_exe_prng_34_io_out_11),
    .io_out_12(rand_exe_prng_34_io_out_12),
    .io_out_13(rand_exe_prng_34_io_out_13),
    .io_out_14(rand_exe_prng_34_io_out_14),
    .io_out_15(rand_exe_prng_34_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_35 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_35_clock),
    .reset(rand_exe_prng_35_reset),
    .io_out_0(rand_exe_prng_35_io_out_0),
    .io_out_1(rand_exe_prng_35_io_out_1),
    .io_out_2(rand_exe_prng_35_io_out_2),
    .io_out_3(rand_exe_prng_35_io_out_3),
    .io_out_4(rand_exe_prng_35_io_out_4),
    .io_out_5(rand_exe_prng_35_io_out_5),
    .io_out_6(rand_exe_prng_35_io_out_6),
    .io_out_7(rand_exe_prng_35_io_out_7),
    .io_out_8(rand_exe_prng_35_io_out_8),
    .io_out_9(rand_exe_prng_35_io_out_9),
    .io_out_10(rand_exe_prng_35_io_out_10),
    .io_out_11(rand_exe_prng_35_io_out_11),
    .io_out_12(rand_exe_prng_35_io_out_12),
    .io_out_13(rand_exe_prng_35_io_out_13),
    .io_out_14(rand_exe_prng_35_io_out_14),
    .io_out_15(rand_exe_prng_35_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_36 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_36_clock),
    .reset(rand_exe_prng_36_reset),
    .io_out_0(rand_exe_prng_36_io_out_0),
    .io_out_1(rand_exe_prng_36_io_out_1),
    .io_out_2(rand_exe_prng_36_io_out_2),
    .io_out_3(rand_exe_prng_36_io_out_3),
    .io_out_4(rand_exe_prng_36_io_out_4),
    .io_out_5(rand_exe_prng_36_io_out_5),
    .io_out_6(rand_exe_prng_36_io_out_6),
    .io_out_7(rand_exe_prng_36_io_out_7),
    .io_out_8(rand_exe_prng_36_io_out_8),
    .io_out_9(rand_exe_prng_36_io_out_9),
    .io_out_10(rand_exe_prng_36_io_out_10),
    .io_out_11(rand_exe_prng_36_io_out_11),
    .io_out_12(rand_exe_prng_36_io_out_12),
    .io_out_13(rand_exe_prng_36_io_out_13),
    .io_out_14(rand_exe_prng_36_io_out_14),
    .io_out_15(rand_exe_prng_36_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_37 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_37_clock),
    .reset(rand_exe_prng_37_reset),
    .io_out_0(rand_exe_prng_37_io_out_0),
    .io_out_1(rand_exe_prng_37_io_out_1),
    .io_out_2(rand_exe_prng_37_io_out_2),
    .io_out_3(rand_exe_prng_37_io_out_3),
    .io_out_4(rand_exe_prng_37_io_out_4),
    .io_out_5(rand_exe_prng_37_io_out_5),
    .io_out_6(rand_exe_prng_37_io_out_6),
    .io_out_7(rand_exe_prng_37_io_out_7),
    .io_out_8(rand_exe_prng_37_io_out_8),
    .io_out_9(rand_exe_prng_37_io_out_9),
    .io_out_10(rand_exe_prng_37_io_out_10),
    .io_out_11(rand_exe_prng_37_io_out_11),
    .io_out_12(rand_exe_prng_37_io_out_12),
    .io_out_13(rand_exe_prng_37_io_out_13),
    .io_out_14(rand_exe_prng_37_io_out_14),
    .io_out_15(rand_exe_prng_37_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_38 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_38_clock),
    .reset(rand_exe_prng_38_reset),
    .io_out_0(rand_exe_prng_38_io_out_0),
    .io_out_1(rand_exe_prng_38_io_out_1),
    .io_out_2(rand_exe_prng_38_io_out_2),
    .io_out_3(rand_exe_prng_38_io_out_3),
    .io_out_4(rand_exe_prng_38_io_out_4),
    .io_out_5(rand_exe_prng_38_io_out_5),
    .io_out_6(rand_exe_prng_38_io_out_6),
    .io_out_7(rand_exe_prng_38_io_out_7),
    .io_out_8(rand_exe_prng_38_io_out_8),
    .io_out_9(rand_exe_prng_38_io_out_9),
    .io_out_10(rand_exe_prng_38_io_out_10),
    .io_out_11(rand_exe_prng_38_io_out_11),
    .io_out_12(rand_exe_prng_38_io_out_12),
    .io_out_13(rand_exe_prng_38_io_out_13),
    .io_out_14(rand_exe_prng_38_io_out_14),
    .io_out_15(rand_exe_prng_38_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_39 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_39_clock),
    .reset(rand_exe_prng_39_reset),
    .io_out_0(rand_exe_prng_39_io_out_0),
    .io_out_1(rand_exe_prng_39_io_out_1),
    .io_out_2(rand_exe_prng_39_io_out_2),
    .io_out_3(rand_exe_prng_39_io_out_3),
    .io_out_4(rand_exe_prng_39_io_out_4),
    .io_out_5(rand_exe_prng_39_io_out_5),
    .io_out_6(rand_exe_prng_39_io_out_6),
    .io_out_7(rand_exe_prng_39_io_out_7),
    .io_out_8(rand_exe_prng_39_io_out_8),
    .io_out_9(rand_exe_prng_39_io_out_9),
    .io_out_10(rand_exe_prng_39_io_out_10),
    .io_out_11(rand_exe_prng_39_io_out_11),
    .io_out_12(rand_exe_prng_39_io_out_12),
    .io_out_13(rand_exe_prng_39_io_out_13),
    .io_out_14(rand_exe_prng_39_io_out_14),
    .io_out_15(rand_exe_prng_39_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_40 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_40_clock),
    .reset(rand_exe_prng_40_reset),
    .io_out_0(rand_exe_prng_40_io_out_0),
    .io_out_1(rand_exe_prng_40_io_out_1),
    .io_out_2(rand_exe_prng_40_io_out_2),
    .io_out_3(rand_exe_prng_40_io_out_3),
    .io_out_4(rand_exe_prng_40_io_out_4),
    .io_out_5(rand_exe_prng_40_io_out_5),
    .io_out_6(rand_exe_prng_40_io_out_6),
    .io_out_7(rand_exe_prng_40_io_out_7),
    .io_out_8(rand_exe_prng_40_io_out_8),
    .io_out_9(rand_exe_prng_40_io_out_9),
    .io_out_10(rand_exe_prng_40_io_out_10),
    .io_out_11(rand_exe_prng_40_io_out_11),
    .io_out_12(rand_exe_prng_40_io_out_12),
    .io_out_13(rand_exe_prng_40_io_out_13),
    .io_out_14(rand_exe_prng_40_io_out_14),
    .io_out_15(rand_exe_prng_40_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_41 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_41_clock),
    .reset(rand_exe_prng_41_reset),
    .io_out_0(rand_exe_prng_41_io_out_0),
    .io_out_1(rand_exe_prng_41_io_out_1),
    .io_out_2(rand_exe_prng_41_io_out_2),
    .io_out_3(rand_exe_prng_41_io_out_3),
    .io_out_4(rand_exe_prng_41_io_out_4),
    .io_out_5(rand_exe_prng_41_io_out_5),
    .io_out_6(rand_exe_prng_41_io_out_6),
    .io_out_7(rand_exe_prng_41_io_out_7),
    .io_out_8(rand_exe_prng_41_io_out_8),
    .io_out_9(rand_exe_prng_41_io_out_9),
    .io_out_10(rand_exe_prng_41_io_out_10),
    .io_out_11(rand_exe_prng_41_io_out_11),
    .io_out_12(rand_exe_prng_41_io_out_12),
    .io_out_13(rand_exe_prng_41_io_out_13),
    .io_out_14(rand_exe_prng_41_io_out_14),
    .io_out_15(rand_exe_prng_41_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_42 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_42_clock),
    .reset(rand_exe_prng_42_reset),
    .io_out_0(rand_exe_prng_42_io_out_0),
    .io_out_1(rand_exe_prng_42_io_out_1),
    .io_out_2(rand_exe_prng_42_io_out_2),
    .io_out_3(rand_exe_prng_42_io_out_3),
    .io_out_4(rand_exe_prng_42_io_out_4),
    .io_out_5(rand_exe_prng_42_io_out_5),
    .io_out_6(rand_exe_prng_42_io_out_6),
    .io_out_7(rand_exe_prng_42_io_out_7),
    .io_out_8(rand_exe_prng_42_io_out_8),
    .io_out_9(rand_exe_prng_42_io_out_9),
    .io_out_10(rand_exe_prng_42_io_out_10),
    .io_out_11(rand_exe_prng_42_io_out_11),
    .io_out_12(rand_exe_prng_42_io_out_12),
    .io_out_13(rand_exe_prng_42_io_out_13),
    .io_out_14(rand_exe_prng_42_io_out_14),
    .io_out_15(rand_exe_prng_42_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_43 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_43_clock),
    .reset(rand_exe_prng_43_reset),
    .io_out_0(rand_exe_prng_43_io_out_0),
    .io_out_1(rand_exe_prng_43_io_out_1),
    .io_out_2(rand_exe_prng_43_io_out_2),
    .io_out_3(rand_exe_prng_43_io_out_3),
    .io_out_4(rand_exe_prng_43_io_out_4),
    .io_out_5(rand_exe_prng_43_io_out_5),
    .io_out_6(rand_exe_prng_43_io_out_6),
    .io_out_7(rand_exe_prng_43_io_out_7),
    .io_out_8(rand_exe_prng_43_io_out_8),
    .io_out_9(rand_exe_prng_43_io_out_9),
    .io_out_10(rand_exe_prng_43_io_out_10),
    .io_out_11(rand_exe_prng_43_io_out_11),
    .io_out_12(rand_exe_prng_43_io_out_12),
    .io_out_13(rand_exe_prng_43_io_out_13),
    .io_out_14(rand_exe_prng_43_io_out_14),
    .io_out_15(rand_exe_prng_43_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_44 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_44_clock),
    .reset(rand_exe_prng_44_reset),
    .io_out_0(rand_exe_prng_44_io_out_0),
    .io_out_1(rand_exe_prng_44_io_out_1),
    .io_out_2(rand_exe_prng_44_io_out_2),
    .io_out_3(rand_exe_prng_44_io_out_3),
    .io_out_4(rand_exe_prng_44_io_out_4),
    .io_out_5(rand_exe_prng_44_io_out_5),
    .io_out_6(rand_exe_prng_44_io_out_6),
    .io_out_7(rand_exe_prng_44_io_out_7),
    .io_out_8(rand_exe_prng_44_io_out_8),
    .io_out_9(rand_exe_prng_44_io_out_9),
    .io_out_10(rand_exe_prng_44_io_out_10),
    .io_out_11(rand_exe_prng_44_io_out_11),
    .io_out_12(rand_exe_prng_44_io_out_12),
    .io_out_13(rand_exe_prng_44_io_out_13),
    .io_out_14(rand_exe_prng_44_io_out_14),
    .io_out_15(rand_exe_prng_44_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_45 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_45_clock),
    .reset(rand_exe_prng_45_reset),
    .io_out_0(rand_exe_prng_45_io_out_0),
    .io_out_1(rand_exe_prng_45_io_out_1),
    .io_out_2(rand_exe_prng_45_io_out_2),
    .io_out_3(rand_exe_prng_45_io_out_3),
    .io_out_4(rand_exe_prng_45_io_out_4),
    .io_out_5(rand_exe_prng_45_io_out_5),
    .io_out_6(rand_exe_prng_45_io_out_6),
    .io_out_7(rand_exe_prng_45_io_out_7),
    .io_out_8(rand_exe_prng_45_io_out_8),
    .io_out_9(rand_exe_prng_45_io_out_9),
    .io_out_10(rand_exe_prng_45_io_out_10),
    .io_out_11(rand_exe_prng_45_io_out_11),
    .io_out_12(rand_exe_prng_45_io_out_12),
    .io_out_13(rand_exe_prng_45_io_out_13),
    .io_out_14(rand_exe_prng_45_io_out_14),
    .io_out_15(rand_exe_prng_45_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_46 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_46_clock),
    .reset(rand_exe_prng_46_reset),
    .io_out_0(rand_exe_prng_46_io_out_0),
    .io_out_1(rand_exe_prng_46_io_out_1),
    .io_out_2(rand_exe_prng_46_io_out_2),
    .io_out_3(rand_exe_prng_46_io_out_3),
    .io_out_4(rand_exe_prng_46_io_out_4),
    .io_out_5(rand_exe_prng_46_io_out_5),
    .io_out_6(rand_exe_prng_46_io_out_6),
    .io_out_7(rand_exe_prng_46_io_out_7),
    .io_out_8(rand_exe_prng_46_io_out_8),
    .io_out_9(rand_exe_prng_46_io_out_9),
    .io_out_10(rand_exe_prng_46_io_out_10),
    .io_out_11(rand_exe_prng_46_io_out_11),
    .io_out_12(rand_exe_prng_46_io_out_12),
    .io_out_13(rand_exe_prng_46_io_out_13),
    .io_out_14(rand_exe_prng_46_io_out_14),
    .io_out_15(rand_exe_prng_46_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_47 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_47_clock),
    .reset(rand_exe_prng_47_reset),
    .io_out_0(rand_exe_prng_47_io_out_0),
    .io_out_1(rand_exe_prng_47_io_out_1),
    .io_out_2(rand_exe_prng_47_io_out_2),
    .io_out_3(rand_exe_prng_47_io_out_3),
    .io_out_4(rand_exe_prng_47_io_out_4),
    .io_out_5(rand_exe_prng_47_io_out_5),
    .io_out_6(rand_exe_prng_47_io_out_6),
    .io_out_7(rand_exe_prng_47_io_out_7),
    .io_out_8(rand_exe_prng_47_io_out_8),
    .io_out_9(rand_exe_prng_47_io_out_9),
    .io_out_10(rand_exe_prng_47_io_out_10),
    .io_out_11(rand_exe_prng_47_io_out_11),
    .io_out_12(rand_exe_prng_47_io_out_12),
    .io_out_13(rand_exe_prng_47_io_out_13),
    .io_out_14(rand_exe_prng_47_io_out_14),
    .io_out_15(rand_exe_prng_47_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_48 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_48_clock),
    .reset(rand_exe_prng_48_reset),
    .io_out_0(rand_exe_prng_48_io_out_0),
    .io_out_1(rand_exe_prng_48_io_out_1),
    .io_out_2(rand_exe_prng_48_io_out_2),
    .io_out_3(rand_exe_prng_48_io_out_3),
    .io_out_4(rand_exe_prng_48_io_out_4),
    .io_out_5(rand_exe_prng_48_io_out_5),
    .io_out_6(rand_exe_prng_48_io_out_6),
    .io_out_7(rand_exe_prng_48_io_out_7),
    .io_out_8(rand_exe_prng_48_io_out_8),
    .io_out_9(rand_exe_prng_48_io_out_9),
    .io_out_10(rand_exe_prng_48_io_out_10),
    .io_out_11(rand_exe_prng_48_io_out_11),
    .io_out_12(rand_exe_prng_48_io_out_12),
    .io_out_13(rand_exe_prng_48_io_out_13),
    .io_out_14(rand_exe_prng_48_io_out_14),
    .io_out_15(rand_exe_prng_48_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_49 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_49_clock),
    .reset(rand_exe_prng_49_reset),
    .io_out_0(rand_exe_prng_49_io_out_0),
    .io_out_1(rand_exe_prng_49_io_out_1),
    .io_out_2(rand_exe_prng_49_io_out_2),
    .io_out_3(rand_exe_prng_49_io_out_3),
    .io_out_4(rand_exe_prng_49_io_out_4),
    .io_out_5(rand_exe_prng_49_io_out_5),
    .io_out_6(rand_exe_prng_49_io_out_6),
    .io_out_7(rand_exe_prng_49_io_out_7),
    .io_out_8(rand_exe_prng_49_io_out_8),
    .io_out_9(rand_exe_prng_49_io_out_9),
    .io_out_10(rand_exe_prng_49_io_out_10),
    .io_out_11(rand_exe_prng_49_io_out_11),
    .io_out_12(rand_exe_prng_49_io_out_12),
    .io_out_13(rand_exe_prng_49_io_out_13),
    .io_out_14(rand_exe_prng_49_io_out_14),
    .io_out_15(rand_exe_prng_49_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_50 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_50_clock),
    .reset(rand_exe_prng_50_reset),
    .io_out_0(rand_exe_prng_50_io_out_0),
    .io_out_1(rand_exe_prng_50_io_out_1),
    .io_out_2(rand_exe_prng_50_io_out_2),
    .io_out_3(rand_exe_prng_50_io_out_3),
    .io_out_4(rand_exe_prng_50_io_out_4),
    .io_out_5(rand_exe_prng_50_io_out_5),
    .io_out_6(rand_exe_prng_50_io_out_6),
    .io_out_7(rand_exe_prng_50_io_out_7),
    .io_out_8(rand_exe_prng_50_io_out_8),
    .io_out_9(rand_exe_prng_50_io_out_9),
    .io_out_10(rand_exe_prng_50_io_out_10),
    .io_out_11(rand_exe_prng_50_io_out_11),
    .io_out_12(rand_exe_prng_50_io_out_12),
    .io_out_13(rand_exe_prng_50_io_out_13),
    .io_out_14(rand_exe_prng_50_io_out_14),
    .io_out_15(rand_exe_prng_50_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_51 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_51_clock),
    .reset(rand_exe_prng_51_reset),
    .io_out_0(rand_exe_prng_51_io_out_0),
    .io_out_1(rand_exe_prng_51_io_out_1),
    .io_out_2(rand_exe_prng_51_io_out_2),
    .io_out_3(rand_exe_prng_51_io_out_3),
    .io_out_4(rand_exe_prng_51_io_out_4),
    .io_out_5(rand_exe_prng_51_io_out_5),
    .io_out_6(rand_exe_prng_51_io_out_6),
    .io_out_7(rand_exe_prng_51_io_out_7),
    .io_out_8(rand_exe_prng_51_io_out_8),
    .io_out_9(rand_exe_prng_51_io_out_9),
    .io_out_10(rand_exe_prng_51_io_out_10),
    .io_out_11(rand_exe_prng_51_io_out_11),
    .io_out_12(rand_exe_prng_51_io_out_12),
    .io_out_13(rand_exe_prng_51_io_out_13),
    .io_out_14(rand_exe_prng_51_io_out_14),
    .io_out_15(rand_exe_prng_51_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_52 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_52_clock),
    .reset(rand_exe_prng_52_reset),
    .io_out_0(rand_exe_prng_52_io_out_0),
    .io_out_1(rand_exe_prng_52_io_out_1),
    .io_out_2(rand_exe_prng_52_io_out_2),
    .io_out_3(rand_exe_prng_52_io_out_3),
    .io_out_4(rand_exe_prng_52_io_out_4),
    .io_out_5(rand_exe_prng_52_io_out_5),
    .io_out_6(rand_exe_prng_52_io_out_6),
    .io_out_7(rand_exe_prng_52_io_out_7),
    .io_out_8(rand_exe_prng_52_io_out_8),
    .io_out_9(rand_exe_prng_52_io_out_9),
    .io_out_10(rand_exe_prng_52_io_out_10),
    .io_out_11(rand_exe_prng_52_io_out_11),
    .io_out_12(rand_exe_prng_52_io_out_12),
    .io_out_13(rand_exe_prng_52_io_out_13),
    .io_out_14(rand_exe_prng_52_io_out_14),
    .io_out_15(rand_exe_prng_52_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_53 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_53_clock),
    .reset(rand_exe_prng_53_reset),
    .io_out_0(rand_exe_prng_53_io_out_0),
    .io_out_1(rand_exe_prng_53_io_out_1),
    .io_out_2(rand_exe_prng_53_io_out_2),
    .io_out_3(rand_exe_prng_53_io_out_3),
    .io_out_4(rand_exe_prng_53_io_out_4),
    .io_out_5(rand_exe_prng_53_io_out_5),
    .io_out_6(rand_exe_prng_53_io_out_6),
    .io_out_7(rand_exe_prng_53_io_out_7),
    .io_out_8(rand_exe_prng_53_io_out_8),
    .io_out_9(rand_exe_prng_53_io_out_9),
    .io_out_10(rand_exe_prng_53_io_out_10),
    .io_out_11(rand_exe_prng_53_io_out_11),
    .io_out_12(rand_exe_prng_53_io_out_12),
    .io_out_13(rand_exe_prng_53_io_out_13),
    .io_out_14(rand_exe_prng_53_io_out_14),
    .io_out_15(rand_exe_prng_53_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_54 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_54_clock),
    .reset(rand_exe_prng_54_reset),
    .io_out_0(rand_exe_prng_54_io_out_0),
    .io_out_1(rand_exe_prng_54_io_out_1),
    .io_out_2(rand_exe_prng_54_io_out_2),
    .io_out_3(rand_exe_prng_54_io_out_3),
    .io_out_4(rand_exe_prng_54_io_out_4),
    .io_out_5(rand_exe_prng_54_io_out_5),
    .io_out_6(rand_exe_prng_54_io_out_6),
    .io_out_7(rand_exe_prng_54_io_out_7),
    .io_out_8(rand_exe_prng_54_io_out_8),
    .io_out_9(rand_exe_prng_54_io_out_9),
    .io_out_10(rand_exe_prng_54_io_out_10),
    .io_out_11(rand_exe_prng_54_io_out_11),
    .io_out_12(rand_exe_prng_54_io_out_12),
    .io_out_13(rand_exe_prng_54_io_out_13),
    .io_out_14(rand_exe_prng_54_io_out_14),
    .io_out_15(rand_exe_prng_54_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_55 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_55_clock),
    .reset(rand_exe_prng_55_reset),
    .io_out_0(rand_exe_prng_55_io_out_0),
    .io_out_1(rand_exe_prng_55_io_out_1),
    .io_out_2(rand_exe_prng_55_io_out_2),
    .io_out_3(rand_exe_prng_55_io_out_3),
    .io_out_4(rand_exe_prng_55_io_out_4),
    .io_out_5(rand_exe_prng_55_io_out_5),
    .io_out_6(rand_exe_prng_55_io_out_6),
    .io_out_7(rand_exe_prng_55_io_out_7),
    .io_out_8(rand_exe_prng_55_io_out_8),
    .io_out_9(rand_exe_prng_55_io_out_9),
    .io_out_10(rand_exe_prng_55_io_out_10),
    .io_out_11(rand_exe_prng_55_io_out_11),
    .io_out_12(rand_exe_prng_55_io_out_12),
    .io_out_13(rand_exe_prng_55_io_out_13),
    .io_out_14(rand_exe_prng_55_io_out_14),
    .io_out_15(rand_exe_prng_55_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_56 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_56_clock),
    .reset(rand_exe_prng_56_reset),
    .io_out_0(rand_exe_prng_56_io_out_0),
    .io_out_1(rand_exe_prng_56_io_out_1),
    .io_out_2(rand_exe_prng_56_io_out_2),
    .io_out_3(rand_exe_prng_56_io_out_3),
    .io_out_4(rand_exe_prng_56_io_out_4),
    .io_out_5(rand_exe_prng_56_io_out_5),
    .io_out_6(rand_exe_prng_56_io_out_6),
    .io_out_7(rand_exe_prng_56_io_out_7),
    .io_out_8(rand_exe_prng_56_io_out_8),
    .io_out_9(rand_exe_prng_56_io_out_9),
    .io_out_10(rand_exe_prng_56_io_out_10),
    .io_out_11(rand_exe_prng_56_io_out_11),
    .io_out_12(rand_exe_prng_56_io_out_12),
    .io_out_13(rand_exe_prng_56_io_out_13),
    .io_out_14(rand_exe_prng_56_io_out_14),
    .io_out_15(rand_exe_prng_56_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_57 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_57_clock),
    .reset(rand_exe_prng_57_reset),
    .io_out_0(rand_exe_prng_57_io_out_0),
    .io_out_1(rand_exe_prng_57_io_out_1),
    .io_out_2(rand_exe_prng_57_io_out_2),
    .io_out_3(rand_exe_prng_57_io_out_3),
    .io_out_4(rand_exe_prng_57_io_out_4),
    .io_out_5(rand_exe_prng_57_io_out_5),
    .io_out_6(rand_exe_prng_57_io_out_6),
    .io_out_7(rand_exe_prng_57_io_out_7),
    .io_out_8(rand_exe_prng_57_io_out_8),
    .io_out_9(rand_exe_prng_57_io_out_9),
    .io_out_10(rand_exe_prng_57_io_out_10),
    .io_out_11(rand_exe_prng_57_io_out_11),
    .io_out_12(rand_exe_prng_57_io_out_12),
    .io_out_13(rand_exe_prng_57_io_out_13),
    .io_out_14(rand_exe_prng_57_io_out_14),
    .io_out_15(rand_exe_prng_57_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_58 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_58_clock),
    .reset(rand_exe_prng_58_reset),
    .io_out_0(rand_exe_prng_58_io_out_0),
    .io_out_1(rand_exe_prng_58_io_out_1),
    .io_out_2(rand_exe_prng_58_io_out_2),
    .io_out_3(rand_exe_prng_58_io_out_3),
    .io_out_4(rand_exe_prng_58_io_out_4),
    .io_out_5(rand_exe_prng_58_io_out_5),
    .io_out_6(rand_exe_prng_58_io_out_6),
    .io_out_7(rand_exe_prng_58_io_out_7),
    .io_out_8(rand_exe_prng_58_io_out_8),
    .io_out_9(rand_exe_prng_58_io_out_9),
    .io_out_10(rand_exe_prng_58_io_out_10),
    .io_out_11(rand_exe_prng_58_io_out_11),
    .io_out_12(rand_exe_prng_58_io_out_12),
    .io_out_13(rand_exe_prng_58_io_out_13),
    .io_out_14(rand_exe_prng_58_io_out_14),
    .io_out_15(rand_exe_prng_58_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_59 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_59_clock),
    .reset(rand_exe_prng_59_reset),
    .io_out_0(rand_exe_prng_59_io_out_0),
    .io_out_1(rand_exe_prng_59_io_out_1),
    .io_out_2(rand_exe_prng_59_io_out_2),
    .io_out_3(rand_exe_prng_59_io_out_3),
    .io_out_4(rand_exe_prng_59_io_out_4),
    .io_out_5(rand_exe_prng_59_io_out_5),
    .io_out_6(rand_exe_prng_59_io_out_6),
    .io_out_7(rand_exe_prng_59_io_out_7),
    .io_out_8(rand_exe_prng_59_io_out_8),
    .io_out_9(rand_exe_prng_59_io_out_9),
    .io_out_10(rand_exe_prng_59_io_out_10),
    .io_out_11(rand_exe_prng_59_io_out_11),
    .io_out_12(rand_exe_prng_59_io_out_12),
    .io_out_13(rand_exe_prng_59_io_out_13),
    .io_out_14(rand_exe_prng_59_io_out_14),
    .io_out_15(rand_exe_prng_59_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_60 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_60_clock),
    .reset(rand_exe_prng_60_reset),
    .io_out_0(rand_exe_prng_60_io_out_0),
    .io_out_1(rand_exe_prng_60_io_out_1),
    .io_out_2(rand_exe_prng_60_io_out_2),
    .io_out_3(rand_exe_prng_60_io_out_3),
    .io_out_4(rand_exe_prng_60_io_out_4),
    .io_out_5(rand_exe_prng_60_io_out_5),
    .io_out_6(rand_exe_prng_60_io_out_6),
    .io_out_7(rand_exe_prng_60_io_out_7),
    .io_out_8(rand_exe_prng_60_io_out_8),
    .io_out_9(rand_exe_prng_60_io_out_9),
    .io_out_10(rand_exe_prng_60_io_out_10),
    .io_out_11(rand_exe_prng_60_io_out_11),
    .io_out_12(rand_exe_prng_60_io_out_12),
    .io_out_13(rand_exe_prng_60_io_out_13),
    .io_out_14(rand_exe_prng_60_io_out_14),
    .io_out_15(rand_exe_prng_60_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_61 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_61_clock),
    .reset(rand_exe_prng_61_reset),
    .io_out_0(rand_exe_prng_61_io_out_0),
    .io_out_1(rand_exe_prng_61_io_out_1),
    .io_out_2(rand_exe_prng_61_io_out_2),
    .io_out_3(rand_exe_prng_61_io_out_3),
    .io_out_4(rand_exe_prng_61_io_out_4),
    .io_out_5(rand_exe_prng_61_io_out_5),
    .io_out_6(rand_exe_prng_61_io_out_6),
    .io_out_7(rand_exe_prng_61_io_out_7),
    .io_out_8(rand_exe_prng_61_io_out_8),
    .io_out_9(rand_exe_prng_61_io_out_9),
    .io_out_10(rand_exe_prng_61_io_out_10),
    .io_out_11(rand_exe_prng_61_io_out_11),
    .io_out_12(rand_exe_prng_61_io_out_12),
    .io_out_13(rand_exe_prng_61_io_out_13),
    .io_out_14(rand_exe_prng_61_io_out_14),
    .io_out_15(rand_exe_prng_61_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_62 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_62_clock),
    .reset(rand_exe_prng_62_reset),
    .io_out_0(rand_exe_prng_62_io_out_0),
    .io_out_1(rand_exe_prng_62_io_out_1),
    .io_out_2(rand_exe_prng_62_io_out_2),
    .io_out_3(rand_exe_prng_62_io_out_3),
    .io_out_4(rand_exe_prng_62_io_out_4),
    .io_out_5(rand_exe_prng_62_io_out_5),
    .io_out_6(rand_exe_prng_62_io_out_6),
    .io_out_7(rand_exe_prng_62_io_out_7),
    .io_out_8(rand_exe_prng_62_io_out_8),
    .io_out_9(rand_exe_prng_62_io_out_9),
    .io_out_10(rand_exe_prng_62_io_out_10),
    .io_out_11(rand_exe_prng_62_io_out_11),
    .io_out_12(rand_exe_prng_62_io_out_12),
    .io_out_13(rand_exe_prng_62_io_out_13),
    .io_out_14(rand_exe_prng_62_io_out_14),
    .io_out_15(rand_exe_prng_62_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_63 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_63_clock),
    .reset(rand_exe_prng_63_reset),
    .io_out_0(rand_exe_prng_63_io_out_0),
    .io_out_1(rand_exe_prng_63_io_out_1),
    .io_out_2(rand_exe_prng_63_io_out_2),
    .io_out_3(rand_exe_prng_63_io_out_3),
    .io_out_4(rand_exe_prng_63_io_out_4),
    .io_out_5(rand_exe_prng_63_io_out_5),
    .io_out_6(rand_exe_prng_63_io_out_6),
    .io_out_7(rand_exe_prng_63_io_out_7),
    .io_out_8(rand_exe_prng_63_io_out_8),
    .io_out_9(rand_exe_prng_63_io_out_9),
    .io_out_10(rand_exe_prng_63_io_out_10),
    .io_out_11(rand_exe_prng_63_io_out_11),
    .io_out_12(rand_exe_prng_63_io_out_12),
    .io_out_13(rand_exe_prng_63_io_out_13),
    .io_out_14(rand_exe_prng_63_io_out_14),
    .io_out_15(rand_exe_prng_63_io_out_15)
  );
  assign io_phv_out_data_0 = rand_0[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_1 = rand_0[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_2 = rand_1[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_3 = rand_1[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_4 = rand_2[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_5 = rand_2[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_6 = rand_3[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_7 = rand_3[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_8 = rand_4[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_9 = rand_4[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_10 = rand_5[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_11 = rand_5[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_12 = rand_6[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_13 = rand_6[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_14 = rand_7[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_15 = rand_7[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_16 = rand_8[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_17 = rand_8[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_18 = rand_9[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_19 = rand_9[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_20 = rand_10[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_21 = rand_10[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_22 = rand_11[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_23 = rand_11[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_24 = rand_12[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_25 = rand_12[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_26 = rand_13[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_27 = rand_13[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_28 = rand_14[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_29 = rand_14[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_30 = rand_15[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_31 = rand_15[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_32 = rand_16[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_33 = rand_16[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_34 = rand_17[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_35 = rand_17[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_36 = rand_18[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_37 = rand_18[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_38 = rand_19[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_39 = rand_19[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_40 = rand_20[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_41 = rand_20[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_42 = rand_21[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_43 = rand_21[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_44 = rand_22[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_45 = rand_22[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_46 = rand_23[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_47 = rand_23[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_48 = rand_24[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_49 = rand_24[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_50 = rand_25[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_51 = rand_25[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_52 = rand_26[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_53 = rand_26[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_54 = rand_27[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_55 = rand_27[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_56 = rand_28[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_57 = rand_28[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_58 = rand_29[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_59 = rand_29[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_60 = rand_30[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_61 = rand_30[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_62 = rand_31[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_63 = rand_31[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_64 = rand_32[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_65 = rand_32[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_66 = rand_33[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_67 = rand_33[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_68 = rand_34[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_69 = rand_34[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_70 = rand_35[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_71 = rand_35[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_72 = rand_36[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_73 = rand_36[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_74 = rand_37[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_75 = rand_37[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_76 = rand_38[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_77 = rand_38[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_78 = rand_39[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_79 = rand_39[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_80 = rand_40[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_81 = rand_40[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_82 = rand_41[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_83 = rand_41[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_84 = rand_42[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_85 = rand_42[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_86 = rand_43[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_87 = rand_43[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_88 = rand_44[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_89 = rand_44[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_90 = rand_45[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_91 = rand_45[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_92 = rand_46[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_93 = rand_46[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_94 = rand_47[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_95 = rand_47[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_96 = rand_48[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_97 = rand_48[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_98 = rand_49[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_99 = rand_49[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_100 = rand_50[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_101 = rand_50[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_102 = rand_51[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_103 = rand_51[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_104 = rand_52[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_105 = rand_52[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_106 = rand_53[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_107 = rand_53[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_108 = rand_54[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_109 = rand_54[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_110 = rand_55[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_111 = rand_55[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_112 = rand_56[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_113 = rand_56[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_114 = rand_57[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_115 = rand_57[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_116 = rand_58[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_117 = rand_58[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_118 = rand_59[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_119 = rand_59[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_120 = rand_60[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_121 = rand_60[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_122 = rand_61[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_123 = rand_61[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_124 = rand_62[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_125 = rand_62[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_126 = rand_63[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_127 = rand_63[7:0]; // @[inport.scala 19:42]
  assign rand_exe_prng_clock = clock;
  assign rand_exe_prng_reset = reset;
  assign rand_exe_prng_1_clock = clock;
  assign rand_exe_prng_1_reset = reset;
  assign rand_exe_prng_2_clock = clock;
  assign rand_exe_prng_2_reset = reset;
  assign rand_exe_prng_3_clock = clock;
  assign rand_exe_prng_3_reset = reset;
  assign rand_exe_prng_4_clock = clock;
  assign rand_exe_prng_4_reset = reset;
  assign rand_exe_prng_5_clock = clock;
  assign rand_exe_prng_5_reset = reset;
  assign rand_exe_prng_6_clock = clock;
  assign rand_exe_prng_6_reset = reset;
  assign rand_exe_prng_7_clock = clock;
  assign rand_exe_prng_7_reset = reset;
  assign rand_exe_prng_8_clock = clock;
  assign rand_exe_prng_8_reset = reset;
  assign rand_exe_prng_9_clock = clock;
  assign rand_exe_prng_9_reset = reset;
  assign rand_exe_prng_10_clock = clock;
  assign rand_exe_prng_10_reset = reset;
  assign rand_exe_prng_11_clock = clock;
  assign rand_exe_prng_11_reset = reset;
  assign rand_exe_prng_12_clock = clock;
  assign rand_exe_prng_12_reset = reset;
  assign rand_exe_prng_13_clock = clock;
  assign rand_exe_prng_13_reset = reset;
  assign rand_exe_prng_14_clock = clock;
  assign rand_exe_prng_14_reset = reset;
  assign rand_exe_prng_15_clock = clock;
  assign rand_exe_prng_15_reset = reset;
  assign rand_exe_prng_16_clock = clock;
  assign rand_exe_prng_16_reset = reset;
  assign rand_exe_prng_17_clock = clock;
  assign rand_exe_prng_17_reset = reset;
  assign rand_exe_prng_18_clock = clock;
  assign rand_exe_prng_18_reset = reset;
  assign rand_exe_prng_19_clock = clock;
  assign rand_exe_prng_19_reset = reset;
  assign rand_exe_prng_20_clock = clock;
  assign rand_exe_prng_20_reset = reset;
  assign rand_exe_prng_21_clock = clock;
  assign rand_exe_prng_21_reset = reset;
  assign rand_exe_prng_22_clock = clock;
  assign rand_exe_prng_22_reset = reset;
  assign rand_exe_prng_23_clock = clock;
  assign rand_exe_prng_23_reset = reset;
  assign rand_exe_prng_24_clock = clock;
  assign rand_exe_prng_24_reset = reset;
  assign rand_exe_prng_25_clock = clock;
  assign rand_exe_prng_25_reset = reset;
  assign rand_exe_prng_26_clock = clock;
  assign rand_exe_prng_26_reset = reset;
  assign rand_exe_prng_27_clock = clock;
  assign rand_exe_prng_27_reset = reset;
  assign rand_exe_prng_28_clock = clock;
  assign rand_exe_prng_28_reset = reset;
  assign rand_exe_prng_29_clock = clock;
  assign rand_exe_prng_29_reset = reset;
  assign rand_exe_prng_30_clock = clock;
  assign rand_exe_prng_30_reset = reset;
  assign rand_exe_prng_31_clock = clock;
  assign rand_exe_prng_31_reset = reset;
  assign rand_exe_prng_32_clock = clock;
  assign rand_exe_prng_32_reset = reset;
  assign rand_exe_prng_33_clock = clock;
  assign rand_exe_prng_33_reset = reset;
  assign rand_exe_prng_34_clock = clock;
  assign rand_exe_prng_34_reset = reset;
  assign rand_exe_prng_35_clock = clock;
  assign rand_exe_prng_35_reset = reset;
  assign rand_exe_prng_36_clock = clock;
  assign rand_exe_prng_36_reset = reset;
  assign rand_exe_prng_37_clock = clock;
  assign rand_exe_prng_37_reset = reset;
  assign rand_exe_prng_38_clock = clock;
  assign rand_exe_prng_38_reset = reset;
  assign rand_exe_prng_39_clock = clock;
  assign rand_exe_prng_39_reset = reset;
  assign rand_exe_prng_40_clock = clock;
  assign rand_exe_prng_40_reset = reset;
  assign rand_exe_prng_41_clock = clock;
  assign rand_exe_prng_41_reset = reset;
  assign rand_exe_prng_42_clock = clock;
  assign rand_exe_prng_42_reset = reset;
  assign rand_exe_prng_43_clock = clock;
  assign rand_exe_prng_43_reset = reset;
  assign rand_exe_prng_44_clock = clock;
  assign rand_exe_prng_44_reset = reset;
  assign rand_exe_prng_45_clock = clock;
  assign rand_exe_prng_45_reset = reset;
  assign rand_exe_prng_46_clock = clock;
  assign rand_exe_prng_46_reset = reset;
  assign rand_exe_prng_47_clock = clock;
  assign rand_exe_prng_47_reset = reset;
  assign rand_exe_prng_48_clock = clock;
  assign rand_exe_prng_48_reset = reset;
  assign rand_exe_prng_49_clock = clock;
  assign rand_exe_prng_49_reset = reset;
  assign rand_exe_prng_50_clock = clock;
  assign rand_exe_prng_50_reset = reset;
  assign rand_exe_prng_51_clock = clock;
  assign rand_exe_prng_51_reset = reset;
  assign rand_exe_prng_52_clock = clock;
  assign rand_exe_prng_52_reset = reset;
  assign rand_exe_prng_53_clock = clock;
  assign rand_exe_prng_53_reset = reset;
  assign rand_exe_prng_54_clock = clock;
  assign rand_exe_prng_54_reset = reset;
  assign rand_exe_prng_55_clock = clock;
  assign rand_exe_prng_55_reset = reset;
  assign rand_exe_prng_56_clock = clock;
  assign rand_exe_prng_56_reset = reset;
  assign rand_exe_prng_57_clock = clock;
  assign rand_exe_prng_57_reset = reset;
  assign rand_exe_prng_58_clock = clock;
  assign rand_exe_prng_58_reset = reset;
  assign rand_exe_prng_59_clock = clock;
  assign rand_exe_prng_59_reset = reset;
  assign rand_exe_prng_60_clock = clock;
  assign rand_exe_prng_60_reset = reset;
  assign rand_exe_prng_61_clock = clock;
  assign rand_exe_prng_61_reset = reset;
  assign rand_exe_prng_62_clock = clock;
  assign rand_exe_prng_62_reset = reset;
  assign rand_exe_prng_63_clock = clock;
  assign rand_exe_prng_63_reset = reset;
endmodule
