module OutPort(
  input  [7:0]    io_phv_in_data_0,
  input  [7:0]    io_phv_in_data_1,
  input  [7:0]    io_phv_in_data_2,
  input  [7:0]    io_phv_in_data_3,
  input  [7:0]    io_phv_in_data_4,
  input  [7:0]    io_phv_in_data_5,
  input  [7:0]    io_phv_in_data_6,
  input  [7:0]    io_phv_in_data_7,
  input  [7:0]    io_phv_in_data_8,
  input  [7:0]    io_phv_in_data_9,
  input  [7:0]    io_phv_in_data_10,
  input  [7:0]    io_phv_in_data_11,
  input  [7:0]    io_phv_in_data_12,
  input  [7:0]    io_phv_in_data_13,
  input  [7:0]    io_phv_in_data_14,
  input  [7:0]    io_phv_in_data_15,
  input  [7:0]    io_phv_in_data_16,
  input  [7:0]    io_phv_in_data_17,
  input  [7:0]    io_phv_in_data_18,
  input  [7:0]    io_phv_in_data_19,
  input  [7:0]    io_phv_in_data_20,
  input  [7:0]    io_phv_in_data_21,
  input  [7:0]    io_phv_in_data_22,
  input  [7:0]    io_phv_in_data_23,
  input  [7:0]    io_phv_in_data_24,
  input  [7:0]    io_phv_in_data_25,
  input  [7:0]    io_phv_in_data_26,
  input  [7:0]    io_phv_in_data_27,
  input  [7:0]    io_phv_in_data_28,
  input  [7:0]    io_phv_in_data_29,
  input  [7:0]    io_phv_in_data_30,
  input  [7:0]    io_phv_in_data_31,
  input  [7:0]    io_phv_in_data_32,
  input  [7:0]    io_phv_in_data_33,
  input  [7:0]    io_phv_in_data_34,
  input  [7:0]    io_phv_in_data_35,
  input  [7:0]    io_phv_in_data_36,
  input  [7:0]    io_phv_in_data_37,
  input  [7:0]    io_phv_in_data_38,
  input  [7:0]    io_phv_in_data_39,
  input  [7:0]    io_phv_in_data_40,
  input  [7:0]    io_phv_in_data_41,
  input  [7:0]    io_phv_in_data_42,
  input  [7:0]    io_phv_in_data_43,
  input  [7:0]    io_phv_in_data_44,
  input  [7:0]    io_phv_in_data_45,
  input  [7:0]    io_phv_in_data_46,
  input  [7:0]    io_phv_in_data_47,
  input  [7:0]    io_phv_in_data_48,
  input  [7:0]    io_phv_in_data_49,
  input  [7:0]    io_phv_in_data_50,
  input  [7:0]    io_phv_in_data_51,
  input  [7:0]    io_phv_in_data_52,
  input  [7:0]    io_phv_in_data_53,
  input  [7:0]    io_phv_in_data_54,
  input  [7:0]    io_phv_in_data_55,
  input  [7:0]    io_phv_in_data_56,
  input  [7:0]    io_phv_in_data_57,
  input  [7:0]    io_phv_in_data_58,
  input  [7:0]    io_phv_in_data_59,
  input  [7:0]    io_phv_in_data_60,
  input  [7:0]    io_phv_in_data_61,
  input  [7:0]    io_phv_in_data_62,
  input  [7:0]    io_phv_in_data_63,
  input  [7:0]    io_phv_in_data_64,
  input  [7:0]    io_phv_in_data_65,
  input  [7:0]    io_phv_in_data_66,
  input  [7:0]    io_phv_in_data_67,
  input  [7:0]    io_phv_in_data_68,
  input  [7:0]    io_phv_in_data_69,
  input  [7:0]    io_phv_in_data_70,
  input  [7:0]    io_phv_in_data_71,
  input  [7:0]    io_phv_in_data_72,
  input  [7:0]    io_phv_in_data_73,
  input  [7:0]    io_phv_in_data_74,
  input  [7:0]    io_phv_in_data_75,
  input  [7:0]    io_phv_in_data_76,
  input  [7:0]    io_phv_in_data_77,
  input  [7:0]    io_phv_in_data_78,
  input  [7:0]    io_phv_in_data_79,
  input  [7:0]    io_phv_in_data_80,
  input  [7:0]    io_phv_in_data_81,
  input  [7:0]    io_phv_in_data_82,
  input  [7:0]    io_phv_in_data_83,
  input  [7:0]    io_phv_in_data_84,
  input  [7:0]    io_phv_in_data_85,
  input  [7:0]    io_phv_in_data_86,
  input  [7:0]    io_phv_in_data_87,
  input  [7:0]    io_phv_in_data_88,
  input  [7:0]    io_phv_in_data_89,
  input  [7:0]    io_phv_in_data_90,
  input  [7:0]    io_phv_in_data_91,
  input  [7:0]    io_phv_in_data_92,
  input  [7:0]    io_phv_in_data_93,
  input  [7:0]    io_phv_in_data_94,
  input  [7:0]    io_phv_in_data_95,
  input  [7:0]    io_phv_in_data_96,
  input  [7:0]    io_phv_in_data_97,
  input  [7:0]    io_phv_in_data_98,
  input  [7:0]    io_phv_in_data_99,
  input  [7:0]    io_phv_in_data_100,
  input  [7:0]    io_phv_in_data_101,
  input  [7:0]    io_phv_in_data_102,
  input  [7:0]    io_phv_in_data_103,
  input  [7:0]    io_phv_in_data_104,
  input  [7:0]    io_phv_in_data_105,
  input  [7:0]    io_phv_in_data_106,
  input  [7:0]    io_phv_in_data_107,
  input  [7:0]    io_phv_in_data_108,
  input  [7:0]    io_phv_in_data_109,
  input  [7:0]    io_phv_in_data_110,
  input  [7:0]    io_phv_in_data_111,
  input  [7:0]    io_phv_in_data_112,
  input  [7:0]    io_phv_in_data_113,
  input  [7:0]    io_phv_in_data_114,
  input  [7:0]    io_phv_in_data_115,
  input  [7:0]    io_phv_in_data_116,
  input  [7:0]    io_phv_in_data_117,
  input  [7:0]    io_phv_in_data_118,
  input  [7:0]    io_phv_in_data_119,
  input  [7:0]    io_phv_in_data_120,
  input  [7:0]    io_phv_in_data_121,
  input  [7:0]    io_phv_in_data_122,
  input  [7:0]    io_phv_in_data_123,
  input  [7:0]    io_phv_in_data_124,
  input  [7:0]    io_phv_in_data_125,
  input  [7:0]    io_phv_in_data_126,
  input  [7:0]    io_phv_in_data_127,
  input           io_phv_in_valid,
  input           io_phv_in_last,
  output [1023:0] io_data,
  output          io_last,
  output          io_en
);
  wire [79:0] io_data_hi_8 = {io_phv_in_data_127,io_phv_in_data_126,io_phv_in_data_125,io_phv_in_data_124,
    io_phv_in_data_123,io_phv_in_data_122,io_phv_in_data_121,io_phv_in_data_120,io_phv_in_data_119,io_phv_in_data_118}; // @[Cat.scala 30:58]
  wire [151:0] io_data_hi_17 = {io_data_hi_8,io_phv_in_data_117,io_phv_in_data_116,io_phv_in_data_115,io_phv_in_data_114
    ,io_phv_in_data_113,io_phv_in_data_112,io_phv_in_data_111,io_phv_in_data_110,io_phv_in_data_109}; // @[Cat.scala 30:58]
  wire [223:0] io_data_hi_26 = {io_data_hi_17,io_phv_in_data_108,io_phv_in_data_107,io_phv_in_data_106,
    io_phv_in_data_105,io_phv_in_data_104,io_phv_in_data_103,io_phv_in_data_102,io_phv_in_data_101,io_phv_in_data_100}; // @[Cat.scala 30:58]
  wire [295:0] io_data_hi_35 = {io_data_hi_26,io_phv_in_data_99,io_phv_in_data_98,io_phv_in_data_97,io_phv_in_data_96,
    io_phv_in_data_95,io_phv_in_data_94,io_phv_in_data_93,io_phv_in_data_92,io_phv_in_data_91}; // @[Cat.scala 30:58]
  wire [367:0] io_data_hi_44 = {io_data_hi_35,io_phv_in_data_90,io_phv_in_data_89,io_phv_in_data_88,io_phv_in_data_87,
    io_phv_in_data_86,io_phv_in_data_85,io_phv_in_data_84,io_phv_in_data_83,io_phv_in_data_82}; // @[Cat.scala 30:58]
  wire [439:0] io_data_hi_53 = {io_data_hi_44,io_phv_in_data_81,io_phv_in_data_80,io_phv_in_data_79,io_phv_in_data_78,
    io_phv_in_data_77,io_phv_in_data_76,io_phv_in_data_75,io_phv_in_data_74,io_phv_in_data_73}; // @[Cat.scala 30:58]
  wire [511:0] io_data_hi_62 = {io_data_hi_53,io_phv_in_data_72,io_phv_in_data_71,io_phv_in_data_70,io_phv_in_data_69,
    io_phv_in_data_68,io_phv_in_data_67,io_phv_in_data_66,io_phv_in_data_65,io_phv_in_data_64}; // @[Cat.scala 30:58]
  wire [583:0] io_data_hi_71 = {io_data_hi_62,io_phv_in_data_63,io_phv_in_data_62,io_phv_in_data_61,io_phv_in_data_60,
    io_phv_in_data_59,io_phv_in_data_58,io_phv_in_data_57,io_phv_in_data_56,io_phv_in_data_55}; // @[Cat.scala 30:58]
  wire [655:0] io_data_hi_80 = {io_data_hi_71,io_phv_in_data_54,io_phv_in_data_53,io_phv_in_data_52,io_phv_in_data_51,
    io_phv_in_data_50,io_phv_in_data_49,io_phv_in_data_48,io_phv_in_data_47,io_phv_in_data_46}; // @[Cat.scala 30:58]
  wire [727:0] io_data_hi_89 = {io_data_hi_80,io_phv_in_data_45,io_phv_in_data_44,io_phv_in_data_43,io_phv_in_data_42,
    io_phv_in_data_41,io_phv_in_data_40,io_phv_in_data_39,io_phv_in_data_38,io_phv_in_data_37}; // @[Cat.scala 30:58]
  wire [799:0] io_data_hi_98 = {io_data_hi_89,io_phv_in_data_36,io_phv_in_data_35,io_phv_in_data_34,io_phv_in_data_33,
    io_phv_in_data_32,io_phv_in_data_31,io_phv_in_data_30,io_phv_in_data_29,io_phv_in_data_28}; // @[Cat.scala 30:58]
  wire [871:0] io_data_hi_107 = {io_data_hi_98,io_phv_in_data_27,io_phv_in_data_26,io_phv_in_data_25,io_phv_in_data_24,
    io_phv_in_data_23,io_phv_in_data_22,io_phv_in_data_21,io_phv_in_data_20,io_phv_in_data_19}; // @[Cat.scala 30:58]
  wire [943:0] io_data_hi_116 = {io_data_hi_107,io_phv_in_data_18,io_phv_in_data_17,io_phv_in_data_16,io_phv_in_data_15,
    io_phv_in_data_14,io_phv_in_data_13,io_phv_in_data_12,io_phv_in_data_11,io_phv_in_data_10}; // @[Cat.scala 30:58]
  wire [1015:0] io_data_hi_125 = {io_data_hi_116,io_phv_in_data_9,io_phv_in_data_8,io_phv_in_data_7,io_phv_in_data_6,
    io_phv_in_data_5,io_phv_in_data_4,io_phv_in_data_3,io_phv_in_data_2,io_phv_in_data_1}; // @[Cat.scala 30:58]
  assign io_data = {io_data_hi_125,io_phv_in_data_0}; // @[Cat.scala 30:58]
  assign io_last = io_phv_in_last; // @[outport.scala 21:13]
  assign io_en = io_phv_in_valid; // @[outport.scala 20:13]
endmodule
