module MatcherPISA(
  input         clock,
  input  [7:0]  io_pipe_phv_in_data_0,
  input  [7:0]  io_pipe_phv_in_data_1,
  input  [7:0]  io_pipe_phv_in_data_2,
  input  [7:0]  io_pipe_phv_in_data_3,
  input  [7:0]  io_pipe_phv_in_data_4,
  input  [7:0]  io_pipe_phv_in_data_5,
  input  [7:0]  io_pipe_phv_in_data_6,
  input  [7:0]  io_pipe_phv_in_data_7,
  input  [7:0]  io_pipe_phv_in_data_8,
  input  [7:0]  io_pipe_phv_in_data_9,
  input  [7:0]  io_pipe_phv_in_data_10,
  input  [7:0]  io_pipe_phv_in_data_11,
  input  [7:0]  io_pipe_phv_in_data_12,
  input  [7:0]  io_pipe_phv_in_data_13,
  input  [7:0]  io_pipe_phv_in_data_14,
  input  [7:0]  io_pipe_phv_in_data_15,
  input  [7:0]  io_pipe_phv_in_data_16,
  input  [7:0]  io_pipe_phv_in_data_17,
  input  [7:0]  io_pipe_phv_in_data_18,
  input  [7:0]  io_pipe_phv_in_data_19,
  input  [7:0]  io_pipe_phv_in_data_20,
  input  [7:0]  io_pipe_phv_in_data_21,
  input  [7:0]  io_pipe_phv_in_data_22,
  input  [7:0]  io_pipe_phv_in_data_23,
  input  [7:0]  io_pipe_phv_in_data_24,
  input  [7:0]  io_pipe_phv_in_data_25,
  input  [7:0]  io_pipe_phv_in_data_26,
  input  [7:0]  io_pipe_phv_in_data_27,
  input  [7:0]  io_pipe_phv_in_data_28,
  input  [7:0]  io_pipe_phv_in_data_29,
  input  [7:0]  io_pipe_phv_in_data_30,
  input  [7:0]  io_pipe_phv_in_data_31,
  input  [7:0]  io_pipe_phv_in_data_32,
  input  [7:0]  io_pipe_phv_in_data_33,
  input  [7:0]  io_pipe_phv_in_data_34,
  input  [7:0]  io_pipe_phv_in_data_35,
  input  [7:0]  io_pipe_phv_in_data_36,
  input  [7:0]  io_pipe_phv_in_data_37,
  input  [7:0]  io_pipe_phv_in_data_38,
  input  [7:0]  io_pipe_phv_in_data_39,
  input  [7:0]  io_pipe_phv_in_data_40,
  input  [7:0]  io_pipe_phv_in_data_41,
  input  [7:0]  io_pipe_phv_in_data_42,
  input  [7:0]  io_pipe_phv_in_data_43,
  input  [7:0]  io_pipe_phv_in_data_44,
  input  [7:0]  io_pipe_phv_in_data_45,
  input  [7:0]  io_pipe_phv_in_data_46,
  input  [7:0]  io_pipe_phv_in_data_47,
  input  [7:0]  io_pipe_phv_in_data_48,
  input  [7:0]  io_pipe_phv_in_data_49,
  input  [7:0]  io_pipe_phv_in_data_50,
  input  [7:0]  io_pipe_phv_in_data_51,
  input  [7:0]  io_pipe_phv_in_data_52,
  input  [7:0]  io_pipe_phv_in_data_53,
  input  [7:0]  io_pipe_phv_in_data_54,
  input  [7:0]  io_pipe_phv_in_data_55,
  input  [7:0]  io_pipe_phv_in_data_56,
  input  [7:0]  io_pipe_phv_in_data_57,
  input  [7:0]  io_pipe_phv_in_data_58,
  input  [7:0]  io_pipe_phv_in_data_59,
  input  [7:0]  io_pipe_phv_in_data_60,
  input  [7:0]  io_pipe_phv_in_data_61,
  input  [7:0]  io_pipe_phv_in_data_62,
  input  [7:0]  io_pipe_phv_in_data_63,
  input  [7:0]  io_pipe_phv_in_data_64,
  input  [7:0]  io_pipe_phv_in_data_65,
  input  [7:0]  io_pipe_phv_in_data_66,
  input  [7:0]  io_pipe_phv_in_data_67,
  input  [7:0]  io_pipe_phv_in_data_68,
  input  [7:0]  io_pipe_phv_in_data_69,
  input  [7:0]  io_pipe_phv_in_data_70,
  input  [7:0]  io_pipe_phv_in_data_71,
  input  [7:0]  io_pipe_phv_in_data_72,
  input  [7:0]  io_pipe_phv_in_data_73,
  input  [7:0]  io_pipe_phv_in_data_74,
  input  [7:0]  io_pipe_phv_in_data_75,
  input  [7:0]  io_pipe_phv_in_data_76,
  input  [7:0]  io_pipe_phv_in_data_77,
  input  [7:0]  io_pipe_phv_in_data_78,
  input  [7:0]  io_pipe_phv_in_data_79,
  input  [7:0]  io_pipe_phv_in_data_80,
  input  [7:0]  io_pipe_phv_in_data_81,
  input  [7:0]  io_pipe_phv_in_data_82,
  input  [7:0]  io_pipe_phv_in_data_83,
  input  [7:0]  io_pipe_phv_in_data_84,
  input  [7:0]  io_pipe_phv_in_data_85,
  input  [7:0]  io_pipe_phv_in_data_86,
  input  [7:0]  io_pipe_phv_in_data_87,
  input  [7:0]  io_pipe_phv_in_data_88,
  input  [7:0]  io_pipe_phv_in_data_89,
  input  [7:0]  io_pipe_phv_in_data_90,
  input  [7:0]  io_pipe_phv_in_data_91,
  input  [7:0]  io_pipe_phv_in_data_92,
  input  [7:0]  io_pipe_phv_in_data_93,
  input  [7:0]  io_pipe_phv_in_data_94,
  input  [7:0]  io_pipe_phv_in_data_95,
  input  [7:0]  io_pipe_phv_in_data_96,
  input  [7:0]  io_pipe_phv_in_data_97,
  input  [7:0]  io_pipe_phv_in_data_98,
  input  [7:0]  io_pipe_phv_in_data_99,
  input  [7:0]  io_pipe_phv_in_data_100,
  input  [7:0]  io_pipe_phv_in_data_101,
  input  [7:0]  io_pipe_phv_in_data_102,
  input  [7:0]  io_pipe_phv_in_data_103,
  input  [7:0]  io_pipe_phv_in_data_104,
  input  [7:0]  io_pipe_phv_in_data_105,
  input  [7:0]  io_pipe_phv_in_data_106,
  input  [7:0]  io_pipe_phv_in_data_107,
  input  [7:0]  io_pipe_phv_in_data_108,
  input  [7:0]  io_pipe_phv_in_data_109,
  input  [7:0]  io_pipe_phv_in_data_110,
  input  [7:0]  io_pipe_phv_in_data_111,
  input  [7:0]  io_pipe_phv_in_data_112,
  input  [7:0]  io_pipe_phv_in_data_113,
  input  [7:0]  io_pipe_phv_in_data_114,
  input  [7:0]  io_pipe_phv_in_data_115,
  input  [7:0]  io_pipe_phv_in_data_116,
  input  [7:0]  io_pipe_phv_in_data_117,
  input  [7:0]  io_pipe_phv_in_data_118,
  input  [7:0]  io_pipe_phv_in_data_119,
  input  [7:0]  io_pipe_phv_in_data_120,
  input  [7:0]  io_pipe_phv_in_data_121,
  input  [7:0]  io_pipe_phv_in_data_122,
  input  [7:0]  io_pipe_phv_in_data_123,
  input  [7:0]  io_pipe_phv_in_data_124,
  input  [7:0]  io_pipe_phv_in_data_125,
  input  [7:0]  io_pipe_phv_in_data_126,
  input  [7:0]  io_pipe_phv_in_data_127,
  input  [7:0]  io_pipe_phv_in_data_128,
  input  [7:0]  io_pipe_phv_in_data_129,
  input  [7:0]  io_pipe_phv_in_data_130,
  input  [7:0]  io_pipe_phv_in_data_131,
  input  [7:0]  io_pipe_phv_in_data_132,
  input  [7:0]  io_pipe_phv_in_data_133,
  input  [7:0]  io_pipe_phv_in_data_134,
  input  [7:0]  io_pipe_phv_in_data_135,
  input  [7:0]  io_pipe_phv_in_data_136,
  input  [7:0]  io_pipe_phv_in_data_137,
  input  [7:0]  io_pipe_phv_in_data_138,
  input  [7:0]  io_pipe_phv_in_data_139,
  input  [7:0]  io_pipe_phv_in_data_140,
  input  [7:0]  io_pipe_phv_in_data_141,
  input  [7:0]  io_pipe_phv_in_data_142,
  input  [7:0]  io_pipe_phv_in_data_143,
  input  [7:0]  io_pipe_phv_in_data_144,
  input  [7:0]  io_pipe_phv_in_data_145,
  input  [7:0]  io_pipe_phv_in_data_146,
  input  [7:0]  io_pipe_phv_in_data_147,
  input  [7:0]  io_pipe_phv_in_data_148,
  input  [7:0]  io_pipe_phv_in_data_149,
  input  [7:0]  io_pipe_phv_in_data_150,
  input  [7:0]  io_pipe_phv_in_data_151,
  input  [7:0]  io_pipe_phv_in_data_152,
  input  [7:0]  io_pipe_phv_in_data_153,
  input  [7:0]  io_pipe_phv_in_data_154,
  input  [7:0]  io_pipe_phv_in_data_155,
  input  [7:0]  io_pipe_phv_in_data_156,
  input  [7:0]  io_pipe_phv_in_data_157,
  input  [7:0]  io_pipe_phv_in_data_158,
  input  [7:0]  io_pipe_phv_in_data_159,
  input  [7:0]  io_pipe_phv_in_data_160,
  input  [7:0]  io_pipe_phv_in_data_161,
  input  [7:0]  io_pipe_phv_in_data_162,
  input  [7:0]  io_pipe_phv_in_data_163,
  input  [7:0]  io_pipe_phv_in_data_164,
  input  [7:0]  io_pipe_phv_in_data_165,
  input  [7:0]  io_pipe_phv_in_data_166,
  input  [7:0]  io_pipe_phv_in_data_167,
  input  [7:0]  io_pipe_phv_in_data_168,
  input  [7:0]  io_pipe_phv_in_data_169,
  input  [7:0]  io_pipe_phv_in_data_170,
  input  [7:0]  io_pipe_phv_in_data_171,
  input  [7:0]  io_pipe_phv_in_data_172,
  input  [7:0]  io_pipe_phv_in_data_173,
  input  [7:0]  io_pipe_phv_in_data_174,
  input  [7:0]  io_pipe_phv_in_data_175,
  input  [7:0]  io_pipe_phv_in_data_176,
  input  [7:0]  io_pipe_phv_in_data_177,
  input  [7:0]  io_pipe_phv_in_data_178,
  input  [7:0]  io_pipe_phv_in_data_179,
  input  [7:0]  io_pipe_phv_in_data_180,
  input  [7:0]  io_pipe_phv_in_data_181,
  input  [7:0]  io_pipe_phv_in_data_182,
  input  [7:0]  io_pipe_phv_in_data_183,
  input  [7:0]  io_pipe_phv_in_data_184,
  input  [7:0]  io_pipe_phv_in_data_185,
  input  [7:0]  io_pipe_phv_in_data_186,
  input  [7:0]  io_pipe_phv_in_data_187,
  input  [7:0]  io_pipe_phv_in_data_188,
  input  [7:0]  io_pipe_phv_in_data_189,
  input  [7:0]  io_pipe_phv_in_data_190,
  input  [7:0]  io_pipe_phv_in_data_191,
  input  [7:0]  io_pipe_phv_in_data_192,
  input  [7:0]  io_pipe_phv_in_data_193,
  input  [7:0]  io_pipe_phv_in_data_194,
  input  [7:0]  io_pipe_phv_in_data_195,
  input  [7:0]  io_pipe_phv_in_data_196,
  input  [7:0]  io_pipe_phv_in_data_197,
  input  [7:0]  io_pipe_phv_in_data_198,
  input  [7:0]  io_pipe_phv_in_data_199,
  input  [7:0]  io_pipe_phv_in_data_200,
  input  [7:0]  io_pipe_phv_in_data_201,
  input  [7:0]  io_pipe_phv_in_data_202,
  input  [7:0]  io_pipe_phv_in_data_203,
  input  [7:0]  io_pipe_phv_in_data_204,
  input  [7:0]  io_pipe_phv_in_data_205,
  input  [7:0]  io_pipe_phv_in_data_206,
  input  [7:0]  io_pipe_phv_in_data_207,
  input  [7:0]  io_pipe_phv_in_data_208,
  input  [7:0]  io_pipe_phv_in_data_209,
  input  [7:0]  io_pipe_phv_in_data_210,
  input  [7:0]  io_pipe_phv_in_data_211,
  input  [7:0]  io_pipe_phv_in_data_212,
  input  [7:0]  io_pipe_phv_in_data_213,
  input  [7:0]  io_pipe_phv_in_data_214,
  input  [7:0]  io_pipe_phv_in_data_215,
  input  [7:0]  io_pipe_phv_in_data_216,
  input  [7:0]  io_pipe_phv_in_data_217,
  input  [7:0]  io_pipe_phv_in_data_218,
  input  [7:0]  io_pipe_phv_in_data_219,
  input  [7:0]  io_pipe_phv_in_data_220,
  input  [7:0]  io_pipe_phv_in_data_221,
  input  [7:0]  io_pipe_phv_in_data_222,
  input  [7:0]  io_pipe_phv_in_data_223,
  input  [7:0]  io_pipe_phv_in_data_224,
  input  [7:0]  io_pipe_phv_in_data_225,
  input  [7:0]  io_pipe_phv_in_data_226,
  input  [7:0]  io_pipe_phv_in_data_227,
  input  [7:0]  io_pipe_phv_in_data_228,
  input  [7:0]  io_pipe_phv_in_data_229,
  input  [7:0]  io_pipe_phv_in_data_230,
  input  [7:0]  io_pipe_phv_in_data_231,
  input  [7:0]  io_pipe_phv_in_data_232,
  input  [7:0]  io_pipe_phv_in_data_233,
  input  [7:0]  io_pipe_phv_in_data_234,
  input  [7:0]  io_pipe_phv_in_data_235,
  input  [7:0]  io_pipe_phv_in_data_236,
  input  [7:0]  io_pipe_phv_in_data_237,
  input  [7:0]  io_pipe_phv_in_data_238,
  input  [7:0]  io_pipe_phv_in_data_239,
  input  [7:0]  io_pipe_phv_in_data_240,
  input  [7:0]  io_pipe_phv_in_data_241,
  input  [7:0]  io_pipe_phv_in_data_242,
  input  [7:0]  io_pipe_phv_in_data_243,
  input  [7:0]  io_pipe_phv_in_data_244,
  input  [7:0]  io_pipe_phv_in_data_245,
  input  [7:0]  io_pipe_phv_in_data_246,
  input  [7:0]  io_pipe_phv_in_data_247,
  input  [7:0]  io_pipe_phv_in_data_248,
  input  [7:0]  io_pipe_phv_in_data_249,
  input  [7:0]  io_pipe_phv_in_data_250,
  input  [7:0]  io_pipe_phv_in_data_251,
  input  [7:0]  io_pipe_phv_in_data_252,
  input  [7:0]  io_pipe_phv_in_data_253,
  input  [7:0]  io_pipe_phv_in_data_254,
  input  [7:0]  io_pipe_phv_in_data_255,
  input  [3:0]  io_pipe_phv_in_next_processor_id,
  input         io_pipe_phv_in_next_config_id,
  input         io_pipe_phv_in_is_valid_processor,
  output [7:0]  io_pipe_phv_out_data_0,
  output [7:0]  io_pipe_phv_out_data_1,
  output [7:0]  io_pipe_phv_out_data_2,
  output [7:0]  io_pipe_phv_out_data_3,
  output [7:0]  io_pipe_phv_out_data_4,
  output [7:0]  io_pipe_phv_out_data_5,
  output [7:0]  io_pipe_phv_out_data_6,
  output [7:0]  io_pipe_phv_out_data_7,
  output [7:0]  io_pipe_phv_out_data_8,
  output [7:0]  io_pipe_phv_out_data_9,
  output [7:0]  io_pipe_phv_out_data_10,
  output [7:0]  io_pipe_phv_out_data_11,
  output [7:0]  io_pipe_phv_out_data_12,
  output [7:0]  io_pipe_phv_out_data_13,
  output [7:0]  io_pipe_phv_out_data_14,
  output [7:0]  io_pipe_phv_out_data_15,
  output [7:0]  io_pipe_phv_out_data_16,
  output [7:0]  io_pipe_phv_out_data_17,
  output [7:0]  io_pipe_phv_out_data_18,
  output [7:0]  io_pipe_phv_out_data_19,
  output [7:0]  io_pipe_phv_out_data_20,
  output [7:0]  io_pipe_phv_out_data_21,
  output [7:0]  io_pipe_phv_out_data_22,
  output [7:0]  io_pipe_phv_out_data_23,
  output [7:0]  io_pipe_phv_out_data_24,
  output [7:0]  io_pipe_phv_out_data_25,
  output [7:0]  io_pipe_phv_out_data_26,
  output [7:0]  io_pipe_phv_out_data_27,
  output [7:0]  io_pipe_phv_out_data_28,
  output [7:0]  io_pipe_phv_out_data_29,
  output [7:0]  io_pipe_phv_out_data_30,
  output [7:0]  io_pipe_phv_out_data_31,
  output [7:0]  io_pipe_phv_out_data_32,
  output [7:0]  io_pipe_phv_out_data_33,
  output [7:0]  io_pipe_phv_out_data_34,
  output [7:0]  io_pipe_phv_out_data_35,
  output [7:0]  io_pipe_phv_out_data_36,
  output [7:0]  io_pipe_phv_out_data_37,
  output [7:0]  io_pipe_phv_out_data_38,
  output [7:0]  io_pipe_phv_out_data_39,
  output [7:0]  io_pipe_phv_out_data_40,
  output [7:0]  io_pipe_phv_out_data_41,
  output [7:0]  io_pipe_phv_out_data_42,
  output [7:0]  io_pipe_phv_out_data_43,
  output [7:0]  io_pipe_phv_out_data_44,
  output [7:0]  io_pipe_phv_out_data_45,
  output [7:0]  io_pipe_phv_out_data_46,
  output [7:0]  io_pipe_phv_out_data_47,
  output [7:0]  io_pipe_phv_out_data_48,
  output [7:0]  io_pipe_phv_out_data_49,
  output [7:0]  io_pipe_phv_out_data_50,
  output [7:0]  io_pipe_phv_out_data_51,
  output [7:0]  io_pipe_phv_out_data_52,
  output [7:0]  io_pipe_phv_out_data_53,
  output [7:0]  io_pipe_phv_out_data_54,
  output [7:0]  io_pipe_phv_out_data_55,
  output [7:0]  io_pipe_phv_out_data_56,
  output [7:0]  io_pipe_phv_out_data_57,
  output [7:0]  io_pipe_phv_out_data_58,
  output [7:0]  io_pipe_phv_out_data_59,
  output [7:0]  io_pipe_phv_out_data_60,
  output [7:0]  io_pipe_phv_out_data_61,
  output [7:0]  io_pipe_phv_out_data_62,
  output [7:0]  io_pipe_phv_out_data_63,
  output [7:0]  io_pipe_phv_out_data_64,
  output [7:0]  io_pipe_phv_out_data_65,
  output [7:0]  io_pipe_phv_out_data_66,
  output [7:0]  io_pipe_phv_out_data_67,
  output [7:0]  io_pipe_phv_out_data_68,
  output [7:0]  io_pipe_phv_out_data_69,
  output [7:0]  io_pipe_phv_out_data_70,
  output [7:0]  io_pipe_phv_out_data_71,
  output [7:0]  io_pipe_phv_out_data_72,
  output [7:0]  io_pipe_phv_out_data_73,
  output [7:0]  io_pipe_phv_out_data_74,
  output [7:0]  io_pipe_phv_out_data_75,
  output [7:0]  io_pipe_phv_out_data_76,
  output [7:0]  io_pipe_phv_out_data_77,
  output [7:0]  io_pipe_phv_out_data_78,
  output [7:0]  io_pipe_phv_out_data_79,
  output [7:0]  io_pipe_phv_out_data_80,
  output [7:0]  io_pipe_phv_out_data_81,
  output [7:0]  io_pipe_phv_out_data_82,
  output [7:0]  io_pipe_phv_out_data_83,
  output [7:0]  io_pipe_phv_out_data_84,
  output [7:0]  io_pipe_phv_out_data_85,
  output [7:0]  io_pipe_phv_out_data_86,
  output [7:0]  io_pipe_phv_out_data_87,
  output [7:0]  io_pipe_phv_out_data_88,
  output [7:0]  io_pipe_phv_out_data_89,
  output [7:0]  io_pipe_phv_out_data_90,
  output [7:0]  io_pipe_phv_out_data_91,
  output [7:0]  io_pipe_phv_out_data_92,
  output [7:0]  io_pipe_phv_out_data_93,
  output [7:0]  io_pipe_phv_out_data_94,
  output [7:0]  io_pipe_phv_out_data_95,
  output [7:0]  io_pipe_phv_out_data_96,
  output [7:0]  io_pipe_phv_out_data_97,
  output [7:0]  io_pipe_phv_out_data_98,
  output [7:0]  io_pipe_phv_out_data_99,
  output [7:0]  io_pipe_phv_out_data_100,
  output [7:0]  io_pipe_phv_out_data_101,
  output [7:0]  io_pipe_phv_out_data_102,
  output [7:0]  io_pipe_phv_out_data_103,
  output [7:0]  io_pipe_phv_out_data_104,
  output [7:0]  io_pipe_phv_out_data_105,
  output [7:0]  io_pipe_phv_out_data_106,
  output [7:0]  io_pipe_phv_out_data_107,
  output [7:0]  io_pipe_phv_out_data_108,
  output [7:0]  io_pipe_phv_out_data_109,
  output [7:0]  io_pipe_phv_out_data_110,
  output [7:0]  io_pipe_phv_out_data_111,
  output [7:0]  io_pipe_phv_out_data_112,
  output [7:0]  io_pipe_phv_out_data_113,
  output [7:0]  io_pipe_phv_out_data_114,
  output [7:0]  io_pipe_phv_out_data_115,
  output [7:0]  io_pipe_phv_out_data_116,
  output [7:0]  io_pipe_phv_out_data_117,
  output [7:0]  io_pipe_phv_out_data_118,
  output [7:0]  io_pipe_phv_out_data_119,
  output [7:0]  io_pipe_phv_out_data_120,
  output [7:0]  io_pipe_phv_out_data_121,
  output [7:0]  io_pipe_phv_out_data_122,
  output [7:0]  io_pipe_phv_out_data_123,
  output [7:0]  io_pipe_phv_out_data_124,
  output [7:0]  io_pipe_phv_out_data_125,
  output [7:0]  io_pipe_phv_out_data_126,
  output [7:0]  io_pipe_phv_out_data_127,
  output [7:0]  io_pipe_phv_out_data_128,
  output [7:0]  io_pipe_phv_out_data_129,
  output [7:0]  io_pipe_phv_out_data_130,
  output [7:0]  io_pipe_phv_out_data_131,
  output [7:0]  io_pipe_phv_out_data_132,
  output [7:0]  io_pipe_phv_out_data_133,
  output [7:0]  io_pipe_phv_out_data_134,
  output [7:0]  io_pipe_phv_out_data_135,
  output [7:0]  io_pipe_phv_out_data_136,
  output [7:0]  io_pipe_phv_out_data_137,
  output [7:0]  io_pipe_phv_out_data_138,
  output [7:0]  io_pipe_phv_out_data_139,
  output [7:0]  io_pipe_phv_out_data_140,
  output [7:0]  io_pipe_phv_out_data_141,
  output [7:0]  io_pipe_phv_out_data_142,
  output [7:0]  io_pipe_phv_out_data_143,
  output [7:0]  io_pipe_phv_out_data_144,
  output [7:0]  io_pipe_phv_out_data_145,
  output [7:0]  io_pipe_phv_out_data_146,
  output [7:0]  io_pipe_phv_out_data_147,
  output [7:0]  io_pipe_phv_out_data_148,
  output [7:0]  io_pipe_phv_out_data_149,
  output [7:0]  io_pipe_phv_out_data_150,
  output [7:0]  io_pipe_phv_out_data_151,
  output [7:0]  io_pipe_phv_out_data_152,
  output [7:0]  io_pipe_phv_out_data_153,
  output [7:0]  io_pipe_phv_out_data_154,
  output [7:0]  io_pipe_phv_out_data_155,
  output [7:0]  io_pipe_phv_out_data_156,
  output [7:0]  io_pipe_phv_out_data_157,
  output [7:0]  io_pipe_phv_out_data_158,
  output [7:0]  io_pipe_phv_out_data_159,
  output [7:0]  io_pipe_phv_out_data_160,
  output [7:0]  io_pipe_phv_out_data_161,
  output [7:0]  io_pipe_phv_out_data_162,
  output [7:0]  io_pipe_phv_out_data_163,
  output [7:0]  io_pipe_phv_out_data_164,
  output [7:0]  io_pipe_phv_out_data_165,
  output [7:0]  io_pipe_phv_out_data_166,
  output [7:0]  io_pipe_phv_out_data_167,
  output [7:0]  io_pipe_phv_out_data_168,
  output [7:0]  io_pipe_phv_out_data_169,
  output [7:0]  io_pipe_phv_out_data_170,
  output [7:0]  io_pipe_phv_out_data_171,
  output [7:0]  io_pipe_phv_out_data_172,
  output [7:0]  io_pipe_phv_out_data_173,
  output [7:0]  io_pipe_phv_out_data_174,
  output [7:0]  io_pipe_phv_out_data_175,
  output [7:0]  io_pipe_phv_out_data_176,
  output [7:0]  io_pipe_phv_out_data_177,
  output [7:0]  io_pipe_phv_out_data_178,
  output [7:0]  io_pipe_phv_out_data_179,
  output [7:0]  io_pipe_phv_out_data_180,
  output [7:0]  io_pipe_phv_out_data_181,
  output [7:0]  io_pipe_phv_out_data_182,
  output [7:0]  io_pipe_phv_out_data_183,
  output [7:0]  io_pipe_phv_out_data_184,
  output [7:0]  io_pipe_phv_out_data_185,
  output [7:0]  io_pipe_phv_out_data_186,
  output [7:0]  io_pipe_phv_out_data_187,
  output [7:0]  io_pipe_phv_out_data_188,
  output [7:0]  io_pipe_phv_out_data_189,
  output [7:0]  io_pipe_phv_out_data_190,
  output [7:0]  io_pipe_phv_out_data_191,
  output [7:0]  io_pipe_phv_out_data_192,
  output [7:0]  io_pipe_phv_out_data_193,
  output [7:0]  io_pipe_phv_out_data_194,
  output [7:0]  io_pipe_phv_out_data_195,
  output [7:0]  io_pipe_phv_out_data_196,
  output [7:0]  io_pipe_phv_out_data_197,
  output [7:0]  io_pipe_phv_out_data_198,
  output [7:0]  io_pipe_phv_out_data_199,
  output [7:0]  io_pipe_phv_out_data_200,
  output [7:0]  io_pipe_phv_out_data_201,
  output [7:0]  io_pipe_phv_out_data_202,
  output [7:0]  io_pipe_phv_out_data_203,
  output [7:0]  io_pipe_phv_out_data_204,
  output [7:0]  io_pipe_phv_out_data_205,
  output [7:0]  io_pipe_phv_out_data_206,
  output [7:0]  io_pipe_phv_out_data_207,
  output [7:0]  io_pipe_phv_out_data_208,
  output [7:0]  io_pipe_phv_out_data_209,
  output [7:0]  io_pipe_phv_out_data_210,
  output [7:0]  io_pipe_phv_out_data_211,
  output [7:0]  io_pipe_phv_out_data_212,
  output [7:0]  io_pipe_phv_out_data_213,
  output [7:0]  io_pipe_phv_out_data_214,
  output [7:0]  io_pipe_phv_out_data_215,
  output [7:0]  io_pipe_phv_out_data_216,
  output [7:0]  io_pipe_phv_out_data_217,
  output [7:0]  io_pipe_phv_out_data_218,
  output [7:0]  io_pipe_phv_out_data_219,
  output [7:0]  io_pipe_phv_out_data_220,
  output [7:0]  io_pipe_phv_out_data_221,
  output [7:0]  io_pipe_phv_out_data_222,
  output [7:0]  io_pipe_phv_out_data_223,
  output [7:0]  io_pipe_phv_out_data_224,
  output [7:0]  io_pipe_phv_out_data_225,
  output [7:0]  io_pipe_phv_out_data_226,
  output [7:0]  io_pipe_phv_out_data_227,
  output [7:0]  io_pipe_phv_out_data_228,
  output [7:0]  io_pipe_phv_out_data_229,
  output [7:0]  io_pipe_phv_out_data_230,
  output [7:0]  io_pipe_phv_out_data_231,
  output [7:0]  io_pipe_phv_out_data_232,
  output [7:0]  io_pipe_phv_out_data_233,
  output [7:0]  io_pipe_phv_out_data_234,
  output [7:0]  io_pipe_phv_out_data_235,
  output [7:0]  io_pipe_phv_out_data_236,
  output [7:0]  io_pipe_phv_out_data_237,
  output [7:0]  io_pipe_phv_out_data_238,
  output [7:0]  io_pipe_phv_out_data_239,
  output [7:0]  io_pipe_phv_out_data_240,
  output [7:0]  io_pipe_phv_out_data_241,
  output [7:0]  io_pipe_phv_out_data_242,
  output [7:0]  io_pipe_phv_out_data_243,
  output [7:0]  io_pipe_phv_out_data_244,
  output [7:0]  io_pipe_phv_out_data_245,
  output [7:0]  io_pipe_phv_out_data_246,
  output [7:0]  io_pipe_phv_out_data_247,
  output [7:0]  io_pipe_phv_out_data_248,
  output [7:0]  io_pipe_phv_out_data_249,
  output [7:0]  io_pipe_phv_out_data_250,
  output [7:0]  io_pipe_phv_out_data_251,
  output [7:0]  io_pipe_phv_out_data_252,
  output [7:0]  io_pipe_phv_out_data_253,
  output [7:0]  io_pipe_phv_out_data_254,
  output [7:0]  io_pipe_phv_out_data_255,
  output [3:0]  io_pipe_phv_out_next_processor_id,
  output        io_pipe_phv_out_next_config_id,
  output        io_pipe_phv_out_is_valid_processor,
  input         io_mod_en,
  input         io_mod_config_id,
  input         io_mod_key_mod_en,
  input  [2:0]  io_mod_key_mod_group_index,
  input  [1:0]  io_mod_key_mod_group_config,
  input         io_mod_key_mod_group_mask_0,
  input         io_mod_key_mod_group_mask_1,
  input         io_mod_key_mod_group_mask_2,
  input         io_mod_key_mod_group_mask_3,
  input  [7:0]  io_mod_key_mod_group_id_0,
  input  [7:0]  io_mod_key_mod_group_id_1,
  input  [7:0]  io_mod_key_mod_group_id_2,
  input  [7:0]  io_mod_key_mod_group_id_3,
  input  [4:0]  io_mod_table_mod_table_depth,
  input  [4:0]  io_mod_table_mod_table_width,
  input         io_mod_w_en,
  input  [3:0]  io_mod_w_sram_id,
  input  [7:0]  io_mod_w_addr,
  input  [63:0] io_mod_w_data,
  output        io_hit,
  output [63:0] io_match_value
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
`endif // RANDOMIZE_REG_INIT
  wire  pipe1_clock; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_0; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_1; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_2; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_3; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_4; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_5; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_6; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_7; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_8; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_9; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_10; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_11; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_12; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_13; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_14; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_15; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_16; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_17; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_18; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_19; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_20; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_21; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_22; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_23; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_24; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_25; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_26; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_27; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_28; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_29; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_30; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_31; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_32; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_33; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_34; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_35; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_36; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_37; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_38; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_39; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_40; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_41; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_42; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_43; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_44; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_45; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_46; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_47; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_48; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_49; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_50; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_51; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_52; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_53; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_54; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_55; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_56; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_57; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_58; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_59; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_60; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_61; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_62; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_63; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_64; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_65; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_66; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_67; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_68; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_69; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_70; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_71; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_72; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_73; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_74; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_75; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_76; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_77; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_78; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_79; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_80; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_81; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_82; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_83; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_84; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_85; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_86; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_87; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_88; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_89; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_90; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_91; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_92; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_93; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_94; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_95; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_96; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_97; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_98; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_99; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_100; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_101; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_102; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_103; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_104; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_105; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_106; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_107; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_108; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_109; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_110; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_111; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_112; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_113; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_114; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_115; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_116; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_117; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_118; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_119; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_120; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_121; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_122; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_123; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_124; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_125; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_126; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_127; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_128; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_129; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_130; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_131; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_132; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_133; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_134; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_135; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_136; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_137; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_138; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_139; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_140; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_141; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_142; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_143; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_144; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_145; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_146; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_147; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_148; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_149; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_150; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_151; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_152; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_153; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_154; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_155; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_156; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_157; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_158; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_159; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_160; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_161; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_162; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_163; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_164; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_165; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_166; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_167; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_168; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_169; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_170; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_171; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_172; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_173; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_174; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_175; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_176; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_177; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_178; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_179; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_180; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_181; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_182; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_183; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_184; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_185; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_186; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_187; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_188; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_189; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_190; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_191; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_192; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_193; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_194; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_195; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_196; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_197; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_198; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_199; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_200; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_201; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_202; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_203; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_204; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_205; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_206; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_207; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_208; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_209; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_210; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_211; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_212; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_213; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_214; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_215; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_216; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_217; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_218; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_219; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_220; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_221; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_222; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_223; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_224; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_225; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_226; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_227; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_228; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_229; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_230; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_231; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_232; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_233; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_234; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_235; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_236; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_237; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_238; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_239; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_240; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_241; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_242; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_243; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_244; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_245; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_246; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_247; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_248; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_249; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_250; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_251; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_252; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_253; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_254; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_255; // @[matcher_pisa.scala 333:23]
  wire [3:0] pipe1_io_pipe_phv_in_next_processor_id; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_pipe_phv_in_next_config_id; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_pipe_phv_in_is_valid_processor; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_0; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_1; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_2; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_3; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_4; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_5; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_6; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_7; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_8; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_9; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_10; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_11; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_12; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_13; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_14; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_15; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_16; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_17; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_18; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_19; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_20; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_21; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_22; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_23; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_24; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_25; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_26; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_27; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_28; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_29; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_30; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_31; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_32; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_33; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_34; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_35; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_36; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_37; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_38; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_39; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_40; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_41; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_42; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_43; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_44; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_45; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_46; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_47; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_48; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_49; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_50; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_51; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_52; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_53; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_54; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_55; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_56; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_57; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_58; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_59; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_60; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_61; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_62; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_63; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_64; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_65; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_66; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_67; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_68; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_69; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_70; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_71; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_72; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_73; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_74; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_75; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_76; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_77; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_78; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_79; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_80; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_81; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_82; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_83; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_84; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_85; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_86; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_87; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_88; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_89; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_90; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_91; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_92; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_93; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_94; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_95; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_96; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_97; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_98; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_99; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_100; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_101; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_102; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_103; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_104; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_105; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_106; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_107; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_108; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_109; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_110; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_111; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_112; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_113; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_114; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_115; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_116; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_117; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_118; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_119; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_120; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_121; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_122; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_123; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_124; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_125; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_126; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_127; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_128; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_129; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_130; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_131; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_132; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_133; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_134; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_135; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_136; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_137; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_138; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_139; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_140; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_141; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_142; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_143; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_144; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_145; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_146; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_147; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_148; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_149; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_150; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_151; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_152; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_153; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_154; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_155; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_156; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_157; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_158; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_159; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_160; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_161; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_162; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_163; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_164; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_165; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_166; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_167; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_168; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_169; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_170; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_171; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_172; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_173; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_174; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_175; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_176; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_177; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_178; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_179; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_180; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_181; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_182; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_183; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_184; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_185; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_186; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_187; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_188; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_189; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_190; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_191; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_192; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_193; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_194; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_195; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_196; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_197; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_198; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_199; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_200; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_201; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_202; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_203; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_204; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_205; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_206; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_207; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_208; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_209; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_210; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_211; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_212; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_213; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_214; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_215; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_216; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_217; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_218; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_219; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_220; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_221; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_222; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_223; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_224; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_225; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_226; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_227; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_228; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_229; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_230; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_231; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_232; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_233; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_234; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_235; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_236; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_237; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_238; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_239; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_240; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_241; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_242; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_243; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_244; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_245; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_246; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_247; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_248; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_249; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_250; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_251; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_252; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_253; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_254; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_255; // @[matcher_pisa.scala 333:23]
  wire [3:0] pipe1_io_pipe_phv_out_next_processor_id; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_pipe_phv_out_next_config_id; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_pipe_phv_out_is_valid_processor; // @[matcher_pisa.scala 333:23]
  wire [1:0] pipe1_io_key_config_0_field_config_0; // @[matcher_pisa.scala 333:23]
  wire [1:0] pipe1_io_key_config_0_field_config_1; // @[matcher_pisa.scala 333:23]
  wire [1:0] pipe1_io_key_config_0_field_config_2; // @[matcher_pisa.scala 333:23]
  wire [1:0] pipe1_io_key_config_0_field_config_3; // @[matcher_pisa.scala 333:23]
  wire [1:0] pipe1_io_key_config_0_field_config_4; // @[matcher_pisa.scala 333:23]
  wire [1:0] pipe1_io_key_config_0_field_config_5; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_0_field_mask_0_0; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_0_field_mask_0_1; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_0_field_mask_0_2; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_0_field_mask_0_3; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_0_field_mask_1_0; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_0_field_mask_1_1; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_0_field_mask_1_2; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_0_field_mask_1_3; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_0_field_mask_2_0; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_0_field_mask_2_1; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_0_field_mask_2_2; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_0_field_mask_2_3; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_0_field_mask_3_0; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_0_field_mask_3_1; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_0_field_mask_3_2; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_0_field_mask_3_3; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_0_field_mask_4_0; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_0_field_mask_4_1; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_0_field_mask_4_2; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_0_field_mask_4_3; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_0_field_mask_5_0; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_0_field_mask_5_1; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_0_field_mask_5_2; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_0_field_mask_5_3; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_0_field_id_0_0; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_0_field_id_0_1; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_0_field_id_0_2; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_0_field_id_0_3; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_0_field_id_1_0; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_0_field_id_1_1; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_0_field_id_1_2; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_0_field_id_1_3; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_0_field_id_2_0; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_0_field_id_2_1; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_0_field_id_2_2; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_0_field_id_2_3; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_0_field_id_3_0; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_0_field_id_3_1; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_0_field_id_3_2; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_0_field_id_3_3; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_0_field_id_4_0; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_0_field_id_4_1; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_0_field_id_4_2; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_0_field_id_4_3; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_0_field_id_5_0; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_0_field_id_5_1; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_0_field_id_5_2; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_0_field_id_5_3; // @[matcher_pisa.scala 333:23]
  wire [1:0] pipe1_io_key_config_1_field_config_0; // @[matcher_pisa.scala 333:23]
  wire [1:0] pipe1_io_key_config_1_field_config_1; // @[matcher_pisa.scala 333:23]
  wire [1:0] pipe1_io_key_config_1_field_config_2; // @[matcher_pisa.scala 333:23]
  wire [1:0] pipe1_io_key_config_1_field_config_3; // @[matcher_pisa.scala 333:23]
  wire [1:0] pipe1_io_key_config_1_field_config_4; // @[matcher_pisa.scala 333:23]
  wire [1:0] pipe1_io_key_config_1_field_config_5; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_1_field_mask_0_0; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_1_field_mask_0_1; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_1_field_mask_0_2; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_1_field_mask_0_3; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_1_field_mask_1_0; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_1_field_mask_1_1; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_1_field_mask_1_2; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_1_field_mask_1_3; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_1_field_mask_2_0; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_1_field_mask_2_1; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_1_field_mask_2_2; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_1_field_mask_2_3; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_1_field_mask_3_0; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_1_field_mask_3_1; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_1_field_mask_3_2; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_1_field_mask_3_3; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_1_field_mask_4_0; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_1_field_mask_4_1; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_1_field_mask_4_2; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_1_field_mask_4_3; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_1_field_mask_5_0; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_1_field_mask_5_1; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_1_field_mask_5_2; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_1_field_mask_5_3; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_1_field_id_0_0; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_1_field_id_0_1; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_1_field_id_0_2; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_1_field_id_0_3; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_1_field_id_1_0; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_1_field_id_1_1; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_1_field_id_1_2; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_1_field_id_1_3; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_1_field_id_2_0; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_1_field_id_2_1; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_1_field_id_2_2; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_1_field_id_2_3; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_1_field_id_3_0; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_1_field_id_3_1; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_1_field_id_3_2; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_1_field_id_3_3; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_1_field_id_4_0; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_1_field_id_4_1; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_1_field_id_4_2; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_1_field_id_4_3; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_1_field_id_5_0; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_1_field_id_5_1; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_1_field_id_5_2; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_1_field_id_5_3; // @[matcher_pisa.scala 333:23]
  wire [191:0] pipe1_io_match_key; // @[matcher_pisa.scala 333:23]
  wire  pipe2_clock; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_0; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_1; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_2; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_3; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_4; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_5; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_6; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_7; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_8; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_9; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_10; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_11; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_12; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_13; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_14; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_15; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_16; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_17; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_18; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_19; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_20; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_21; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_22; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_23; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_24; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_25; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_26; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_27; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_28; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_29; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_30; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_31; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_32; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_33; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_34; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_35; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_36; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_37; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_38; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_39; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_40; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_41; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_42; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_43; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_44; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_45; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_46; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_47; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_48; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_49; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_50; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_51; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_52; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_53; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_54; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_55; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_56; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_57; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_58; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_59; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_60; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_61; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_62; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_63; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_64; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_65; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_66; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_67; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_68; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_69; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_70; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_71; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_72; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_73; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_74; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_75; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_76; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_77; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_78; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_79; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_80; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_81; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_82; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_83; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_84; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_85; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_86; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_87; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_88; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_89; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_90; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_91; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_92; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_93; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_94; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_95; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_96; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_97; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_98; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_99; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_100; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_101; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_102; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_103; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_104; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_105; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_106; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_107; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_108; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_109; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_110; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_111; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_112; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_113; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_114; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_115; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_116; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_117; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_118; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_119; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_120; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_121; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_122; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_123; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_124; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_125; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_126; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_127; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_128; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_129; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_130; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_131; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_132; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_133; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_134; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_135; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_136; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_137; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_138; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_139; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_140; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_141; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_142; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_143; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_144; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_145; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_146; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_147; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_148; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_149; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_150; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_151; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_152; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_153; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_154; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_155; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_156; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_157; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_158; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_159; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_160; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_161; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_162; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_163; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_164; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_165; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_166; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_167; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_168; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_169; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_170; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_171; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_172; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_173; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_174; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_175; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_176; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_177; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_178; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_179; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_180; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_181; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_182; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_183; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_184; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_185; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_186; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_187; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_188; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_189; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_190; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_191; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_192; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_193; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_194; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_195; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_196; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_197; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_198; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_199; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_200; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_201; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_202; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_203; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_204; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_205; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_206; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_207; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_208; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_209; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_210; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_211; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_212; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_213; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_214; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_215; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_216; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_217; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_218; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_219; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_220; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_221; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_222; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_223; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_224; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_225; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_226; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_227; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_228; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_229; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_230; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_231; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_232; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_233; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_234; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_235; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_236; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_237; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_238; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_239; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_240; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_241; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_242; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_243; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_244; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_245; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_246; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_247; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_248; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_249; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_250; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_251; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_252; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_253; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_254; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_255; // @[matcher_pisa.scala 334:23]
  wire [3:0] pipe2_io_pipe_phv_in_next_processor_id; // @[matcher_pisa.scala 334:23]
  wire  pipe2_io_pipe_phv_in_next_config_id; // @[matcher_pisa.scala 334:23]
  wire  pipe2_io_pipe_phv_in_is_valid_processor; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_0; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_1; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_2; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_3; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_4; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_5; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_6; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_7; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_8; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_9; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_10; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_11; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_12; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_13; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_14; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_15; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_16; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_17; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_18; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_19; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_20; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_21; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_22; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_23; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_24; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_25; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_26; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_27; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_28; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_29; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_30; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_31; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_32; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_33; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_34; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_35; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_36; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_37; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_38; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_39; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_40; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_41; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_42; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_43; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_44; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_45; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_46; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_47; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_48; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_49; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_50; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_51; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_52; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_53; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_54; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_55; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_56; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_57; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_58; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_59; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_60; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_61; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_62; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_63; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_64; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_65; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_66; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_67; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_68; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_69; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_70; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_71; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_72; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_73; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_74; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_75; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_76; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_77; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_78; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_79; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_80; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_81; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_82; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_83; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_84; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_85; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_86; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_87; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_88; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_89; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_90; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_91; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_92; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_93; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_94; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_95; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_96; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_97; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_98; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_99; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_100; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_101; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_102; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_103; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_104; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_105; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_106; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_107; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_108; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_109; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_110; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_111; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_112; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_113; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_114; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_115; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_116; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_117; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_118; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_119; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_120; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_121; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_122; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_123; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_124; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_125; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_126; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_127; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_128; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_129; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_130; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_131; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_132; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_133; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_134; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_135; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_136; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_137; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_138; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_139; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_140; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_141; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_142; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_143; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_144; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_145; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_146; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_147; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_148; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_149; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_150; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_151; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_152; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_153; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_154; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_155; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_156; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_157; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_158; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_159; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_160; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_161; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_162; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_163; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_164; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_165; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_166; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_167; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_168; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_169; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_170; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_171; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_172; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_173; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_174; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_175; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_176; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_177; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_178; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_179; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_180; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_181; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_182; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_183; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_184; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_185; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_186; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_187; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_188; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_189; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_190; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_191; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_192; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_193; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_194; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_195; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_196; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_197; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_198; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_199; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_200; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_201; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_202; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_203; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_204; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_205; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_206; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_207; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_208; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_209; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_210; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_211; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_212; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_213; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_214; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_215; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_216; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_217; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_218; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_219; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_220; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_221; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_222; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_223; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_224; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_225; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_226; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_227; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_228; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_229; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_230; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_231; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_232; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_233; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_234; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_235; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_236; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_237; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_238; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_239; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_240; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_241; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_242; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_243; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_244; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_245; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_246; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_247; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_248; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_249; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_250; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_251; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_252; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_253; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_254; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_255; // @[matcher_pisa.scala 334:23]
  wire [3:0] pipe2_io_pipe_phv_out_next_processor_id; // @[matcher_pisa.scala 334:23]
  wire  pipe2_io_pipe_phv_out_next_config_id; // @[matcher_pisa.scala 334:23]
  wire  pipe2_io_pipe_phv_out_is_valid_processor; // @[matcher_pisa.scala 334:23]
  wire  pipe2_io_mod_hash_depth_mod; // @[matcher_pisa.scala 334:23]
  wire  pipe2_io_mod_config_id; // @[matcher_pisa.scala 334:23]
  wire [3:0] pipe2_io_mod_hash_depth; // @[matcher_pisa.scala 334:23]
  wire [191:0] pipe2_io_key_in; // @[matcher_pisa.scala 334:23]
  wire [191:0] pipe2_io_key_out; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_hash_val; // @[matcher_pisa.scala 334:23]
  wire [3:0] pipe2_io_hash_val_cs; // @[matcher_pisa.scala 334:23]
  wire  pipe3_clock; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_0; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_1; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_2; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_3; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_4; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_5; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_6; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_7; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_8; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_9; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_10; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_11; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_12; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_13; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_14; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_15; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_16; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_17; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_18; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_19; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_20; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_21; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_22; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_23; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_24; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_25; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_26; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_27; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_28; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_29; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_30; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_31; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_32; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_33; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_34; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_35; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_36; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_37; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_38; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_39; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_40; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_41; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_42; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_43; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_44; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_45; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_46; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_47; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_48; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_49; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_50; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_51; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_52; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_53; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_54; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_55; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_56; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_57; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_58; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_59; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_60; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_61; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_62; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_63; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_64; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_65; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_66; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_67; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_68; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_69; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_70; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_71; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_72; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_73; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_74; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_75; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_76; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_77; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_78; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_79; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_80; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_81; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_82; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_83; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_84; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_85; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_86; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_87; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_88; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_89; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_90; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_91; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_92; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_93; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_94; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_95; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_96; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_97; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_98; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_99; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_100; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_101; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_102; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_103; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_104; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_105; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_106; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_107; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_108; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_109; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_110; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_111; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_112; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_113; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_114; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_115; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_116; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_117; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_118; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_119; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_120; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_121; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_122; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_123; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_124; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_125; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_126; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_127; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_128; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_129; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_130; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_131; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_132; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_133; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_134; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_135; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_136; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_137; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_138; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_139; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_140; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_141; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_142; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_143; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_144; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_145; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_146; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_147; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_148; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_149; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_150; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_151; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_152; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_153; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_154; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_155; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_156; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_157; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_158; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_159; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_160; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_161; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_162; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_163; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_164; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_165; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_166; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_167; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_168; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_169; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_170; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_171; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_172; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_173; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_174; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_175; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_176; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_177; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_178; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_179; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_180; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_181; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_182; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_183; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_184; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_185; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_186; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_187; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_188; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_189; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_190; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_191; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_192; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_193; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_194; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_195; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_196; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_197; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_198; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_199; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_200; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_201; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_202; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_203; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_204; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_205; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_206; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_207; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_208; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_209; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_210; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_211; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_212; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_213; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_214; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_215; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_216; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_217; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_218; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_219; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_220; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_221; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_222; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_223; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_224; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_225; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_226; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_227; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_228; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_229; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_230; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_231; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_232; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_233; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_234; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_235; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_236; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_237; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_238; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_239; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_240; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_241; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_242; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_243; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_244; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_245; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_246; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_247; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_248; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_249; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_250; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_251; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_252; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_253; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_254; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_255; // @[matcher_pisa.scala 335:23]
  wire [3:0] pipe3_io_pipe_phv_in_next_processor_id; // @[matcher_pisa.scala 335:23]
  wire  pipe3_io_pipe_phv_in_next_config_id; // @[matcher_pisa.scala 335:23]
  wire  pipe3_io_pipe_phv_in_is_valid_processor; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_0; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_1; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_2; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_3; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_4; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_5; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_6; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_7; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_8; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_9; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_10; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_11; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_12; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_13; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_14; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_15; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_16; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_17; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_18; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_19; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_20; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_21; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_22; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_23; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_24; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_25; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_26; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_27; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_28; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_29; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_30; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_31; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_32; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_33; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_34; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_35; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_36; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_37; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_38; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_39; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_40; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_41; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_42; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_43; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_44; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_45; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_46; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_47; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_48; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_49; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_50; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_51; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_52; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_53; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_54; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_55; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_56; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_57; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_58; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_59; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_60; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_61; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_62; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_63; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_64; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_65; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_66; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_67; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_68; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_69; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_70; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_71; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_72; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_73; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_74; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_75; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_76; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_77; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_78; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_79; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_80; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_81; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_82; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_83; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_84; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_85; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_86; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_87; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_88; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_89; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_90; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_91; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_92; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_93; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_94; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_95; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_96; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_97; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_98; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_99; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_100; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_101; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_102; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_103; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_104; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_105; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_106; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_107; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_108; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_109; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_110; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_111; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_112; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_113; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_114; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_115; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_116; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_117; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_118; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_119; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_120; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_121; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_122; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_123; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_124; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_125; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_126; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_127; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_128; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_129; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_130; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_131; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_132; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_133; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_134; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_135; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_136; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_137; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_138; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_139; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_140; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_141; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_142; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_143; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_144; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_145; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_146; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_147; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_148; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_149; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_150; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_151; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_152; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_153; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_154; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_155; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_156; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_157; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_158; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_159; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_160; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_161; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_162; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_163; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_164; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_165; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_166; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_167; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_168; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_169; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_170; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_171; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_172; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_173; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_174; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_175; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_176; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_177; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_178; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_179; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_180; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_181; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_182; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_183; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_184; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_185; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_186; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_187; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_188; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_189; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_190; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_191; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_192; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_193; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_194; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_195; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_196; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_197; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_198; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_199; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_200; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_201; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_202; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_203; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_204; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_205; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_206; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_207; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_208; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_209; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_210; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_211; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_212; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_213; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_214; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_215; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_216; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_217; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_218; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_219; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_220; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_221; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_222; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_223; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_224; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_225; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_226; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_227; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_228; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_229; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_230; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_231; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_232; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_233; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_234; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_235; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_236; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_237; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_238; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_239; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_240; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_241; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_242; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_243; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_244; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_245; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_246; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_247; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_248; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_249; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_250; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_251; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_252; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_253; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_254; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_255; // @[matcher_pisa.scala 335:23]
  wire [3:0] pipe3_io_pipe_phv_out_next_processor_id; // @[matcher_pisa.scala 335:23]
  wire  pipe3_io_pipe_phv_out_next_config_id; // @[matcher_pisa.scala 335:23]
  wire  pipe3_io_pipe_phv_out_is_valid_processor; // @[matcher_pisa.scala 335:23]
  wire [4:0] pipe3_io_table_config_0_table_depth; // @[matcher_pisa.scala 335:23]
  wire [4:0] pipe3_io_table_config_0_table_width; // @[matcher_pisa.scala 335:23]
  wire [4:0] pipe3_io_table_config_1_table_depth; // @[matcher_pisa.scala 335:23]
  wire [4:0] pipe3_io_table_config_1_table_width; // @[matcher_pisa.scala 335:23]
  wire [191:0] pipe3_io_key_in; // @[matcher_pisa.scala 335:23]
  wire [191:0] pipe3_io_key_out; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_addr_in; // @[matcher_pisa.scala 335:23]
  wire [3:0] pipe3_io_cs_in; // @[matcher_pisa.scala 335:23]
  wire [255:0] pipe3_io_data_out; // @[matcher_pisa.scala 335:23]
  wire  pipe3_io_w_en; // @[matcher_pisa.scala 335:23]
  wire [3:0] pipe3_io_w_sram_id; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_w_addr; // @[matcher_pisa.scala 335:23]
  wire [63:0] pipe3_io_w_data; // @[matcher_pisa.scala 335:23]
  wire  pipe4_clock; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_0; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_1; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_2; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_3; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_4; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_5; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_6; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_7; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_8; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_9; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_10; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_11; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_12; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_13; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_14; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_15; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_16; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_17; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_18; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_19; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_20; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_21; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_22; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_23; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_24; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_25; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_26; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_27; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_28; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_29; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_30; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_31; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_32; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_33; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_34; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_35; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_36; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_37; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_38; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_39; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_40; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_41; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_42; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_43; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_44; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_45; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_46; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_47; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_48; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_49; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_50; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_51; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_52; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_53; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_54; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_55; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_56; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_57; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_58; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_59; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_60; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_61; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_62; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_63; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_64; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_65; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_66; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_67; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_68; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_69; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_70; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_71; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_72; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_73; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_74; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_75; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_76; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_77; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_78; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_79; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_80; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_81; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_82; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_83; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_84; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_85; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_86; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_87; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_88; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_89; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_90; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_91; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_92; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_93; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_94; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_95; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_96; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_97; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_98; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_99; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_100; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_101; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_102; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_103; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_104; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_105; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_106; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_107; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_108; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_109; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_110; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_111; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_112; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_113; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_114; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_115; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_116; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_117; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_118; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_119; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_120; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_121; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_122; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_123; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_124; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_125; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_126; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_127; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_128; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_129; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_130; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_131; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_132; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_133; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_134; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_135; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_136; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_137; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_138; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_139; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_140; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_141; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_142; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_143; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_144; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_145; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_146; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_147; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_148; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_149; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_150; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_151; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_152; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_153; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_154; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_155; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_156; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_157; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_158; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_159; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_160; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_161; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_162; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_163; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_164; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_165; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_166; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_167; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_168; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_169; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_170; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_171; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_172; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_173; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_174; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_175; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_176; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_177; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_178; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_179; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_180; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_181; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_182; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_183; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_184; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_185; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_186; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_187; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_188; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_189; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_190; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_191; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_192; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_193; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_194; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_195; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_196; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_197; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_198; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_199; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_200; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_201; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_202; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_203; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_204; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_205; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_206; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_207; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_208; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_209; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_210; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_211; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_212; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_213; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_214; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_215; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_216; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_217; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_218; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_219; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_220; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_221; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_222; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_223; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_224; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_225; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_226; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_227; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_228; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_229; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_230; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_231; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_232; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_233; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_234; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_235; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_236; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_237; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_238; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_239; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_240; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_241; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_242; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_243; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_244; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_245; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_246; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_247; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_248; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_249; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_250; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_251; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_252; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_253; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_254; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_255; // @[matcher_pisa.scala 336:23]
  wire [3:0] pipe4_io_pipe_phv_in_next_processor_id; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_pipe_phv_in_next_config_id; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_pipe_phv_in_is_valid_processor; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_0; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_1; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_2; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_3; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_4; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_5; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_6; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_7; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_8; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_9; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_10; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_11; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_12; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_13; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_14; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_15; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_16; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_17; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_18; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_19; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_20; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_21; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_22; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_23; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_24; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_25; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_26; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_27; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_28; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_29; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_30; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_31; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_32; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_33; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_34; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_35; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_36; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_37; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_38; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_39; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_40; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_41; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_42; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_43; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_44; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_45; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_46; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_47; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_48; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_49; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_50; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_51; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_52; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_53; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_54; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_55; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_56; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_57; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_58; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_59; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_60; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_61; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_62; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_63; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_64; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_65; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_66; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_67; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_68; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_69; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_70; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_71; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_72; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_73; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_74; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_75; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_76; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_77; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_78; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_79; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_80; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_81; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_82; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_83; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_84; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_85; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_86; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_87; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_88; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_89; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_90; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_91; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_92; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_93; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_94; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_95; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_96; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_97; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_98; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_99; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_100; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_101; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_102; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_103; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_104; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_105; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_106; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_107; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_108; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_109; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_110; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_111; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_112; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_113; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_114; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_115; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_116; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_117; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_118; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_119; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_120; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_121; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_122; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_123; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_124; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_125; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_126; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_127; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_128; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_129; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_130; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_131; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_132; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_133; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_134; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_135; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_136; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_137; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_138; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_139; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_140; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_141; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_142; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_143; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_144; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_145; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_146; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_147; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_148; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_149; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_150; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_151; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_152; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_153; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_154; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_155; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_156; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_157; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_158; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_159; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_160; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_161; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_162; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_163; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_164; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_165; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_166; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_167; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_168; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_169; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_170; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_171; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_172; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_173; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_174; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_175; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_176; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_177; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_178; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_179; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_180; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_181; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_182; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_183; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_184; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_185; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_186; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_187; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_188; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_189; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_190; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_191; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_192; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_193; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_194; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_195; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_196; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_197; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_198; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_199; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_200; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_201; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_202; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_203; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_204; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_205; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_206; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_207; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_208; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_209; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_210; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_211; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_212; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_213; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_214; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_215; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_216; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_217; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_218; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_219; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_220; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_221; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_222; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_223; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_224; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_225; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_226; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_227; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_228; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_229; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_230; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_231; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_232; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_233; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_234; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_235; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_236; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_237; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_238; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_239; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_240; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_241; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_242; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_243; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_244; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_245; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_246; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_247; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_248; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_249; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_250; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_251; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_252; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_253; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_254; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_255; // @[matcher_pisa.scala 336:23]
  wire [3:0] pipe4_io_pipe_phv_out_next_processor_id; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_pipe_phv_out_next_config_id; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_pipe_phv_out_is_valid_processor; // @[matcher_pisa.scala 336:23]
  wire [1:0] pipe4_io_key_config_0_field_config_0; // @[matcher_pisa.scala 336:23]
  wire [1:0] pipe4_io_key_config_0_field_config_1; // @[matcher_pisa.scala 336:23]
  wire [1:0] pipe4_io_key_config_0_field_config_2; // @[matcher_pisa.scala 336:23]
  wire [1:0] pipe4_io_key_config_0_field_config_3; // @[matcher_pisa.scala 336:23]
  wire [1:0] pipe4_io_key_config_0_field_config_4; // @[matcher_pisa.scala 336:23]
  wire [1:0] pipe4_io_key_config_0_field_config_5; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_0_field_mask_0_0; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_0_field_mask_0_1; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_0_field_mask_0_2; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_0_field_mask_0_3; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_0_field_mask_1_0; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_0_field_mask_1_1; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_0_field_mask_1_2; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_0_field_mask_1_3; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_0_field_mask_2_0; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_0_field_mask_2_1; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_0_field_mask_2_2; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_0_field_mask_2_3; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_0_field_mask_3_0; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_0_field_mask_3_1; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_0_field_mask_3_2; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_0_field_mask_3_3; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_0_field_mask_4_0; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_0_field_mask_4_1; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_0_field_mask_4_2; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_0_field_mask_4_3; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_0_field_mask_5_0; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_0_field_mask_5_1; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_0_field_mask_5_2; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_0_field_mask_5_3; // @[matcher_pisa.scala 336:23]
  wire [1:0] pipe4_io_key_config_1_field_config_0; // @[matcher_pisa.scala 336:23]
  wire [1:0] pipe4_io_key_config_1_field_config_1; // @[matcher_pisa.scala 336:23]
  wire [1:0] pipe4_io_key_config_1_field_config_2; // @[matcher_pisa.scala 336:23]
  wire [1:0] pipe4_io_key_config_1_field_config_3; // @[matcher_pisa.scala 336:23]
  wire [1:0] pipe4_io_key_config_1_field_config_4; // @[matcher_pisa.scala 336:23]
  wire [1:0] pipe4_io_key_config_1_field_config_5; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_1_field_mask_0_0; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_1_field_mask_0_1; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_1_field_mask_0_2; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_1_field_mask_0_3; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_1_field_mask_1_0; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_1_field_mask_1_1; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_1_field_mask_1_2; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_1_field_mask_1_3; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_1_field_mask_2_0; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_1_field_mask_2_1; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_1_field_mask_2_2; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_1_field_mask_2_3; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_1_field_mask_3_0; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_1_field_mask_3_1; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_1_field_mask_3_2; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_1_field_mask_3_3; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_1_field_mask_4_0; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_1_field_mask_4_1; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_1_field_mask_4_2; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_1_field_mask_4_3; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_1_field_mask_5_0; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_1_field_mask_5_1; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_1_field_mask_5_2; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_1_field_mask_5_3; // @[matcher_pisa.scala 336:23]
  wire [191:0] pipe4_io_key_in; // @[matcher_pisa.scala 336:23]
  wire [255:0] pipe4_io_data_in; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_hit; // @[matcher_pisa.scala 336:23]
  wire [63:0] pipe4_io_match_value; // @[matcher_pisa.scala 336:23]
  reg [1:0] key_config_0_field_config_0; // @[matcher_pisa.scala 70:25]
  reg [1:0] key_config_0_field_config_1; // @[matcher_pisa.scala 70:25]
  reg [1:0] key_config_0_field_config_2; // @[matcher_pisa.scala 70:25]
  reg [1:0] key_config_0_field_config_3; // @[matcher_pisa.scala 70:25]
  reg [1:0] key_config_0_field_config_4; // @[matcher_pisa.scala 70:25]
  reg [1:0] key_config_0_field_config_5; // @[matcher_pisa.scala 70:25]
  reg  key_config_0_field_mask_0_0; // @[matcher_pisa.scala 70:25]
  reg  key_config_0_field_mask_0_1; // @[matcher_pisa.scala 70:25]
  reg  key_config_0_field_mask_0_2; // @[matcher_pisa.scala 70:25]
  reg  key_config_0_field_mask_0_3; // @[matcher_pisa.scala 70:25]
  reg  key_config_0_field_mask_1_0; // @[matcher_pisa.scala 70:25]
  reg  key_config_0_field_mask_1_1; // @[matcher_pisa.scala 70:25]
  reg  key_config_0_field_mask_1_2; // @[matcher_pisa.scala 70:25]
  reg  key_config_0_field_mask_1_3; // @[matcher_pisa.scala 70:25]
  reg  key_config_0_field_mask_2_0; // @[matcher_pisa.scala 70:25]
  reg  key_config_0_field_mask_2_1; // @[matcher_pisa.scala 70:25]
  reg  key_config_0_field_mask_2_2; // @[matcher_pisa.scala 70:25]
  reg  key_config_0_field_mask_2_3; // @[matcher_pisa.scala 70:25]
  reg  key_config_0_field_mask_3_0; // @[matcher_pisa.scala 70:25]
  reg  key_config_0_field_mask_3_1; // @[matcher_pisa.scala 70:25]
  reg  key_config_0_field_mask_3_2; // @[matcher_pisa.scala 70:25]
  reg  key_config_0_field_mask_3_3; // @[matcher_pisa.scala 70:25]
  reg  key_config_0_field_mask_4_0; // @[matcher_pisa.scala 70:25]
  reg  key_config_0_field_mask_4_1; // @[matcher_pisa.scala 70:25]
  reg  key_config_0_field_mask_4_2; // @[matcher_pisa.scala 70:25]
  reg  key_config_0_field_mask_4_3; // @[matcher_pisa.scala 70:25]
  reg  key_config_0_field_mask_5_0; // @[matcher_pisa.scala 70:25]
  reg  key_config_0_field_mask_5_1; // @[matcher_pisa.scala 70:25]
  reg  key_config_0_field_mask_5_2; // @[matcher_pisa.scala 70:25]
  reg  key_config_0_field_mask_5_3; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_0_field_id_0_0; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_0_field_id_0_1; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_0_field_id_0_2; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_0_field_id_0_3; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_0_field_id_1_0; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_0_field_id_1_1; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_0_field_id_1_2; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_0_field_id_1_3; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_0_field_id_2_0; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_0_field_id_2_1; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_0_field_id_2_2; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_0_field_id_2_3; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_0_field_id_3_0; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_0_field_id_3_1; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_0_field_id_3_2; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_0_field_id_3_3; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_0_field_id_4_0; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_0_field_id_4_1; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_0_field_id_4_2; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_0_field_id_4_3; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_0_field_id_5_0; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_0_field_id_5_1; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_0_field_id_5_2; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_0_field_id_5_3; // @[matcher_pisa.scala 70:25]
  reg [1:0] key_config_1_field_config_0; // @[matcher_pisa.scala 70:25]
  reg [1:0] key_config_1_field_config_1; // @[matcher_pisa.scala 70:25]
  reg [1:0] key_config_1_field_config_2; // @[matcher_pisa.scala 70:25]
  reg [1:0] key_config_1_field_config_3; // @[matcher_pisa.scala 70:25]
  reg [1:0] key_config_1_field_config_4; // @[matcher_pisa.scala 70:25]
  reg [1:0] key_config_1_field_config_5; // @[matcher_pisa.scala 70:25]
  reg  key_config_1_field_mask_0_0; // @[matcher_pisa.scala 70:25]
  reg  key_config_1_field_mask_0_1; // @[matcher_pisa.scala 70:25]
  reg  key_config_1_field_mask_0_2; // @[matcher_pisa.scala 70:25]
  reg  key_config_1_field_mask_0_3; // @[matcher_pisa.scala 70:25]
  reg  key_config_1_field_mask_1_0; // @[matcher_pisa.scala 70:25]
  reg  key_config_1_field_mask_1_1; // @[matcher_pisa.scala 70:25]
  reg  key_config_1_field_mask_1_2; // @[matcher_pisa.scala 70:25]
  reg  key_config_1_field_mask_1_3; // @[matcher_pisa.scala 70:25]
  reg  key_config_1_field_mask_2_0; // @[matcher_pisa.scala 70:25]
  reg  key_config_1_field_mask_2_1; // @[matcher_pisa.scala 70:25]
  reg  key_config_1_field_mask_2_2; // @[matcher_pisa.scala 70:25]
  reg  key_config_1_field_mask_2_3; // @[matcher_pisa.scala 70:25]
  reg  key_config_1_field_mask_3_0; // @[matcher_pisa.scala 70:25]
  reg  key_config_1_field_mask_3_1; // @[matcher_pisa.scala 70:25]
  reg  key_config_1_field_mask_3_2; // @[matcher_pisa.scala 70:25]
  reg  key_config_1_field_mask_3_3; // @[matcher_pisa.scala 70:25]
  reg  key_config_1_field_mask_4_0; // @[matcher_pisa.scala 70:25]
  reg  key_config_1_field_mask_4_1; // @[matcher_pisa.scala 70:25]
  reg  key_config_1_field_mask_4_2; // @[matcher_pisa.scala 70:25]
  reg  key_config_1_field_mask_4_3; // @[matcher_pisa.scala 70:25]
  reg  key_config_1_field_mask_5_0; // @[matcher_pisa.scala 70:25]
  reg  key_config_1_field_mask_5_1; // @[matcher_pisa.scala 70:25]
  reg  key_config_1_field_mask_5_2; // @[matcher_pisa.scala 70:25]
  reg  key_config_1_field_mask_5_3; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_1_field_id_0_0; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_1_field_id_0_1; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_1_field_id_0_2; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_1_field_id_0_3; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_1_field_id_1_0; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_1_field_id_1_1; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_1_field_id_1_2; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_1_field_id_1_3; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_1_field_id_2_0; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_1_field_id_2_1; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_1_field_id_2_2; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_1_field_id_2_3; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_1_field_id_3_0; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_1_field_id_3_1; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_1_field_id_3_2; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_1_field_id_3_3; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_1_field_id_4_0; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_1_field_id_4_1; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_1_field_id_4_2; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_1_field_id_4_3; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_1_field_id_5_0; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_1_field_id_5_1; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_1_field_id_5_2; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_1_field_id_5_3; // @[matcher_pisa.scala 70:25]
  reg [4:0] table_config_0_table_depth; // @[matcher_pisa.scala 71:27]
  reg [4:0] table_config_0_table_width; // @[matcher_pisa.scala 71:27]
  reg [4:0] table_config_1_table_depth; // @[matcher_pisa.scala 71:27]
  reg [4:0] table_config_1_table_width; // @[matcher_pisa.scala 71:27]
  wire  _GEN_338 = ~io_mod_config_id; // @[matcher_pisa.scala 74:83 matcher_pisa.scala 74:83 matcher_pisa.scala 70:25]
  wire  _GEN_339 = 3'h0 == io_mod_key_mod_group_index; // @[matcher_pisa.scala 74:83 matcher_pisa.scala 74:83 matcher_pisa.scala 70:25]
  wire  _GEN_341 = 3'h1 == io_mod_key_mod_group_index; // @[matcher_pisa.scala 74:83 matcher_pisa.scala 74:83 matcher_pisa.scala 70:25]
  wire  _GEN_343 = 3'h2 == io_mod_key_mod_group_index; // @[matcher_pisa.scala 74:83 matcher_pisa.scala 74:83 matcher_pisa.scala 70:25]
  wire  _GEN_345 = 3'h3 == io_mod_key_mod_group_index; // @[matcher_pisa.scala 74:83 matcher_pisa.scala 74:83 matcher_pisa.scala 70:25]
  wire  _GEN_347 = 3'h4 == io_mod_key_mod_group_index; // @[matcher_pisa.scala 74:83 matcher_pisa.scala 74:83 matcher_pisa.scala 70:25]
  wire  _GEN_349 = 3'h5 == io_mod_key_mod_group_index; // @[matcher_pisa.scala 74:83 matcher_pisa.scala 74:83 matcher_pisa.scala 70:25]
  MatchGetKeyPISA pipe1 ( // @[matcher_pisa.scala 333:23]
    .clock(pipe1_clock),
    .io_pipe_phv_in_data_0(pipe1_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe1_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe1_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe1_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe1_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe1_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe1_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe1_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe1_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe1_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe1_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe1_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe1_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe1_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe1_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe1_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe1_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe1_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe1_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe1_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe1_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe1_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe1_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe1_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe1_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe1_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe1_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe1_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe1_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe1_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe1_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe1_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe1_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe1_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe1_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe1_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe1_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe1_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe1_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe1_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe1_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe1_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe1_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe1_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe1_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe1_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe1_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe1_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe1_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe1_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe1_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe1_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe1_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe1_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe1_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe1_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe1_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe1_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe1_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe1_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe1_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe1_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe1_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe1_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe1_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe1_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe1_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe1_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe1_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe1_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe1_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe1_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe1_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe1_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe1_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe1_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe1_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe1_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe1_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe1_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe1_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe1_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe1_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe1_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe1_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe1_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe1_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe1_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe1_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe1_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe1_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe1_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe1_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe1_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe1_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe1_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe1_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe1_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe1_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe1_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe1_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe1_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe1_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe1_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe1_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe1_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe1_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe1_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe1_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe1_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe1_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe1_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe1_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe1_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe1_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe1_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe1_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe1_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe1_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe1_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe1_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe1_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe1_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe1_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe1_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe1_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe1_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe1_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe1_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe1_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe1_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe1_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe1_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe1_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe1_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe1_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe1_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe1_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe1_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe1_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe1_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe1_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe1_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe1_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe1_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe1_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe1_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe1_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe1_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe1_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe1_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe1_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe1_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe1_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe1_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe1_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe1_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe1_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe1_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe1_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(pipe1_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(pipe1_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(pipe1_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(pipe1_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(pipe1_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(pipe1_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(pipe1_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(pipe1_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(pipe1_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(pipe1_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(pipe1_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(pipe1_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(pipe1_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(pipe1_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(pipe1_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(pipe1_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(pipe1_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(pipe1_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(pipe1_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(pipe1_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(pipe1_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(pipe1_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(pipe1_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(pipe1_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(pipe1_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(pipe1_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(pipe1_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(pipe1_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(pipe1_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(pipe1_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(pipe1_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(pipe1_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(pipe1_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(pipe1_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(pipe1_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(pipe1_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(pipe1_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(pipe1_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(pipe1_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(pipe1_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(pipe1_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(pipe1_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(pipe1_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(pipe1_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(pipe1_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(pipe1_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(pipe1_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(pipe1_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(pipe1_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(pipe1_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(pipe1_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(pipe1_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(pipe1_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(pipe1_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(pipe1_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(pipe1_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(pipe1_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(pipe1_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(pipe1_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(pipe1_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(pipe1_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(pipe1_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(pipe1_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(pipe1_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(pipe1_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(pipe1_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(pipe1_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(pipe1_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(pipe1_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(pipe1_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(pipe1_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(pipe1_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(pipe1_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(pipe1_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(pipe1_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(pipe1_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(pipe1_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(pipe1_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(pipe1_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(pipe1_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(pipe1_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(pipe1_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(pipe1_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(pipe1_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(pipe1_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(pipe1_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(pipe1_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(pipe1_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(pipe1_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(pipe1_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(pipe1_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(pipe1_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(pipe1_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(pipe1_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(pipe1_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(pipe1_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_next_processor_id(pipe1_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe1_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe1_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe1_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe1_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe1_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe1_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe1_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe1_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe1_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe1_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe1_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe1_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe1_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe1_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe1_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe1_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe1_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe1_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe1_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe1_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe1_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe1_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe1_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe1_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe1_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe1_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe1_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe1_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe1_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe1_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe1_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe1_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe1_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe1_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe1_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe1_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe1_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe1_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe1_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe1_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe1_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe1_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe1_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe1_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe1_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe1_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe1_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe1_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe1_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe1_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe1_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe1_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe1_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe1_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe1_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe1_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe1_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe1_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe1_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe1_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe1_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe1_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe1_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe1_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe1_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe1_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe1_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe1_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe1_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe1_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe1_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe1_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe1_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe1_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe1_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe1_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe1_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe1_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe1_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe1_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe1_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe1_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe1_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe1_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe1_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe1_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe1_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe1_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe1_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe1_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe1_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe1_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe1_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe1_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe1_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe1_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe1_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe1_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe1_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe1_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe1_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe1_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe1_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe1_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe1_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe1_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe1_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe1_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe1_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe1_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe1_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe1_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe1_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe1_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe1_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe1_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe1_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe1_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe1_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe1_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe1_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe1_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe1_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe1_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe1_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe1_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe1_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe1_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe1_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe1_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe1_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe1_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe1_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe1_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe1_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe1_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe1_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe1_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe1_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe1_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe1_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe1_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe1_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe1_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe1_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe1_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe1_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe1_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe1_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe1_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe1_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe1_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe1_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe1_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe1_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe1_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe1_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe1_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe1_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe1_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe1_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe1_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(pipe1_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(pipe1_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(pipe1_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(pipe1_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(pipe1_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(pipe1_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(pipe1_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(pipe1_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(pipe1_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(pipe1_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(pipe1_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(pipe1_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(pipe1_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(pipe1_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(pipe1_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(pipe1_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(pipe1_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(pipe1_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(pipe1_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(pipe1_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(pipe1_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(pipe1_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(pipe1_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(pipe1_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(pipe1_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(pipe1_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(pipe1_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(pipe1_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(pipe1_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(pipe1_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(pipe1_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(pipe1_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(pipe1_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(pipe1_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(pipe1_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(pipe1_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(pipe1_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(pipe1_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(pipe1_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(pipe1_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(pipe1_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(pipe1_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(pipe1_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(pipe1_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(pipe1_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(pipe1_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(pipe1_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(pipe1_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(pipe1_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(pipe1_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(pipe1_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(pipe1_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(pipe1_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(pipe1_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(pipe1_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(pipe1_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(pipe1_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(pipe1_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(pipe1_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(pipe1_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(pipe1_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(pipe1_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(pipe1_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(pipe1_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(pipe1_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(pipe1_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(pipe1_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(pipe1_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(pipe1_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(pipe1_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(pipe1_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(pipe1_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(pipe1_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(pipe1_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(pipe1_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(pipe1_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(pipe1_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(pipe1_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(pipe1_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(pipe1_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(pipe1_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(pipe1_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(pipe1_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(pipe1_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(pipe1_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(pipe1_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(pipe1_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(pipe1_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(pipe1_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(pipe1_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(pipe1_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(pipe1_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(pipe1_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(pipe1_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(pipe1_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(pipe1_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_next_processor_id(pipe1_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe1_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe1_io_pipe_phv_out_is_valid_processor),
    .io_key_config_0_field_config_0(pipe1_io_key_config_0_field_config_0),
    .io_key_config_0_field_config_1(pipe1_io_key_config_0_field_config_1),
    .io_key_config_0_field_config_2(pipe1_io_key_config_0_field_config_2),
    .io_key_config_0_field_config_3(pipe1_io_key_config_0_field_config_3),
    .io_key_config_0_field_config_4(pipe1_io_key_config_0_field_config_4),
    .io_key_config_0_field_config_5(pipe1_io_key_config_0_field_config_5),
    .io_key_config_0_field_mask_0_0(pipe1_io_key_config_0_field_mask_0_0),
    .io_key_config_0_field_mask_0_1(pipe1_io_key_config_0_field_mask_0_1),
    .io_key_config_0_field_mask_0_2(pipe1_io_key_config_0_field_mask_0_2),
    .io_key_config_0_field_mask_0_3(pipe1_io_key_config_0_field_mask_0_3),
    .io_key_config_0_field_mask_1_0(pipe1_io_key_config_0_field_mask_1_0),
    .io_key_config_0_field_mask_1_1(pipe1_io_key_config_0_field_mask_1_1),
    .io_key_config_0_field_mask_1_2(pipe1_io_key_config_0_field_mask_1_2),
    .io_key_config_0_field_mask_1_3(pipe1_io_key_config_0_field_mask_1_3),
    .io_key_config_0_field_mask_2_0(pipe1_io_key_config_0_field_mask_2_0),
    .io_key_config_0_field_mask_2_1(pipe1_io_key_config_0_field_mask_2_1),
    .io_key_config_0_field_mask_2_2(pipe1_io_key_config_0_field_mask_2_2),
    .io_key_config_0_field_mask_2_3(pipe1_io_key_config_0_field_mask_2_3),
    .io_key_config_0_field_mask_3_0(pipe1_io_key_config_0_field_mask_3_0),
    .io_key_config_0_field_mask_3_1(pipe1_io_key_config_0_field_mask_3_1),
    .io_key_config_0_field_mask_3_2(pipe1_io_key_config_0_field_mask_3_2),
    .io_key_config_0_field_mask_3_3(pipe1_io_key_config_0_field_mask_3_3),
    .io_key_config_0_field_mask_4_0(pipe1_io_key_config_0_field_mask_4_0),
    .io_key_config_0_field_mask_4_1(pipe1_io_key_config_0_field_mask_4_1),
    .io_key_config_0_field_mask_4_2(pipe1_io_key_config_0_field_mask_4_2),
    .io_key_config_0_field_mask_4_3(pipe1_io_key_config_0_field_mask_4_3),
    .io_key_config_0_field_mask_5_0(pipe1_io_key_config_0_field_mask_5_0),
    .io_key_config_0_field_mask_5_1(pipe1_io_key_config_0_field_mask_5_1),
    .io_key_config_0_field_mask_5_2(pipe1_io_key_config_0_field_mask_5_2),
    .io_key_config_0_field_mask_5_3(pipe1_io_key_config_0_field_mask_5_3),
    .io_key_config_0_field_id_0_0(pipe1_io_key_config_0_field_id_0_0),
    .io_key_config_0_field_id_0_1(pipe1_io_key_config_0_field_id_0_1),
    .io_key_config_0_field_id_0_2(pipe1_io_key_config_0_field_id_0_2),
    .io_key_config_0_field_id_0_3(pipe1_io_key_config_0_field_id_0_3),
    .io_key_config_0_field_id_1_0(pipe1_io_key_config_0_field_id_1_0),
    .io_key_config_0_field_id_1_1(pipe1_io_key_config_0_field_id_1_1),
    .io_key_config_0_field_id_1_2(pipe1_io_key_config_0_field_id_1_2),
    .io_key_config_0_field_id_1_3(pipe1_io_key_config_0_field_id_1_3),
    .io_key_config_0_field_id_2_0(pipe1_io_key_config_0_field_id_2_0),
    .io_key_config_0_field_id_2_1(pipe1_io_key_config_0_field_id_2_1),
    .io_key_config_0_field_id_2_2(pipe1_io_key_config_0_field_id_2_2),
    .io_key_config_0_field_id_2_3(pipe1_io_key_config_0_field_id_2_3),
    .io_key_config_0_field_id_3_0(pipe1_io_key_config_0_field_id_3_0),
    .io_key_config_0_field_id_3_1(pipe1_io_key_config_0_field_id_3_1),
    .io_key_config_0_field_id_3_2(pipe1_io_key_config_0_field_id_3_2),
    .io_key_config_0_field_id_3_3(pipe1_io_key_config_0_field_id_3_3),
    .io_key_config_0_field_id_4_0(pipe1_io_key_config_0_field_id_4_0),
    .io_key_config_0_field_id_4_1(pipe1_io_key_config_0_field_id_4_1),
    .io_key_config_0_field_id_4_2(pipe1_io_key_config_0_field_id_4_2),
    .io_key_config_0_field_id_4_3(pipe1_io_key_config_0_field_id_4_3),
    .io_key_config_0_field_id_5_0(pipe1_io_key_config_0_field_id_5_0),
    .io_key_config_0_field_id_5_1(pipe1_io_key_config_0_field_id_5_1),
    .io_key_config_0_field_id_5_2(pipe1_io_key_config_0_field_id_5_2),
    .io_key_config_0_field_id_5_3(pipe1_io_key_config_0_field_id_5_3),
    .io_key_config_1_field_config_0(pipe1_io_key_config_1_field_config_0),
    .io_key_config_1_field_config_1(pipe1_io_key_config_1_field_config_1),
    .io_key_config_1_field_config_2(pipe1_io_key_config_1_field_config_2),
    .io_key_config_1_field_config_3(pipe1_io_key_config_1_field_config_3),
    .io_key_config_1_field_config_4(pipe1_io_key_config_1_field_config_4),
    .io_key_config_1_field_config_5(pipe1_io_key_config_1_field_config_5),
    .io_key_config_1_field_mask_0_0(pipe1_io_key_config_1_field_mask_0_0),
    .io_key_config_1_field_mask_0_1(pipe1_io_key_config_1_field_mask_0_1),
    .io_key_config_1_field_mask_0_2(pipe1_io_key_config_1_field_mask_0_2),
    .io_key_config_1_field_mask_0_3(pipe1_io_key_config_1_field_mask_0_3),
    .io_key_config_1_field_mask_1_0(pipe1_io_key_config_1_field_mask_1_0),
    .io_key_config_1_field_mask_1_1(pipe1_io_key_config_1_field_mask_1_1),
    .io_key_config_1_field_mask_1_2(pipe1_io_key_config_1_field_mask_1_2),
    .io_key_config_1_field_mask_1_3(pipe1_io_key_config_1_field_mask_1_3),
    .io_key_config_1_field_mask_2_0(pipe1_io_key_config_1_field_mask_2_0),
    .io_key_config_1_field_mask_2_1(pipe1_io_key_config_1_field_mask_2_1),
    .io_key_config_1_field_mask_2_2(pipe1_io_key_config_1_field_mask_2_2),
    .io_key_config_1_field_mask_2_3(pipe1_io_key_config_1_field_mask_2_3),
    .io_key_config_1_field_mask_3_0(pipe1_io_key_config_1_field_mask_3_0),
    .io_key_config_1_field_mask_3_1(pipe1_io_key_config_1_field_mask_3_1),
    .io_key_config_1_field_mask_3_2(pipe1_io_key_config_1_field_mask_3_2),
    .io_key_config_1_field_mask_3_3(pipe1_io_key_config_1_field_mask_3_3),
    .io_key_config_1_field_mask_4_0(pipe1_io_key_config_1_field_mask_4_0),
    .io_key_config_1_field_mask_4_1(pipe1_io_key_config_1_field_mask_4_1),
    .io_key_config_1_field_mask_4_2(pipe1_io_key_config_1_field_mask_4_2),
    .io_key_config_1_field_mask_4_3(pipe1_io_key_config_1_field_mask_4_3),
    .io_key_config_1_field_mask_5_0(pipe1_io_key_config_1_field_mask_5_0),
    .io_key_config_1_field_mask_5_1(pipe1_io_key_config_1_field_mask_5_1),
    .io_key_config_1_field_mask_5_2(pipe1_io_key_config_1_field_mask_5_2),
    .io_key_config_1_field_mask_5_3(pipe1_io_key_config_1_field_mask_5_3),
    .io_key_config_1_field_id_0_0(pipe1_io_key_config_1_field_id_0_0),
    .io_key_config_1_field_id_0_1(pipe1_io_key_config_1_field_id_0_1),
    .io_key_config_1_field_id_0_2(pipe1_io_key_config_1_field_id_0_2),
    .io_key_config_1_field_id_0_3(pipe1_io_key_config_1_field_id_0_3),
    .io_key_config_1_field_id_1_0(pipe1_io_key_config_1_field_id_1_0),
    .io_key_config_1_field_id_1_1(pipe1_io_key_config_1_field_id_1_1),
    .io_key_config_1_field_id_1_2(pipe1_io_key_config_1_field_id_1_2),
    .io_key_config_1_field_id_1_3(pipe1_io_key_config_1_field_id_1_3),
    .io_key_config_1_field_id_2_0(pipe1_io_key_config_1_field_id_2_0),
    .io_key_config_1_field_id_2_1(pipe1_io_key_config_1_field_id_2_1),
    .io_key_config_1_field_id_2_2(pipe1_io_key_config_1_field_id_2_2),
    .io_key_config_1_field_id_2_3(pipe1_io_key_config_1_field_id_2_3),
    .io_key_config_1_field_id_3_0(pipe1_io_key_config_1_field_id_3_0),
    .io_key_config_1_field_id_3_1(pipe1_io_key_config_1_field_id_3_1),
    .io_key_config_1_field_id_3_2(pipe1_io_key_config_1_field_id_3_2),
    .io_key_config_1_field_id_3_3(pipe1_io_key_config_1_field_id_3_3),
    .io_key_config_1_field_id_4_0(pipe1_io_key_config_1_field_id_4_0),
    .io_key_config_1_field_id_4_1(pipe1_io_key_config_1_field_id_4_1),
    .io_key_config_1_field_id_4_2(pipe1_io_key_config_1_field_id_4_2),
    .io_key_config_1_field_id_4_3(pipe1_io_key_config_1_field_id_4_3),
    .io_key_config_1_field_id_5_0(pipe1_io_key_config_1_field_id_5_0),
    .io_key_config_1_field_id_5_1(pipe1_io_key_config_1_field_id_5_1),
    .io_key_config_1_field_id_5_2(pipe1_io_key_config_1_field_id_5_2),
    .io_key_config_1_field_id_5_3(pipe1_io_key_config_1_field_id_5_3),
    .io_match_key(pipe1_io_match_key)
  );
  Hash pipe2 ( // @[matcher_pisa.scala 334:23]
    .clock(pipe2_clock),
    .io_pipe_phv_in_data_0(pipe2_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe2_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe2_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe2_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe2_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe2_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe2_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe2_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe2_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe2_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe2_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe2_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe2_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe2_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe2_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe2_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe2_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe2_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe2_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe2_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe2_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe2_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe2_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe2_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe2_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe2_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe2_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe2_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe2_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe2_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe2_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe2_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe2_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe2_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe2_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe2_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe2_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe2_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe2_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe2_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe2_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe2_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe2_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe2_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe2_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe2_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe2_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe2_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe2_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe2_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe2_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe2_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe2_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe2_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe2_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe2_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe2_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe2_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe2_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe2_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe2_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe2_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe2_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe2_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe2_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe2_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe2_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe2_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe2_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe2_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe2_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe2_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe2_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe2_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe2_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe2_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe2_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe2_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe2_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe2_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe2_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe2_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe2_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe2_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe2_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe2_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe2_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe2_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe2_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe2_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe2_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe2_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe2_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe2_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe2_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe2_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe2_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe2_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe2_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe2_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe2_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe2_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe2_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe2_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe2_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe2_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe2_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe2_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe2_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe2_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe2_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe2_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe2_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe2_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe2_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe2_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe2_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe2_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe2_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe2_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe2_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe2_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe2_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe2_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe2_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe2_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe2_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe2_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe2_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe2_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe2_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe2_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe2_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe2_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe2_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe2_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe2_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe2_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe2_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe2_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe2_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe2_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe2_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe2_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe2_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe2_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe2_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe2_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe2_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe2_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe2_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe2_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe2_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe2_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe2_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe2_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe2_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe2_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe2_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe2_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(pipe2_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(pipe2_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(pipe2_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(pipe2_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(pipe2_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(pipe2_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(pipe2_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(pipe2_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(pipe2_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(pipe2_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(pipe2_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(pipe2_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(pipe2_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(pipe2_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(pipe2_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(pipe2_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(pipe2_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(pipe2_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(pipe2_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(pipe2_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(pipe2_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(pipe2_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(pipe2_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(pipe2_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(pipe2_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(pipe2_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(pipe2_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(pipe2_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(pipe2_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(pipe2_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(pipe2_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(pipe2_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(pipe2_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(pipe2_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(pipe2_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(pipe2_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(pipe2_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(pipe2_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(pipe2_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(pipe2_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(pipe2_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(pipe2_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(pipe2_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(pipe2_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(pipe2_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(pipe2_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(pipe2_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(pipe2_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(pipe2_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(pipe2_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(pipe2_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(pipe2_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(pipe2_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(pipe2_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(pipe2_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(pipe2_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(pipe2_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(pipe2_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(pipe2_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(pipe2_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(pipe2_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(pipe2_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(pipe2_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(pipe2_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(pipe2_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(pipe2_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(pipe2_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(pipe2_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(pipe2_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(pipe2_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(pipe2_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(pipe2_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(pipe2_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(pipe2_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(pipe2_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(pipe2_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(pipe2_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(pipe2_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(pipe2_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(pipe2_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(pipe2_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(pipe2_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(pipe2_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(pipe2_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(pipe2_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(pipe2_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(pipe2_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(pipe2_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(pipe2_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(pipe2_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(pipe2_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(pipe2_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(pipe2_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(pipe2_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(pipe2_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(pipe2_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_next_processor_id(pipe2_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe2_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe2_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe2_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe2_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe2_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe2_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe2_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe2_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe2_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe2_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe2_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe2_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe2_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe2_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe2_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe2_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe2_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe2_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe2_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe2_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe2_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe2_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe2_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe2_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe2_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe2_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe2_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe2_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe2_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe2_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe2_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe2_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe2_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe2_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe2_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe2_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe2_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe2_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe2_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe2_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe2_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe2_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe2_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe2_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe2_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe2_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe2_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe2_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe2_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe2_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe2_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe2_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe2_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe2_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe2_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe2_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe2_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe2_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe2_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe2_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe2_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe2_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe2_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe2_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe2_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe2_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe2_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe2_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe2_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe2_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe2_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe2_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe2_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe2_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe2_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe2_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe2_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe2_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe2_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe2_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe2_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe2_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe2_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe2_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe2_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe2_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe2_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe2_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe2_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe2_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe2_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe2_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe2_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe2_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe2_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe2_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe2_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe2_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe2_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe2_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe2_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe2_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe2_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe2_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe2_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe2_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe2_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe2_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe2_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe2_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe2_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe2_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe2_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe2_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe2_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe2_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe2_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe2_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe2_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe2_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe2_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe2_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe2_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe2_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe2_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe2_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe2_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe2_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe2_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe2_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe2_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe2_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe2_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe2_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe2_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe2_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe2_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe2_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe2_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe2_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe2_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe2_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe2_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe2_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe2_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe2_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe2_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe2_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe2_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe2_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe2_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe2_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe2_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe2_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe2_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe2_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe2_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe2_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe2_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe2_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe2_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe2_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(pipe2_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(pipe2_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(pipe2_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(pipe2_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(pipe2_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(pipe2_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(pipe2_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(pipe2_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(pipe2_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(pipe2_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(pipe2_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(pipe2_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(pipe2_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(pipe2_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(pipe2_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(pipe2_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(pipe2_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(pipe2_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(pipe2_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(pipe2_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(pipe2_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(pipe2_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(pipe2_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(pipe2_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(pipe2_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(pipe2_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(pipe2_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(pipe2_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(pipe2_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(pipe2_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(pipe2_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(pipe2_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(pipe2_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(pipe2_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(pipe2_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(pipe2_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(pipe2_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(pipe2_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(pipe2_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(pipe2_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(pipe2_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(pipe2_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(pipe2_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(pipe2_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(pipe2_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(pipe2_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(pipe2_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(pipe2_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(pipe2_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(pipe2_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(pipe2_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(pipe2_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(pipe2_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(pipe2_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(pipe2_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(pipe2_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(pipe2_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(pipe2_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(pipe2_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(pipe2_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(pipe2_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(pipe2_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(pipe2_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(pipe2_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(pipe2_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(pipe2_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(pipe2_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(pipe2_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(pipe2_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(pipe2_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(pipe2_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(pipe2_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(pipe2_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(pipe2_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(pipe2_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(pipe2_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(pipe2_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(pipe2_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(pipe2_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(pipe2_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(pipe2_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(pipe2_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(pipe2_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(pipe2_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(pipe2_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(pipe2_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(pipe2_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(pipe2_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(pipe2_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(pipe2_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(pipe2_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(pipe2_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(pipe2_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(pipe2_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(pipe2_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(pipe2_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_next_processor_id(pipe2_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe2_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe2_io_pipe_phv_out_is_valid_processor),
    .io_mod_hash_depth_mod(pipe2_io_mod_hash_depth_mod),
    .io_mod_config_id(pipe2_io_mod_config_id),
    .io_mod_hash_depth(pipe2_io_mod_hash_depth),
    .io_key_in(pipe2_io_key_in),
    .io_key_out(pipe2_io_key_out),
    .io_hash_val(pipe2_io_hash_val),
    .io_hash_val_cs(pipe2_io_hash_val_cs)
  );
  MatchReadDataPISA pipe3 ( // @[matcher_pisa.scala 335:23]
    .clock(pipe3_clock),
    .io_pipe_phv_in_data_0(pipe3_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe3_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe3_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe3_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe3_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe3_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe3_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe3_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe3_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe3_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe3_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe3_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe3_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe3_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe3_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe3_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe3_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe3_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe3_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe3_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe3_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe3_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe3_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe3_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe3_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe3_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe3_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe3_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe3_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe3_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe3_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe3_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe3_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe3_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe3_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe3_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe3_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe3_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe3_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe3_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe3_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe3_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe3_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe3_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe3_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe3_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe3_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe3_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe3_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe3_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe3_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe3_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe3_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe3_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe3_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe3_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe3_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe3_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe3_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe3_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe3_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe3_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe3_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe3_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe3_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe3_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe3_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe3_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe3_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe3_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe3_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe3_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe3_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe3_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe3_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe3_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe3_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe3_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe3_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe3_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe3_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe3_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe3_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe3_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe3_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe3_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe3_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe3_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe3_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe3_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe3_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe3_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe3_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe3_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe3_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe3_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe3_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe3_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe3_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe3_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe3_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe3_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe3_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe3_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe3_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe3_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe3_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe3_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe3_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe3_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe3_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe3_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe3_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe3_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe3_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe3_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe3_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe3_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe3_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe3_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe3_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe3_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe3_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe3_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe3_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe3_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe3_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe3_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe3_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe3_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe3_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe3_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe3_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe3_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe3_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe3_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe3_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe3_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe3_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe3_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe3_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe3_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe3_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe3_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe3_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe3_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe3_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe3_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe3_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe3_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe3_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe3_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe3_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe3_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe3_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe3_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe3_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe3_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe3_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe3_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(pipe3_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(pipe3_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(pipe3_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(pipe3_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(pipe3_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(pipe3_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(pipe3_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(pipe3_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(pipe3_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(pipe3_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(pipe3_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(pipe3_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(pipe3_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(pipe3_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(pipe3_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(pipe3_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(pipe3_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(pipe3_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(pipe3_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(pipe3_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(pipe3_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(pipe3_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(pipe3_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(pipe3_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(pipe3_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(pipe3_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(pipe3_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(pipe3_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(pipe3_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(pipe3_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(pipe3_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(pipe3_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(pipe3_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(pipe3_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(pipe3_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(pipe3_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(pipe3_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(pipe3_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(pipe3_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(pipe3_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(pipe3_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(pipe3_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(pipe3_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(pipe3_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(pipe3_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(pipe3_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(pipe3_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(pipe3_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(pipe3_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(pipe3_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(pipe3_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(pipe3_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(pipe3_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(pipe3_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(pipe3_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(pipe3_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(pipe3_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(pipe3_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(pipe3_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(pipe3_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(pipe3_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(pipe3_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(pipe3_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(pipe3_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(pipe3_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(pipe3_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(pipe3_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(pipe3_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(pipe3_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(pipe3_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(pipe3_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(pipe3_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(pipe3_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(pipe3_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(pipe3_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(pipe3_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(pipe3_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(pipe3_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(pipe3_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(pipe3_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(pipe3_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(pipe3_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(pipe3_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(pipe3_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(pipe3_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(pipe3_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(pipe3_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(pipe3_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(pipe3_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(pipe3_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(pipe3_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(pipe3_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(pipe3_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(pipe3_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(pipe3_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(pipe3_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_next_processor_id(pipe3_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe3_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe3_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe3_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe3_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe3_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe3_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe3_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe3_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe3_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe3_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe3_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe3_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe3_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe3_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe3_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe3_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe3_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe3_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe3_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe3_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe3_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe3_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe3_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe3_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe3_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe3_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe3_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe3_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe3_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe3_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe3_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe3_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe3_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe3_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe3_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe3_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe3_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe3_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe3_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe3_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe3_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe3_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe3_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe3_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe3_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe3_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe3_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe3_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe3_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe3_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe3_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe3_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe3_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe3_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe3_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe3_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe3_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe3_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe3_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe3_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe3_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe3_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe3_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe3_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe3_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe3_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe3_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe3_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe3_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe3_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe3_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe3_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe3_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe3_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe3_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe3_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe3_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe3_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe3_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe3_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe3_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe3_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe3_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe3_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe3_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe3_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe3_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe3_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe3_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe3_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe3_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe3_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe3_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe3_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe3_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe3_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe3_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe3_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe3_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe3_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe3_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe3_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe3_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe3_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe3_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe3_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe3_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe3_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe3_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe3_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe3_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe3_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe3_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe3_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe3_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe3_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe3_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe3_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe3_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe3_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe3_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe3_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe3_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe3_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe3_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe3_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe3_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe3_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe3_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe3_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe3_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe3_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe3_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe3_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe3_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe3_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe3_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe3_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe3_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe3_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe3_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe3_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe3_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe3_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe3_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe3_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe3_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe3_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe3_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe3_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe3_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe3_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe3_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe3_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe3_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe3_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe3_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe3_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe3_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe3_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe3_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe3_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(pipe3_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(pipe3_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(pipe3_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(pipe3_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(pipe3_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(pipe3_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(pipe3_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(pipe3_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(pipe3_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(pipe3_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(pipe3_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(pipe3_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(pipe3_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(pipe3_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(pipe3_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(pipe3_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(pipe3_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(pipe3_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(pipe3_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(pipe3_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(pipe3_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(pipe3_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(pipe3_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(pipe3_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(pipe3_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(pipe3_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(pipe3_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(pipe3_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(pipe3_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(pipe3_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(pipe3_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(pipe3_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(pipe3_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(pipe3_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(pipe3_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(pipe3_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(pipe3_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(pipe3_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(pipe3_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(pipe3_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(pipe3_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(pipe3_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(pipe3_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(pipe3_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(pipe3_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(pipe3_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(pipe3_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(pipe3_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(pipe3_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(pipe3_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(pipe3_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(pipe3_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(pipe3_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(pipe3_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(pipe3_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(pipe3_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(pipe3_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(pipe3_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(pipe3_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(pipe3_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(pipe3_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(pipe3_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(pipe3_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(pipe3_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(pipe3_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(pipe3_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(pipe3_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(pipe3_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(pipe3_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(pipe3_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(pipe3_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(pipe3_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(pipe3_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(pipe3_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(pipe3_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(pipe3_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(pipe3_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(pipe3_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(pipe3_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(pipe3_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(pipe3_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(pipe3_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(pipe3_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(pipe3_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(pipe3_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(pipe3_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(pipe3_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(pipe3_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(pipe3_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(pipe3_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(pipe3_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(pipe3_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(pipe3_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(pipe3_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(pipe3_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(pipe3_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_next_processor_id(pipe3_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe3_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe3_io_pipe_phv_out_is_valid_processor),
    .io_table_config_0_table_depth(pipe3_io_table_config_0_table_depth),
    .io_table_config_0_table_width(pipe3_io_table_config_0_table_width),
    .io_table_config_1_table_depth(pipe3_io_table_config_1_table_depth),
    .io_table_config_1_table_width(pipe3_io_table_config_1_table_width),
    .io_key_in(pipe3_io_key_in),
    .io_key_out(pipe3_io_key_out),
    .io_addr_in(pipe3_io_addr_in),
    .io_cs_in(pipe3_io_cs_in),
    .io_data_out(pipe3_io_data_out),
    .io_w_en(pipe3_io_w_en),
    .io_w_sram_id(pipe3_io_w_sram_id),
    .io_w_addr(pipe3_io_w_addr),
    .io_w_data(pipe3_io_w_data)
  );
  MatchResultPISA pipe4 ( // @[matcher_pisa.scala 336:23]
    .clock(pipe4_clock),
    .io_pipe_phv_in_data_0(pipe4_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe4_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe4_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe4_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe4_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe4_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe4_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe4_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe4_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe4_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe4_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe4_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe4_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe4_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe4_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe4_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe4_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe4_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe4_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe4_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe4_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe4_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe4_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe4_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe4_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe4_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe4_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe4_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe4_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe4_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe4_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe4_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe4_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe4_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe4_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe4_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe4_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe4_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe4_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe4_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe4_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe4_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe4_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe4_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe4_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe4_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe4_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe4_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe4_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe4_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe4_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe4_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe4_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe4_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe4_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe4_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe4_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe4_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe4_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe4_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe4_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe4_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe4_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe4_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe4_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe4_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe4_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe4_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe4_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe4_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe4_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe4_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe4_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe4_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe4_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe4_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe4_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe4_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe4_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe4_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe4_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe4_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe4_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe4_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe4_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe4_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe4_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe4_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe4_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe4_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe4_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe4_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe4_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe4_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe4_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe4_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe4_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe4_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe4_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe4_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe4_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe4_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe4_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe4_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe4_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe4_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe4_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe4_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe4_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe4_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe4_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe4_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe4_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe4_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe4_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe4_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe4_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe4_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe4_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe4_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe4_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe4_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe4_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe4_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe4_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe4_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe4_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe4_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe4_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe4_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe4_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe4_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe4_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe4_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe4_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe4_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe4_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe4_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe4_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe4_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe4_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe4_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe4_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe4_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe4_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe4_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe4_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe4_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe4_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe4_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe4_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe4_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe4_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe4_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe4_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe4_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe4_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe4_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe4_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe4_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(pipe4_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(pipe4_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(pipe4_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(pipe4_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(pipe4_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(pipe4_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(pipe4_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(pipe4_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(pipe4_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(pipe4_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(pipe4_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(pipe4_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(pipe4_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(pipe4_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(pipe4_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(pipe4_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(pipe4_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(pipe4_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(pipe4_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(pipe4_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(pipe4_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(pipe4_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(pipe4_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(pipe4_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(pipe4_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(pipe4_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(pipe4_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(pipe4_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(pipe4_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(pipe4_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(pipe4_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(pipe4_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(pipe4_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(pipe4_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(pipe4_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(pipe4_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(pipe4_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(pipe4_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(pipe4_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(pipe4_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(pipe4_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(pipe4_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(pipe4_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(pipe4_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(pipe4_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(pipe4_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(pipe4_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(pipe4_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(pipe4_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(pipe4_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(pipe4_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(pipe4_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(pipe4_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(pipe4_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(pipe4_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(pipe4_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(pipe4_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(pipe4_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(pipe4_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(pipe4_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(pipe4_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(pipe4_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(pipe4_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(pipe4_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(pipe4_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(pipe4_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(pipe4_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(pipe4_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(pipe4_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(pipe4_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(pipe4_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(pipe4_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(pipe4_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(pipe4_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(pipe4_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(pipe4_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(pipe4_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(pipe4_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(pipe4_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(pipe4_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(pipe4_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(pipe4_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(pipe4_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(pipe4_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(pipe4_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(pipe4_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(pipe4_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(pipe4_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(pipe4_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(pipe4_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(pipe4_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(pipe4_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(pipe4_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(pipe4_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(pipe4_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(pipe4_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_next_processor_id(pipe4_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe4_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe4_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe4_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe4_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe4_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe4_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe4_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe4_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe4_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe4_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe4_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe4_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe4_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe4_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe4_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe4_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe4_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe4_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe4_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe4_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe4_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe4_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe4_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe4_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe4_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe4_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe4_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe4_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe4_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe4_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe4_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe4_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe4_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe4_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe4_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe4_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe4_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe4_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe4_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe4_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe4_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe4_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe4_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe4_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe4_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe4_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe4_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe4_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe4_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe4_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe4_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe4_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe4_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe4_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe4_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe4_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe4_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe4_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe4_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe4_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe4_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe4_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe4_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe4_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe4_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe4_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe4_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe4_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe4_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe4_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe4_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe4_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe4_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe4_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe4_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe4_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe4_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe4_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe4_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe4_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe4_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe4_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe4_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe4_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe4_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe4_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe4_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe4_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe4_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe4_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe4_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe4_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe4_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe4_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe4_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe4_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe4_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe4_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe4_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe4_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe4_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe4_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe4_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe4_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe4_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe4_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe4_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe4_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe4_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe4_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe4_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe4_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe4_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe4_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe4_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe4_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe4_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe4_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe4_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe4_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe4_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe4_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe4_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe4_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe4_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe4_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe4_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe4_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe4_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe4_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe4_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe4_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe4_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe4_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe4_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe4_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe4_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe4_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe4_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe4_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe4_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe4_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe4_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe4_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe4_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe4_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe4_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe4_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe4_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe4_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe4_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe4_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe4_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe4_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe4_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe4_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe4_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe4_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe4_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe4_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe4_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe4_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(pipe4_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(pipe4_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(pipe4_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(pipe4_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(pipe4_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(pipe4_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(pipe4_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(pipe4_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(pipe4_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(pipe4_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(pipe4_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(pipe4_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(pipe4_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(pipe4_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(pipe4_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(pipe4_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(pipe4_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(pipe4_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(pipe4_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(pipe4_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(pipe4_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(pipe4_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(pipe4_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(pipe4_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(pipe4_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(pipe4_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(pipe4_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(pipe4_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(pipe4_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(pipe4_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(pipe4_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(pipe4_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(pipe4_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(pipe4_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(pipe4_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(pipe4_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(pipe4_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(pipe4_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(pipe4_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(pipe4_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(pipe4_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(pipe4_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(pipe4_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(pipe4_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(pipe4_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(pipe4_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(pipe4_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(pipe4_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(pipe4_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(pipe4_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(pipe4_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(pipe4_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(pipe4_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(pipe4_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(pipe4_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(pipe4_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(pipe4_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(pipe4_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(pipe4_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(pipe4_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(pipe4_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(pipe4_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(pipe4_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(pipe4_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(pipe4_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(pipe4_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(pipe4_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(pipe4_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(pipe4_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(pipe4_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(pipe4_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(pipe4_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(pipe4_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(pipe4_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(pipe4_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(pipe4_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(pipe4_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(pipe4_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(pipe4_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(pipe4_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(pipe4_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(pipe4_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(pipe4_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(pipe4_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(pipe4_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(pipe4_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(pipe4_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(pipe4_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(pipe4_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(pipe4_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(pipe4_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(pipe4_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(pipe4_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(pipe4_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(pipe4_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(pipe4_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_next_processor_id(pipe4_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe4_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe4_io_pipe_phv_out_is_valid_processor),
    .io_key_config_0_field_config_0(pipe4_io_key_config_0_field_config_0),
    .io_key_config_0_field_config_1(pipe4_io_key_config_0_field_config_1),
    .io_key_config_0_field_config_2(pipe4_io_key_config_0_field_config_2),
    .io_key_config_0_field_config_3(pipe4_io_key_config_0_field_config_3),
    .io_key_config_0_field_config_4(pipe4_io_key_config_0_field_config_4),
    .io_key_config_0_field_config_5(pipe4_io_key_config_0_field_config_5),
    .io_key_config_0_field_mask_0_0(pipe4_io_key_config_0_field_mask_0_0),
    .io_key_config_0_field_mask_0_1(pipe4_io_key_config_0_field_mask_0_1),
    .io_key_config_0_field_mask_0_2(pipe4_io_key_config_0_field_mask_0_2),
    .io_key_config_0_field_mask_0_3(pipe4_io_key_config_0_field_mask_0_3),
    .io_key_config_0_field_mask_1_0(pipe4_io_key_config_0_field_mask_1_0),
    .io_key_config_0_field_mask_1_1(pipe4_io_key_config_0_field_mask_1_1),
    .io_key_config_0_field_mask_1_2(pipe4_io_key_config_0_field_mask_1_2),
    .io_key_config_0_field_mask_1_3(pipe4_io_key_config_0_field_mask_1_3),
    .io_key_config_0_field_mask_2_0(pipe4_io_key_config_0_field_mask_2_0),
    .io_key_config_0_field_mask_2_1(pipe4_io_key_config_0_field_mask_2_1),
    .io_key_config_0_field_mask_2_2(pipe4_io_key_config_0_field_mask_2_2),
    .io_key_config_0_field_mask_2_3(pipe4_io_key_config_0_field_mask_2_3),
    .io_key_config_0_field_mask_3_0(pipe4_io_key_config_0_field_mask_3_0),
    .io_key_config_0_field_mask_3_1(pipe4_io_key_config_0_field_mask_3_1),
    .io_key_config_0_field_mask_3_2(pipe4_io_key_config_0_field_mask_3_2),
    .io_key_config_0_field_mask_3_3(pipe4_io_key_config_0_field_mask_3_3),
    .io_key_config_0_field_mask_4_0(pipe4_io_key_config_0_field_mask_4_0),
    .io_key_config_0_field_mask_4_1(pipe4_io_key_config_0_field_mask_4_1),
    .io_key_config_0_field_mask_4_2(pipe4_io_key_config_0_field_mask_4_2),
    .io_key_config_0_field_mask_4_3(pipe4_io_key_config_0_field_mask_4_3),
    .io_key_config_0_field_mask_5_0(pipe4_io_key_config_0_field_mask_5_0),
    .io_key_config_0_field_mask_5_1(pipe4_io_key_config_0_field_mask_5_1),
    .io_key_config_0_field_mask_5_2(pipe4_io_key_config_0_field_mask_5_2),
    .io_key_config_0_field_mask_5_3(pipe4_io_key_config_0_field_mask_5_3),
    .io_key_config_1_field_config_0(pipe4_io_key_config_1_field_config_0),
    .io_key_config_1_field_config_1(pipe4_io_key_config_1_field_config_1),
    .io_key_config_1_field_config_2(pipe4_io_key_config_1_field_config_2),
    .io_key_config_1_field_config_3(pipe4_io_key_config_1_field_config_3),
    .io_key_config_1_field_config_4(pipe4_io_key_config_1_field_config_4),
    .io_key_config_1_field_config_5(pipe4_io_key_config_1_field_config_5),
    .io_key_config_1_field_mask_0_0(pipe4_io_key_config_1_field_mask_0_0),
    .io_key_config_1_field_mask_0_1(pipe4_io_key_config_1_field_mask_0_1),
    .io_key_config_1_field_mask_0_2(pipe4_io_key_config_1_field_mask_0_2),
    .io_key_config_1_field_mask_0_3(pipe4_io_key_config_1_field_mask_0_3),
    .io_key_config_1_field_mask_1_0(pipe4_io_key_config_1_field_mask_1_0),
    .io_key_config_1_field_mask_1_1(pipe4_io_key_config_1_field_mask_1_1),
    .io_key_config_1_field_mask_1_2(pipe4_io_key_config_1_field_mask_1_2),
    .io_key_config_1_field_mask_1_3(pipe4_io_key_config_1_field_mask_1_3),
    .io_key_config_1_field_mask_2_0(pipe4_io_key_config_1_field_mask_2_0),
    .io_key_config_1_field_mask_2_1(pipe4_io_key_config_1_field_mask_2_1),
    .io_key_config_1_field_mask_2_2(pipe4_io_key_config_1_field_mask_2_2),
    .io_key_config_1_field_mask_2_3(pipe4_io_key_config_1_field_mask_2_3),
    .io_key_config_1_field_mask_3_0(pipe4_io_key_config_1_field_mask_3_0),
    .io_key_config_1_field_mask_3_1(pipe4_io_key_config_1_field_mask_3_1),
    .io_key_config_1_field_mask_3_2(pipe4_io_key_config_1_field_mask_3_2),
    .io_key_config_1_field_mask_3_3(pipe4_io_key_config_1_field_mask_3_3),
    .io_key_config_1_field_mask_4_0(pipe4_io_key_config_1_field_mask_4_0),
    .io_key_config_1_field_mask_4_1(pipe4_io_key_config_1_field_mask_4_1),
    .io_key_config_1_field_mask_4_2(pipe4_io_key_config_1_field_mask_4_2),
    .io_key_config_1_field_mask_4_3(pipe4_io_key_config_1_field_mask_4_3),
    .io_key_config_1_field_mask_5_0(pipe4_io_key_config_1_field_mask_5_0),
    .io_key_config_1_field_mask_5_1(pipe4_io_key_config_1_field_mask_5_1),
    .io_key_config_1_field_mask_5_2(pipe4_io_key_config_1_field_mask_5_2),
    .io_key_config_1_field_mask_5_3(pipe4_io_key_config_1_field_mask_5_3),
    .io_key_in(pipe4_io_key_in),
    .io_data_in(pipe4_io_data_in),
    .io_hit(pipe4_io_hit),
    .io_match_value(pipe4_io_match_value)
  );
  assign io_pipe_phv_out_data_0 = pipe4_io_pipe_phv_out_data_0; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_1 = pipe4_io_pipe_phv_out_data_1; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_2 = pipe4_io_pipe_phv_out_data_2; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_3 = pipe4_io_pipe_phv_out_data_3; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_4 = pipe4_io_pipe_phv_out_data_4; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_5 = pipe4_io_pipe_phv_out_data_5; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_6 = pipe4_io_pipe_phv_out_data_6; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_7 = pipe4_io_pipe_phv_out_data_7; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_8 = pipe4_io_pipe_phv_out_data_8; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_9 = pipe4_io_pipe_phv_out_data_9; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_10 = pipe4_io_pipe_phv_out_data_10; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_11 = pipe4_io_pipe_phv_out_data_11; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_12 = pipe4_io_pipe_phv_out_data_12; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_13 = pipe4_io_pipe_phv_out_data_13; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_14 = pipe4_io_pipe_phv_out_data_14; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_15 = pipe4_io_pipe_phv_out_data_15; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_16 = pipe4_io_pipe_phv_out_data_16; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_17 = pipe4_io_pipe_phv_out_data_17; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_18 = pipe4_io_pipe_phv_out_data_18; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_19 = pipe4_io_pipe_phv_out_data_19; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_20 = pipe4_io_pipe_phv_out_data_20; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_21 = pipe4_io_pipe_phv_out_data_21; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_22 = pipe4_io_pipe_phv_out_data_22; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_23 = pipe4_io_pipe_phv_out_data_23; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_24 = pipe4_io_pipe_phv_out_data_24; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_25 = pipe4_io_pipe_phv_out_data_25; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_26 = pipe4_io_pipe_phv_out_data_26; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_27 = pipe4_io_pipe_phv_out_data_27; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_28 = pipe4_io_pipe_phv_out_data_28; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_29 = pipe4_io_pipe_phv_out_data_29; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_30 = pipe4_io_pipe_phv_out_data_30; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_31 = pipe4_io_pipe_phv_out_data_31; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_32 = pipe4_io_pipe_phv_out_data_32; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_33 = pipe4_io_pipe_phv_out_data_33; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_34 = pipe4_io_pipe_phv_out_data_34; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_35 = pipe4_io_pipe_phv_out_data_35; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_36 = pipe4_io_pipe_phv_out_data_36; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_37 = pipe4_io_pipe_phv_out_data_37; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_38 = pipe4_io_pipe_phv_out_data_38; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_39 = pipe4_io_pipe_phv_out_data_39; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_40 = pipe4_io_pipe_phv_out_data_40; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_41 = pipe4_io_pipe_phv_out_data_41; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_42 = pipe4_io_pipe_phv_out_data_42; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_43 = pipe4_io_pipe_phv_out_data_43; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_44 = pipe4_io_pipe_phv_out_data_44; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_45 = pipe4_io_pipe_phv_out_data_45; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_46 = pipe4_io_pipe_phv_out_data_46; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_47 = pipe4_io_pipe_phv_out_data_47; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_48 = pipe4_io_pipe_phv_out_data_48; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_49 = pipe4_io_pipe_phv_out_data_49; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_50 = pipe4_io_pipe_phv_out_data_50; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_51 = pipe4_io_pipe_phv_out_data_51; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_52 = pipe4_io_pipe_phv_out_data_52; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_53 = pipe4_io_pipe_phv_out_data_53; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_54 = pipe4_io_pipe_phv_out_data_54; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_55 = pipe4_io_pipe_phv_out_data_55; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_56 = pipe4_io_pipe_phv_out_data_56; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_57 = pipe4_io_pipe_phv_out_data_57; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_58 = pipe4_io_pipe_phv_out_data_58; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_59 = pipe4_io_pipe_phv_out_data_59; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_60 = pipe4_io_pipe_phv_out_data_60; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_61 = pipe4_io_pipe_phv_out_data_61; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_62 = pipe4_io_pipe_phv_out_data_62; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_63 = pipe4_io_pipe_phv_out_data_63; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_64 = pipe4_io_pipe_phv_out_data_64; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_65 = pipe4_io_pipe_phv_out_data_65; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_66 = pipe4_io_pipe_phv_out_data_66; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_67 = pipe4_io_pipe_phv_out_data_67; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_68 = pipe4_io_pipe_phv_out_data_68; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_69 = pipe4_io_pipe_phv_out_data_69; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_70 = pipe4_io_pipe_phv_out_data_70; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_71 = pipe4_io_pipe_phv_out_data_71; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_72 = pipe4_io_pipe_phv_out_data_72; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_73 = pipe4_io_pipe_phv_out_data_73; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_74 = pipe4_io_pipe_phv_out_data_74; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_75 = pipe4_io_pipe_phv_out_data_75; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_76 = pipe4_io_pipe_phv_out_data_76; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_77 = pipe4_io_pipe_phv_out_data_77; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_78 = pipe4_io_pipe_phv_out_data_78; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_79 = pipe4_io_pipe_phv_out_data_79; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_80 = pipe4_io_pipe_phv_out_data_80; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_81 = pipe4_io_pipe_phv_out_data_81; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_82 = pipe4_io_pipe_phv_out_data_82; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_83 = pipe4_io_pipe_phv_out_data_83; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_84 = pipe4_io_pipe_phv_out_data_84; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_85 = pipe4_io_pipe_phv_out_data_85; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_86 = pipe4_io_pipe_phv_out_data_86; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_87 = pipe4_io_pipe_phv_out_data_87; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_88 = pipe4_io_pipe_phv_out_data_88; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_89 = pipe4_io_pipe_phv_out_data_89; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_90 = pipe4_io_pipe_phv_out_data_90; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_91 = pipe4_io_pipe_phv_out_data_91; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_92 = pipe4_io_pipe_phv_out_data_92; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_93 = pipe4_io_pipe_phv_out_data_93; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_94 = pipe4_io_pipe_phv_out_data_94; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_95 = pipe4_io_pipe_phv_out_data_95; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_96 = pipe4_io_pipe_phv_out_data_96; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_97 = pipe4_io_pipe_phv_out_data_97; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_98 = pipe4_io_pipe_phv_out_data_98; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_99 = pipe4_io_pipe_phv_out_data_99; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_100 = pipe4_io_pipe_phv_out_data_100; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_101 = pipe4_io_pipe_phv_out_data_101; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_102 = pipe4_io_pipe_phv_out_data_102; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_103 = pipe4_io_pipe_phv_out_data_103; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_104 = pipe4_io_pipe_phv_out_data_104; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_105 = pipe4_io_pipe_phv_out_data_105; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_106 = pipe4_io_pipe_phv_out_data_106; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_107 = pipe4_io_pipe_phv_out_data_107; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_108 = pipe4_io_pipe_phv_out_data_108; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_109 = pipe4_io_pipe_phv_out_data_109; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_110 = pipe4_io_pipe_phv_out_data_110; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_111 = pipe4_io_pipe_phv_out_data_111; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_112 = pipe4_io_pipe_phv_out_data_112; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_113 = pipe4_io_pipe_phv_out_data_113; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_114 = pipe4_io_pipe_phv_out_data_114; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_115 = pipe4_io_pipe_phv_out_data_115; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_116 = pipe4_io_pipe_phv_out_data_116; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_117 = pipe4_io_pipe_phv_out_data_117; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_118 = pipe4_io_pipe_phv_out_data_118; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_119 = pipe4_io_pipe_phv_out_data_119; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_120 = pipe4_io_pipe_phv_out_data_120; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_121 = pipe4_io_pipe_phv_out_data_121; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_122 = pipe4_io_pipe_phv_out_data_122; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_123 = pipe4_io_pipe_phv_out_data_123; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_124 = pipe4_io_pipe_phv_out_data_124; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_125 = pipe4_io_pipe_phv_out_data_125; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_126 = pipe4_io_pipe_phv_out_data_126; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_127 = pipe4_io_pipe_phv_out_data_127; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_128 = pipe4_io_pipe_phv_out_data_128; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_129 = pipe4_io_pipe_phv_out_data_129; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_130 = pipe4_io_pipe_phv_out_data_130; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_131 = pipe4_io_pipe_phv_out_data_131; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_132 = pipe4_io_pipe_phv_out_data_132; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_133 = pipe4_io_pipe_phv_out_data_133; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_134 = pipe4_io_pipe_phv_out_data_134; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_135 = pipe4_io_pipe_phv_out_data_135; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_136 = pipe4_io_pipe_phv_out_data_136; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_137 = pipe4_io_pipe_phv_out_data_137; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_138 = pipe4_io_pipe_phv_out_data_138; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_139 = pipe4_io_pipe_phv_out_data_139; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_140 = pipe4_io_pipe_phv_out_data_140; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_141 = pipe4_io_pipe_phv_out_data_141; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_142 = pipe4_io_pipe_phv_out_data_142; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_143 = pipe4_io_pipe_phv_out_data_143; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_144 = pipe4_io_pipe_phv_out_data_144; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_145 = pipe4_io_pipe_phv_out_data_145; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_146 = pipe4_io_pipe_phv_out_data_146; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_147 = pipe4_io_pipe_phv_out_data_147; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_148 = pipe4_io_pipe_phv_out_data_148; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_149 = pipe4_io_pipe_phv_out_data_149; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_150 = pipe4_io_pipe_phv_out_data_150; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_151 = pipe4_io_pipe_phv_out_data_151; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_152 = pipe4_io_pipe_phv_out_data_152; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_153 = pipe4_io_pipe_phv_out_data_153; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_154 = pipe4_io_pipe_phv_out_data_154; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_155 = pipe4_io_pipe_phv_out_data_155; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_156 = pipe4_io_pipe_phv_out_data_156; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_157 = pipe4_io_pipe_phv_out_data_157; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_158 = pipe4_io_pipe_phv_out_data_158; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_159 = pipe4_io_pipe_phv_out_data_159; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_160 = pipe4_io_pipe_phv_out_data_160; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_161 = pipe4_io_pipe_phv_out_data_161; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_162 = pipe4_io_pipe_phv_out_data_162; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_163 = pipe4_io_pipe_phv_out_data_163; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_164 = pipe4_io_pipe_phv_out_data_164; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_165 = pipe4_io_pipe_phv_out_data_165; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_166 = pipe4_io_pipe_phv_out_data_166; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_167 = pipe4_io_pipe_phv_out_data_167; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_168 = pipe4_io_pipe_phv_out_data_168; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_169 = pipe4_io_pipe_phv_out_data_169; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_170 = pipe4_io_pipe_phv_out_data_170; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_171 = pipe4_io_pipe_phv_out_data_171; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_172 = pipe4_io_pipe_phv_out_data_172; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_173 = pipe4_io_pipe_phv_out_data_173; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_174 = pipe4_io_pipe_phv_out_data_174; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_175 = pipe4_io_pipe_phv_out_data_175; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_176 = pipe4_io_pipe_phv_out_data_176; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_177 = pipe4_io_pipe_phv_out_data_177; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_178 = pipe4_io_pipe_phv_out_data_178; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_179 = pipe4_io_pipe_phv_out_data_179; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_180 = pipe4_io_pipe_phv_out_data_180; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_181 = pipe4_io_pipe_phv_out_data_181; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_182 = pipe4_io_pipe_phv_out_data_182; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_183 = pipe4_io_pipe_phv_out_data_183; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_184 = pipe4_io_pipe_phv_out_data_184; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_185 = pipe4_io_pipe_phv_out_data_185; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_186 = pipe4_io_pipe_phv_out_data_186; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_187 = pipe4_io_pipe_phv_out_data_187; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_188 = pipe4_io_pipe_phv_out_data_188; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_189 = pipe4_io_pipe_phv_out_data_189; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_190 = pipe4_io_pipe_phv_out_data_190; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_191 = pipe4_io_pipe_phv_out_data_191; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_192 = pipe4_io_pipe_phv_out_data_192; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_193 = pipe4_io_pipe_phv_out_data_193; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_194 = pipe4_io_pipe_phv_out_data_194; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_195 = pipe4_io_pipe_phv_out_data_195; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_196 = pipe4_io_pipe_phv_out_data_196; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_197 = pipe4_io_pipe_phv_out_data_197; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_198 = pipe4_io_pipe_phv_out_data_198; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_199 = pipe4_io_pipe_phv_out_data_199; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_200 = pipe4_io_pipe_phv_out_data_200; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_201 = pipe4_io_pipe_phv_out_data_201; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_202 = pipe4_io_pipe_phv_out_data_202; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_203 = pipe4_io_pipe_phv_out_data_203; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_204 = pipe4_io_pipe_phv_out_data_204; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_205 = pipe4_io_pipe_phv_out_data_205; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_206 = pipe4_io_pipe_phv_out_data_206; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_207 = pipe4_io_pipe_phv_out_data_207; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_208 = pipe4_io_pipe_phv_out_data_208; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_209 = pipe4_io_pipe_phv_out_data_209; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_210 = pipe4_io_pipe_phv_out_data_210; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_211 = pipe4_io_pipe_phv_out_data_211; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_212 = pipe4_io_pipe_phv_out_data_212; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_213 = pipe4_io_pipe_phv_out_data_213; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_214 = pipe4_io_pipe_phv_out_data_214; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_215 = pipe4_io_pipe_phv_out_data_215; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_216 = pipe4_io_pipe_phv_out_data_216; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_217 = pipe4_io_pipe_phv_out_data_217; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_218 = pipe4_io_pipe_phv_out_data_218; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_219 = pipe4_io_pipe_phv_out_data_219; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_220 = pipe4_io_pipe_phv_out_data_220; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_221 = pipe4_io_pipe_phv_out_data_221; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_222 = pipe4_io_pipe_phv_out_data_222; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_223 = pipe4_io_pipe_phv_out_data_223; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_224 = pipe4_io_pipe_phv_out_data_224; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_225 = pipe4_io_pipe_phv_out_data_225; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_226 = pipe4_io_pipe_phv_out_data_226; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_227 = pipe4_io_pipe_phv_out_data_227; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_228 = pipe4_io_pipe_phv_out_data_228; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_229 = pipe4_io_pipe_phv_out_data_229; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_230 = pipe4_io_pipe_phv_out_data_230; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_231 = pipe4_io_pipe_phv_out_data_231; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_232 = pipe4_io_pipe_phv_out_data_232; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_233 = pipe4_io_pipe_phv_out_data_233; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_234 = pipe4_io_pipe_phv_out_data_234; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_235 = pipe4_io_pipe_phv_out_data_235; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_236 = pipe4_io_pipe_phv_out_data_236; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_237 = pipe4_io_pipe_phv_out_data_237; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_238 = pipe4_io_pipe_phv_out_data_238; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_239 = pipe4_io_pipe_phv_out_data_239; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_240 = pipe4_io_pipe_phv_out_data_240; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_241 = pipe4_io_pipe_phv_out_data_241; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_242 = pipe4_io_pipe_phv_out_data_242; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_243 = pipe4_io_pipe_phv_out_data_243; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_244 = pipe4_io_pipe_phv_out_data_244; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_245 = pipe4_io_pipe_phv_out_data_245; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_246 = pipe4_io_pipe_phv_out_data_246; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_247 = pipe4_io_pipe_phv_out_data_247; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_248 = pipe4_io_pipe_phv_out_data_248; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_249 = pipe4_io_pipe_phv_out_data_249; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_250 = pipe4_io_pipe_phv_out_data_250; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_251 = pipe4_io_pipe_phv_out_data_251; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_252 = pipe4_io_pipe_phv_out_data_252; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_253 = pipe4_io_pipe_phv_out_data_253; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_254 = pipe4_io_pipe_phv_out_data_254; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_255 = pipe4_io_pipe_phv_out_data_255; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_next_processor_id = pipe4_io_pipe_phv_out_next_processor_id; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_next_config_id = pipe4_io_pipe_phv_out_next_config_id; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_is_valid_processor = pipe4_io_pipe_phv_out_is_valid_processor; // @[matcher_pisa.scala 359:26]
  assign io_hit = pipe4_io_hit; // @[matcher_pisa.scala 360:26]
  assign io_match_value = pipe4_io_match_value; // @[matcher_pisa.scala 361:26]
  assign pipe1_clock = clock;
  assign pipe1_io_pipe_phv_in_data_0 = io_pipe_phv_in_data_0; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_1 = io_pipe_phv_in_data_1; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_2 = io_pipe_phv_in_data_2; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_3 = io_pipe_phv_in_data_3; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_4 = io_pipe_phv_in_data_4; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_5 = io_pipe_phv_in_data_5; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_6 = io_pipe_phv_in_data_6; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_7 = io_pipe_phv_in_data_7; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_8 = io_pipe_phv_in_data_8; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_9 = io_pipe_phv_in_data_9; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_10 = io_pipe_phv_in_data_10; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_11 = io_pipe_phv_in_data_11; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_12 = io_pipe_phv_in_data_12; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_13 = io_pipe_phv_in_data_13; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_14 = io_pipe_phv_in_data_14; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_15 = io_pipe_phv_in_data_15; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_16 = io_pipe_phv_in_data_16; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_17 = io_pipe_phv_in_data_17; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_18 = io_pipe_phv_in_data_18; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_19 = io_pipe_phv_in_data_19; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_20 = io_pipe_phv_in_data_20; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_21 = io_pipe_phv_in_data_21; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_22 = io_pipe_phv_in_data_22; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_23 = io_pipe_phv_in_data_23; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_24 = io_pipe_phv_in_data_24; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_25 = io_pipe_phv_in_data_25; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_26 = io_pipe_phv_in_data_26; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_27 = io_pipe_phv_in_data_27; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_28 = io_pipe_phv_in_data_28; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_29 = io_pipe_phv_in_data_29; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_30 = io_pipe_phv_in_data_30; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_31 = io_pipe_phv_in_data_31; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_32 = io_pipe_phv_in_data_32; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_33 = io_pipe_phv_in_data_33; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_34 = io_pipe_phv_in_data_34; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_35 = io_pipe_phv_in_data_35; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_36 = io_pipe_phv_in_data_36; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_37 = io_pipe_phv_in_data_37; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_38 = io_pipe_phv_in_data_38; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_39 = io_pipe_phv_in_data_39; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_40 = io_pipe_phv_in_data_40; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_41 = io_pipe_phv_in_data_41; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_42 = io_pipe_phv_in_data_42; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_43 = io_pipe_phv_in_data_43; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_44 = io_pipe_phv_in_data_44; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_45 = io_pipe_phv_in_data_45; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_46 = io_pipe_phv_in_data_46; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_47 = io_pipe_phv_in_data_47; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_48 = io_pipe_phv_in_data_48; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_49 = io_pipe_phv_in_data_49; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_50 = io_pipe_phv_in_data_50; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_51 = io_pipe_phv_in_data_51; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_52 = io_pipe_phv_in_data_52; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_53 = io_pipe_phv_in_data_53; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_54 = io_pipe_phv_in_data_54; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_55 = io_pipe_phv_in_data_55; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_56 = io_pipe_phv_in_data_56; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_57 = io_pipe_phv_in_data_57; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_58 = io_pipe_phv_in_data_58; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_59 = io_pipe_phv_in_data_59; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_60 = io_pipe_phv_in_data_60; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_61 = io_pipe_phv_in_data_61; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_62 = io_pipe_phv_in_data_62; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_63 = io_pipe_phv_in_data_63; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_64 = io_pipe_phv_in_data_64; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_65 = io_pipe_phv_in_data_65; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_66 = io_pipe_phv_in_data_66; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_67 = io_pipe_phv_in_data_67; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_68 = io_pipe_phv_in_data_68; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_69 = io_pipe_phv_in_data_69; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_70 = io_pipe_phv_in_data_70; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_71 = io_pipe_phv_in_data_71; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_72 = io_pipe_phv_in_data_72; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_73 = io_pipe_phv_in_data_73; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_74 = io_pipe_phv_in_data_74; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_75 = io_pipe_phv_in_data_75; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_76 = io_pipe_phv_in_data_76; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_77 = io_pipe_phv_in_data_77; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_78 = io_pipe_phv_in_data_78; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_79 = io_pipe_phv_in_data_79; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_80 = io_pipe_phv_in_data_80; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_81 = io_pipe_phv_in_data_81; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_82 = io_pipe_phv_in_data_82; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_83 = io_pipe_phv_in_data_83; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_84 = io_pipe_phv_in_data_84; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_85 = io_pipe_phv_in_data_85; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_86 = io_pipe_phv_in_data_86; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_87 = io_pipe_phv_in_data_87; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_88 = io_pipe_phv_in_data_88; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_89 = io_pipe_phv_in_data_89; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_90 = io_pipe_phv_in_data_90; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_91 = io_pipe_phv_in_data_91; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_92 = io_pipe_phv_in_data_92; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_93 = io_pipe_phv_in_data_93; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_94 = io_pipe_phv_in_data_94; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_95 = io_pipe_phv_in_data_95; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_96 = io_pipe_phv_in_data_96; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_97 = io_pipe_phv_in_data_97; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_98 = io_pipe_phv_in_data_98; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_99 = io_pipe_phv_in_data_99; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_100 = io_pipe_phv_in_data_100; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_101 = io_pipe_phv_in_data_101; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_102 = io_pipe_phv_in_data_102; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_103 = io_pipe_phv_in_data_103; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_104 = io_pipe_phv_in_data_104; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_105 = io_pipe_phv_in_data_105; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_106 = io_pipe_phv_in_data_106; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_107 = io_pipe_phv_in_data_107; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_108 = io_pipe_phv_in_data_108; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_109 = io_pipe_phv_in_data_109; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_110 = io_pipe_phv_in_data_110; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_111 = io_pipe_phv_in_data_111; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_112 = io_pipe_phv_in_data_112; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_113 = io_pipe_phv_in_data_113; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_114 = io_pipe_phv_in_data_114; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_115 = io_pipe_phv_in_data_115; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_116 = io_pipe_phv_in_data_116; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_117 = io_pipe_phv_in_data_117; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_118 = io_pipe_phv_in_data_118; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_119 = io_pipe_phv_in_data_119; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_120 = io_pipe_phv_in_data_120; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_121 = io_pipe_phv_in_data_121; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_122 = io_pipe_phv_in_data_122; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_123 = io_pipe_phv_in_data_123; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_124 = io_pipe_phv_in_data_124; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_125 = io_pipe_phv_in_data_125; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_126 = io_pipe_phv_in_data_126; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_127 = io_pipe_phv_in_data_127; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_128 = io_pipe_phv_in_data_128; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_129 = io_pipe_phv_in_data_129; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_130 = io_pipe_phv_in_data_130; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_131 = io_pipe_phv_in_data_131; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_132 = io_pipe_phv_in_data_132; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_133 = io_pipe_phv_in_data_133; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_134 = io_pipe_phv_in_data_134; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_135 = io_pipe_phv_in_data_135; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_136 = io_pipe_phv_in_data_136; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_137 = io_pipe_phv_in_data_137; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_138 = io_pipe_phv_in_data_138; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_139 = io_pipe_phv_in_data_139; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_140 = io_pipe_phv_in_data_140; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_141 = io_pipe_phv_in_data_141; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_142 = io_pipe_phv_in_data_142; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_143 = io_pipe_phv_in_data_143; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_144 = io_pipe_phv_in_data_144; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_145 = io_pipe_phv_in_data_145; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_146 = io_pipe_phv_in_data_146; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_147 = io_pipe_phv_in_data_147; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_148 = io_pipe_phv_in_data_148; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_149 = io_pipe_phv_in_data_149; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_150 = io_pipe_phv_in_data_150; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_151 = io_pipe_phv_in_data_151; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_152 = io_pipe_phv_in_data_152; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_153 = io_pipe_phv_in_data_153; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_154 = io_pipe_phv_in_data_154; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_155 = io_pipe_phv_in_data_155; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_156 = io_pipe_phv_in_data_156; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_157 = io_pipe_phv_in_data_157; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_158 = io_pipe_phv_in_data_158; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_159 = io_pipe_phv_in_data_159; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_160 = io_pipe_phv_in_data_160; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_161 = io_pipe_phv_in_data_161; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_162 = io_pipe_phv_in_data_162; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_163 = io_pipe_phv_in_data_163; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_164 = io_pipe_phv_in_data_164; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_165 = io_pipe_phv_in_data_165; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_166 = io_pipe_phv_in_data_166; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_167 = io_pipe_phv_in_data_167; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_168 = io_pipe_phv_in_data_168; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_169 = io_pipe_phv_in_data_169; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_170 = io_pipe_phv_in_data_170; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_171 = io_pipe_phv_in_data_171; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_172 = io_pipe_phv_in_data_172; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_173 = io_pipe_phv_in_data_173; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_174 = io_pipe_phv_in_data_174; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_175 = io_pipe_phv_in_data_175; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_176 = io_pipe_phv_in_data_176; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_177 = io_pipe_phv_in_data_177; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_178 = io_pipe_phv_in_data_178; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_179 = io_pipe_phv_in_data_179; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_180 = io_pipe_phv_in_data_180; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_181 = io_pipe_phv_in_data_181; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_182 = io_pipe_phv_in_data_182; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_183 = io_pipe_phv_in_data_183; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_184 = io_pipe_phv_in_data_184; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_185 = io_pipe_phv_in_data_185; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_186 = io_pipe_phv_in_data_186; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_187 = io_pipe_phv_in_data_187; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_188 = io_pipe_phv_in_data_188; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_189 = io_pipe_phv_in_data_189; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_190 = io_pipe_phv_in_data_190; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_191 = io_pipe_phv_in_data_191; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_192 = io_pipe_phv_in_data_192; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_193 = io_pipe_phv_in_data_193; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_194 = io_pipe_phv_in_data_194; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_195 = io_pipe_phv_in_data_195; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_196 = io_pipe_phv_in_data_196; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_197 = io_pipe_phv_in_data_197; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_198 = io_pipe_phv_in_data_198; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_199 = io_pipe_phv_in_data_199; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_200 = io_pipe_phv_in_data_200; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_201 = io_pipe_phv_in_data_201; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_202 = io_pipe_phv_in_data_202; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_203 = io_pipe_phv_in_data_203; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_204 = io_pipe_phv_in_data_204; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_205 = io_pipe_phv_in_data_205; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_206 = io_pipe_phv_in_data_206; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_207 = io_pipe_phv_in_data_207; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_208 = io_pipe_phv_in_data_208; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_209 = io_pipe_phv_in_data_209; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_210 = io_pipe_phv_in_data_210; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_211 = io_pipe_phv_in_data_211; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_212 = io_pipe_phv_in_data_212; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_213 = io_pipe_phv_in_data_213; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_214 = io_pipe_phv_in_data_214; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_215 = io_pipe_phv_in_data_215; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_216 = io_pipe_phv_in_data_216; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_217 = io_pipe_phv_in_data_217; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_218 = io_pipe_phv_in_data_218; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_219 = io_pipe_phv_in_data_219; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_220 = io_pipe_phv_in_data_220; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_221 = io_pipe_phv_in_data_221; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_222 = io_pipe_phv_in_data_222; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_223 = io_pipe_phv_in_data_223; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_224 = io_pipe_phv_in_data_224; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_225 = io_pipe_phv_in_data_225; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_226 = io_pipe_phv_in_data_226; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_227 = io_pipe_phv_in_data_227; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_228 = io_pipe_phv_in_data_228; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_229 = io_pipe_phv_in_data_229; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_230 = io_pipe_phv_in_data_230; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_231 = io_pipe_phv_in_data_231; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_232 = io_pipe_phv_in_data_232; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_233 = io_pipe_phv_in_data_233; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_234 = io_pipe_phv_in_data_234; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_235 = io_pipe_phv_in_data_235; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_236 = io_pipe_phv_in_data_236; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_237 = io_pipe_phv_in_data_237; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_238 = io_pipe_phv_in_data_238; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_239 = io_pipe_phv_in_data_239; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_240 = io_pipe_phv_in_data_240; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_241 = io_pipe_phv_in_data_241; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_242 = io_pipe_phv_in_data_242; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_243 = io_pipe_phv_in_data_243; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_244 = io_pipe_phv_in_data_244; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_245 = io_pipe_phv_in_data_245; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_246 = io_pipe_phv_in_data_246; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_247 = io_pipe_phv_in_data_247; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_248 = io_pipe_phv_in_data_248; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_249 = io_pipe_phv_in_data_249; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_250 = io_pipe_phv_in_data_250; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_251 = io_pipe_phv_in_data_251; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_252 = io_pipe_phv_in_data_252; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_253 = io_pipe_phv_in_data_253; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_254 = io_pipe_phv_in_data_254; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_255 = io_pipe_phv_in_data_255; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_next_processor_id = io_pipe_phv_in_next_processor_id; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_next_config_id = io_pipe_phv_in_next_config_id; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_is_valid_processor = io_pipe_phv_in_is_valid_processor; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_key_config_0_field_config_0 = key_config_0_field_config_0; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_config_1 = key_config_0_field_config_1; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_config_2 = key_config_0_field_config_2; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_config_3 = key_config_0_field_config_3; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_config_4 = key_config_0_field_config_4; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_config_5 = key_config_0_field_config_5; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_mask_0_0 = key_config_0_field_mask_0_0; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_mask_0_1 = key_config_0_field_mask_0_1; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_mask_0_2 = key_config_0_field_mask_0_2; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_mask_0_3 = key_config_0_field_mask_0_3; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_mask_1_0 = key_config_0_field_mask_1_0; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_mask_1_1 = key_config_0_field_mask_1_1; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_mask_1_2 = key_config_0_field_mask_1_2; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_mask_1_3 = key_config_0_field_mask_1_3; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_mask_2_0 = key_config_0_field_mask_2_0; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_mask_2_1 = key_config_0_field_mask_2_1; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_mask_2_2 = key_config_0_field_mask_2_2; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_mask_2_3 = key_config_0_field_mask_2_3; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_mask_3_0 = key_config_0_field_mask_3_0; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_mask_3_1 = key_config_0_field_mask_3_1; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_mask_3_2 = key_config_0_field_mask_3_2; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_mask_3_3 = key_config_0_field_mask_3_3; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_mask_4_0 = key_config_0_field_mask_4_0; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_mask_4_1 = key_config_0_field_mask_4_1; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_mask_4_2 = key_config_0_field_mask_4_2; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_mask_4_3 = key_config_0_field_mask_4_3; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_mask_5_0 = key_config_0_field_mask_5_0; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_mask_5_1 = key_config_0_field_mask_5_1; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_mask_5_2 = key_config_0_field_mask_5_2; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_mask_5_3 = key_config_0_field_mask_5_3; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_id_0_0 = key_config_0_field_id_0_0; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_id_0_1 = key_config_0_field_id_0_1; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_id_0_2 = key_config_0_field_id_0_2; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_id_0_3 = key_config_0_field_id_0_3; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_id_1_0 = key_config_0_field_id_1_0; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_id_1_1 = key_config_0_field_id_1_1; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_id_1_2 = key_config_0_field_id_1_2; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_id_1_3 = key_config_0_field_id_1_3; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_id_2_0 = key_config_0_field_id_2_0; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_id_2_1 = key_config_0_field_id_2_1; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_id_2_2 = key_config_0_field_id_2_2; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_id_2_3 = key_config_0_field_id_2_3; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_id_3_0 = key_config_0_field_id_3_0; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_id_3_1 = key_config_0_field_id_3_1; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_id_3_2 = key_config_0_field_id_3_2; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_id_3_3 = key_config_0_field_id_3_3; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_id_4_0 = key_config_0_field_id_4_0; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_id_4_1 = key_config_0_field_id_4_1; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_id_4_2 = key_config_0_field_id_4_2; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_id_4_3 = key_config_0_field_id_4_3; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_id_5_0 = key_config_0_field_id_5_0; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_id_5_1 = key_config_0_field_id_5_1; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_id_5_2 = key_config_0_field_id_5_2; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_id_5_3 = key_config_0_field_id_5_3; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_config_0 = key_config_1_field_config_0; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_config_1 = key_config_1_field_config_1; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_config_2 = key_config_1_field_config_2; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_config_3 = key_config_1_field_config_3; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_config_4 = key_config_1_field_config_4; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_config_5 = key_config_1_field_config_5; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_mask_0_0 = key_config_1_field_mask_0_0; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_mask_0_1 = key_config_1_field_mask_0_1; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_mask_0_2 = key_config_1_field_mask_0_2; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_mask_0_3 = key_config_1_field_mask_0_3; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_mask_1_0 = key_config_1_field_mask_1_0; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_mask_1_1 = key_config_1_field_mask_1_1; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_mask_1_2 = key_config_1_field_mask_1_2; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_mask_1_3 = key_config_1_field_mask_1_3; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_mask_2_0 = key_config_1_field_mask_2_0; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_mask_2_1 = key_config_1_field_mask_2_1; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_mask_2_2 = key_config_1_field_mask_2_2; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_mask_2_3 = key_config_1_field_mask_2_3; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_mask_3_0 = key_config_1_field_mask_3_0; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_mask_3_1 = key_config_1_field_mask_3_1; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_mask_3_2 = key_config_1_field_mask_3_2; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_mask_3_3 = key_config_1_field_mask_3_3; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_mask_4_0 = key_config_1_field_mask_4_0; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_mask_4_1 = key_config_1_field_mask_4_1; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_mask_4_2 = key_config_1_field_mask_4_2; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_mask_4_3 = key_config_1_field_mask_4_3; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_mask_5_0 = key_config_1_field_mask_5_0; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_mask_5_1 = key_config_1_field_mask_5_1; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_mask_5_2 = key_config_1_field_mask_5_2; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_mask_5_3 = key_config_1_field_mask_5_3; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_id_0_0 = key_config_1_field_id_0_0; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_id_0_1 = key_config_1_field_id_0_1; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_id_0_2 = key_config_1_field_id_0_2; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_id_0_3 = key_config_1_field_id_0_3; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_id_1_0 = key_config_1_field_id_1_0; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_id_1_1 = key_config_1_field_id_1_1; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_id_1_2 = key_config_1_field_id_1_2; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_id_1_3 = key_config_1_field_id_1_3; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_id_2_0 = key_config_1_field_id_2_0; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_id_2_1 = key_config_1_field_id_2_1; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_id_2_2 = key_config_1_field_id_2_2; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_id_2_3 = key_config_1_field_id_2_3; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_id_3_0 = key_config_1_field_id_3_0; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_id_3_1 = key_config_1_field_id_3_1; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_id_3_2 = key_config_1_field_id_3_2; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_id_3_3 = key_config_1_field_id_3_3; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_id_4_0 = key_config_1_field_id_4_0; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_id_4_1 = key_config_1_field_id_4_1; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_id_4_2 = key_config_1_field_id_4_2; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_id_4_3 = key_config_1_field_id_4_3; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_id_5_0 = key_config_1_field_id_5_0; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_id_5_1 = key_config_1_field_id_5_1; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_id_5_2 = key_config_1_field_id_5_2; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_id_5_3 = key_config_1_field_id_5_3; // @[matcher_pisa.scala 339:26]
  assign pipe2_clock = clock;
  assign pipe2_io_pipe_phv_in_data_0 = pipe1_io_pipe_phv_out_data_0; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_1 = pipe1_io_pipe_phv_out_data_1; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_2 = pipe1_io_pipe_phv_out_data_2; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_3 = pipe1_io_pipe_phv_out_data_3; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_4 = pipe1_io_pipe_phv_out_data_4; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_5 = pipe1_io_pipe_phv_out_data_5; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_6 = pipe1_io_pipe_phv_out_data_6; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_7 = pipe1_io_pipe_phv_out_data_7; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_8 = pipe1_io_pipe_phv_out_data_8; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_9 = pipe1_io_pipe_phv_out_data_9; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_10 = pipe1_io_pipe_phv_out_data_10; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_11 = pipe1_io_pipe_phv_out_data_11; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_12 = pipe1_io_pipe_phv_out_data_12; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_13 = pipe1_io_pipe_phv_out_data_13; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_14 = pipe1_io_pipe_phv_out_data_14; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_15 = pipe1_io_pipe_phv_out_data_15; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_16 = pipe1_io_pipe_phv_out_data_16; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_17 = pipe1_io_pipe_phv_out_data_17; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_18 = pipe1_io_pipe_phv_out_data_18; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_19 = pipe1_io_pipe_phv_out_data_19; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_20 = pipe1_io_pipe_phv_out_data_20; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_21 = pipe1_io_pipe_phv_out_data_21; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_22 = pipe1_io_pipe_phv_out_data_22; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_23 = pipe1_io_pipe_phv_out_data_23; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_24 = pipe1_io_pipe_phv_out_data_24; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_25 = pipe1_io_pipe_phv_out_data_25; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_26 = pipe1_io_pipe_phv_out_data_26; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_27 = pipe1_io_pipe_phv_out_data_27; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_28 = pipe1_io_pipe_phv_out_data_28; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_29 = pipe1_io_pipe_phv_out_data_29; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_30 = pipe1_io_pipe_phv_out_data_30; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_31 = pipe1_io_pipe_phv_out_data_31; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_32 = pipe1_io_pipe_phv_out_data_32; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_33 = pipe1_io_pipe_phv_out_data_33; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_34 = pipe1_io_pipe_phv_out_data_34; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_35 = pipe1_io_pipe_phv_out_data_35; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_36 = pipe1_io_pipe_phv_out_data_36; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_37 = pipe1_io_pipe_phv_out_data_37; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_38 = pipe1_io_pipe_phv_out_data_38; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_39 = pipe1_io_pipe_phv_out_data_39; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_40 = pipe1_io_pipe_phv_out_data_40; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_41 = pipe1_io_pipe_phv_out_data_41; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_42 = pipe1_io_pipe_phv_out_data_42; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_43 = pipe1_io_pipe_phv_out_data_43; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_44 = pipe1_io_pipe_phv_out_data_44; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_45 = pipe1_io_pipe_phv_out_data_45; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_46 = pipe1_io_pipe_phv_out_data_46; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_47 = pipe1_io_pipe_phv_out_data_47; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_48 = pipe1_io_pipe_phv_out_data_48; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_49 = pipe1_io_pipe_phv_out_data_49; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_50 = pipe1_io_pipe_phv_out_data_50; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_51 = pipe1_io_pipe_phv_out_data_51; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_52 = pipe1_io_pipe_phv_out_data_52; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_53 = pipe1_io_pipe_phv_out_data_53; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_54 = pipe1_io_pipe_phv_out_data_54; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_55 = pipe1_io_pipe_phv_out_data_55; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_56 = pipe1_io_pipe_phv_out_data_56; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_57 = pipe1_io_pipe_phv_out_data_57; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_58 = pipe1_io_pipe_phv_out_data_58; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_59 = pipe1_io_pipe_phv_out_data_59; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_60 = pipe1_io_pipe_phv_out_data_60; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_61 = pipe1_io_pipe_phv_out_data_61; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_62 = pipe1_io_pipe_phv_out_data_62; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_63 = pipe1_io_pipe_phv_out_data_63; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_64 = pipe1_io_pipe_phv_out_data_64; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_65 = pipe1_io_pipe_phv_out_data_65; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_66 = pipe1_io_pipe_phv_out_data_66; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_67 = pipe1_io_pipe_phv_out_data_67; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_68 = pipe1_io_pipe_phv_out_data_68; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_69 = pipe1_io_pipe_phv_out_data_69; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_70 = pipe1_io_pipe_phv_out_data_70; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_71 = pipe1_io_pipe_phv_out_data_71; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_72 = pipe1_io_pipe_phv_out_data_72; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_73 = pipe1_io_pipe_phv_out_data_73; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_74 = pipe1_io_pipe_phv_out_data_74; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_75 = pipe1_io_pipe_phv_out_data_75; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_76 = pipe1_io_pipe_phv_out_data_76; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_77 = pipe1_io_pipe_phv_out_data_77; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_78 = pipe1_io_pipe_phv_out_data_78; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_79 = pipe1_io_pipe_phv_out_data_79; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_80 = pipe1_io_pipe_phv_out_data_80; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_81 = pipe1_io_pipe_phv_out_data_81; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_82 = pipe1_io_pipe_phv_out_data_82; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_83 = pipe1_io_pipe_phv_out_data_83; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_84 = pipe1_io_pipe_phv_out_data_84; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_85 = pipe1_io_pipe_phv_out_data_85; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_86 = pipe1_io_pipe_phv_out_data_86; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_87 = pipe1_io_pipe_phv_out_data_87; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_88 = pipe1_io_pipe_phv_out_data_88; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_89 = pipe1_io_pipe_phv_out_data_89; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_90 = pipe1_io_pipe_phv_out_data_90; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_91 = pipe1_io_pipe_phv_out_data_91; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_92 = pipe1_io_pipe_phv_out_data_92; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_93 = pipe1_io_pipe_phv_out_data_93; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_94 = pipe1_io_pipe_phv_out_data_94; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_95 = pipe1_io_pipe_phv_out_data_95; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_96 = pipe1_io_pipe_phv_out_data_96; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_97 = pipe1_io_pipe_phv_out_data_97; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_98 = pipe1_io_pipe_phv_out_data_98; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_99 = pipe1_io_pipe_phv_out_data_99; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_100 = pipe1_io_pipe_phv_out_data_100; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_101 = pipe1_io_pipe_phv_out_data_101; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_102 = pipe1_io_pipe_phv_out_data_102; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_103 = pipe1_io_pipe_phv_out_data_103; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_104 = pipe1_io_pipe_phv_out_data_104; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_105 = pipe1_io_pipe_phv_out_data_105; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_106 = pipe1_io_pipe_phv_out_data_106; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_107 = pipe1_io_pipe_phv_out_data_107; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_108 = pipe1_io_pipe_phv_out_data_108; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_109 = pipe1_io_pipe_phv_out_data_109; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_110 = pipe1_io_pipe_phv_out_data_110; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_111 = pipe1_io_pipe_phv_out_data_111; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_112 = pipe1_io_pipe_phv_out_data_112; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_113 = pipe1_io_pipe_phv_out_data_113; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_114 = pipe1_io_pipe_phv_out_data_114; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_115 = pipe1_io_pipe_phv_out_data_115; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_116 = pipe1_io_pipe_phv_out_data_116; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_117 = pipe1_io_pipe_phv_out_data_117; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_118 = pipe1_io_pipe_phv_out_data_118; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_119 = pipe1_io_pipe_phv_out_data_119; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_120 = pipe1_io_pipe_phv_out_data_120; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_121 = pipe1_io_pipe_phv_out_data_121; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_122 = pipe1_io_pipe_phv_out_data_122; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_123 = pipe1_io_pipe_phv_out_data_123; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_124 = pipe1_io_pipe_phv_out_data_124; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_125 = pipe1_io_pipe_phv_out_data_125; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_126 = pipe1_io_pipe_phv_out_data_126; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_127 = pipe1_io_pipe_phv_out_data_127; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_128 = pipe1_io_pipe_phv_out_data_128; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_129 = pipe1_io_pipe_phv_out_data_129; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_130 = pipe1_io_pipe_phv_out_data_130; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_131 = pipe1_io_pipe_phv_out_data_131; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_132 = pipe1_io_pipe_phv_out_data_132; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_133 = pipe1_io_pipe_phv_out_data_133; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_134 = pipe1_io_pipe_phv_out_data_134; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_135 = pipe1_io_pipe_phv_out_data_135; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_136 = pipe1_io_pipe_phv_out_data_136; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_137 = pipe1_io_pipe_phv_out_data_137; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_138 = pipe1_io_pipe_phv_out_data_138; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_139 = pipe1_io_pipe_phv_out_data_139; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_140 = pipe1_io_pipe_phv_out_data_140; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_141 = pipe1_io_pipe_phv_out_data_141; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_142 = pipe1_io_pipe_phv_out_data_142; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_143 = pipe1_io_pipe_phv_out_data_143; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_144 = pipe1_io_pipe_phv_out_data_144; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_145 = pipe1_io_pipe_phv_out_data_145; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_146 = pipe1_io_pipe_phv_out_data_146; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_147 = pipe1_io_pipe_phv_out_data_147; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_148 = pipe1_io_pipe_phv_out_data_148; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_149 = pipe1_io_pipe_phv_out_data_149; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_150 = pipe1_io_pipe_phv_out_data_150; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_151 = pipe1_io_pipe_phv_out_data_151; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_152 = pipe1_io_pipe_phv_out_data_152; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_153 = pipe1_io_pipe_phv_out_data_153; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_154 = pipe1_io_pipe_phv_out_data_154; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_155 = pipe1_io_pipe_phv_out_data_155; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_156 = pipe1_io_pipe_phv_out_data_156; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_157 = pipe1_io_pipe_phv_out_data_157; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_158 = pipe1_io_pipe_phv_out_data_158; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_159 = pipe1_io_pipe_phv_out_data_159; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_160 = pipe1_io_pipe_phv_out_data_160; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_161 = pipe1_io_pipe_phv_out_data_161; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_162 = pipe1_io_pipe_phv_out_data_162; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_163 = pipe1_io_pipe_phv_out_data_163; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_164 = pipe1_io_pipe_phv_out_data_164; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_165 = pipe1_io_pipe_phv_out_data_165; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_166 = pipe1_io_pipe_phv_out_data_166; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_167 = pipe1_io_pipe_phv_out_data_167; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_168 = pipe1_io_pipe_phv_out_data_168; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_169 = pipe1_io_pipe_phv_out_data_169; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_170 = pipe1_io_pipe_phv_out_data_170; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_171 = pipe1_io_pipe_phv_out_data_171; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_172 = pipe1_io_pipe_phv_out_data_172; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_173 = pipe1_io_pipe_phv_out_data_173; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_174 = pipe1_io_pipe_phv_out_data_174; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_175 = pipe1_io_pipe_phv_out_data_175; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_176 = pipe1_io_pipe_phv_out_data_176; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_177 = pipe1_io_pipe_phv_out_data_177; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_178 = pipe1_io_pipe_phv_out_data_178; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_179 = pipe1_io_pipe_phv_out_data_179; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_180 = pipe1_io_pipe_phv_out_data_180; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_181 = pipe1_io_pipe_phv_out_data_181; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_182 = pipe1_io_pipe_phv_out_data_182; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_183 = pipe1_io_pipe_phv_out_data_183; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_184 = pipe1_io_pipe_phv_out_data_184; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_185 = pipe1_io_pipe_phv_out_data_185; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_186 = pipe1_io_pipe_phv_out_data_186; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_187 = pipe1_io_pipe_phv_out_data_187; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_188 = pipe1_io_pipe_phv_out_data_188; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_189 = pipe1_io_pipe_phv_out_data_189; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_190 = pipe1_io_pipe_phv_out_data_190; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_191 = pipe1_io_pipe_phv_out_data_191; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_192 = pipe1_io_pipe_phv_out_data_192; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_193 = pipe1_io_pipe_phv_out_data_193; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_194 = pipe1_io_pipe_phv_out_data_194; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_195 = pipe1_io_pipe_phv_out_data_195; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_196 = pipe1_io_pipe_phv_out_data_196; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_197 = pipe1_io_pipe_phv_out_data_197; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_198 = pipe1_io_pipe_phv_out_data_198; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_199 = pipe1_io_pipe_phv_out_data_199; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_200 = pipe1_io_pipe_phv_out_data_200; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_201 = pipe1_io_pipe_phv_out_data_201; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_202 = pipe1_io_pipe_phv_out_data_202; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_203 = pipe1_io_pipe_phv_out_data_203; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_204 = pipe1_io_pipe_phv_out_data_204; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_205 = pipe1_io_pipe_phv_out_data_205; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_206 = pipe1_io_pipe_phv_out_data_206; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_207 = pipe1_io_pipe_phv_out_data_207; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_208 = pipe1_io_pipe_phv_out_data_208; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_209 = pipe1_io_pipe_phv_out_data_209; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_210 = pipe1_io_pipe_phv_out_data_210; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_211 = pipe1_io_pipe_phv_out_data_211; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_212 = pipe1_io_pipe_phv_out_data_212; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_213 = pipe1_io_pipe_phv_out_data_213; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_214 = pipe1_io_pipe_phv_out_data_214; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_215 = pipe1_io_pipe_phv_out_data_215; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_216 = pipe1_io_pipe_phv_out_data_216; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_217 = pipe1_io_pipe_phv_out_data_217; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_218 = pipe1_io_pipe_phv_out_data_218; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_219 = pipe1_io_pipe_phv_out_data_219; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_220 = pipe1_io_pipe_phv_out_data_220; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_221 = pipe1_io_pipe_phv_out_data_221; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_222 = pipe1_io_pipe_phv_out_data_222; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_223 = pipe1_io_pipe_phv_out_data_223; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_224 = pipe1_io_pipe_phv_out_data_224; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_225 = pipe1_io_pipe_phv_out_data_225; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_226 = pipe1_io_pipe_phv_out_data_226; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_227 = pipe1_io_pipe_phv_out_data_227; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_228 = pipe1_io_pipe_phv_out_data_228; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_229 = pipe1_io_pipe_phv_out_data_229; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_230 = pipe1_io_pipe_phv_out_data_230; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_231 = pipe1_io_pipe_phv_out_data_231; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_232 = pipe1_io_pipe_phv_out_data_232; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_233 = pipe1_io_pipe_phv_out_data_233; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_234 = pipe1_io_pipe_phv_out_data_234; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_235 = pipe1_io_pipe_phv_out_data_235; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_236 = pipe1_io_pipe_phv_out_data_236; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_237 = pipe1_io_pipe_phv_out_data_237; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_238 = pipe1_io_pipe_phv_out_data_238; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_239 = pipe1_io_pipe_phv_out_data_239; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_240 = pipe1_io_pipe_phv_out_data_240; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_241 = pipe1_io_pipe_phv_out_data_241; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_242 = pipe1_io_pipe_phv_out_data_242; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_243 = pipe1_io_pipe_phv_out_data_243; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_244 = pipe1_io_pipe_phv_out_data_244; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_245 = pipe1_io_pipe_phv_out_data_245; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_246 = pipe1_io_pipe_phv_out_data_246; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_247 = pipe1_io_pipe_phv_out_data_247; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_248 = pipe1_io_pipe_phv_out_data_248; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_249 = pipe1_io_pipe_phv_out_data_249; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_250 = pipe1_io_pipe_phv_out_data_250; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_251 = pipe1_io_pipe_phv_out_data_251; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_252 = pipe1_io_pipe_phv_out_data_252; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_253 = pipe1_io_pipe_phv_out_data_253; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_254 = pipe1_io_pipe_phv_out_data_254; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_255 = pipe1_io_pipe_phv_out_data_255; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_next_processor_id = pipe1_io_pipe_phv_out_next_processor_id; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_next_config_id = pipe1_io_pipe_phv_out_next_config_id; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_is_valid_processor = pipe1_io_pipe_phv_out_is_valid_processor; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_mod_hash_depth_mod = io_mod_en; // @[matcher_pisa.scala 342:33]
  assign pipe2_io_mod_config_id = io_mod_config_id; // @[matcher_pisa.scala 343:28]
  assign pipe2_io_mod_hash_depth = io_mod_table_mod_table_depth[3:0]; // @[matcher_pisa.scala 344:29]
  assign pipe2_io_key_in = pipe1_io_match_key; // @[matcher_pisa.scala 345:26]
  assign pipe3_clock = clock;
  assign pipe3_io_pipe_phv_in_data_0 = pipe2_io_pipe_phv_out_data_0; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_1 = pipe2_io_pipe_phv_out_data_1; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_2 = pipe2_io_pipe_phv_out_data_2; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_3 = pipe2_io_pipe_phv_out_data_3; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_4 = pipe2_io_pipe_phv_out_data_4; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_5 = pipe2_io_pipe_phv_out_data_5; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_6 = pipe2_io_pipe_phv_out_data_6; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_7 = pipe2_io_pipe_phv_out_data_7; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_8 = pipe2_io_pipe_phv_out_data_8; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_9 = pipe2_io_pipe_phv_out_data_9; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_10 = pipe2_io_pipe_phv_out_data_10; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_11 = pipe2_io_pipe_phv_out_data_11; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_12 = pipe2_io_pipe_phv_out_data_12; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_13 = pipe2_io_pipe_phv_out_data_13; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_14 = pipe2_io_pipe_phv_out_data_14; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_15 = pipe2_io_pipe_phv_out_data_15; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_16 = pipe2_io_pipe_phv_out_data_16; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_17 = pipe2_io_pipe_phv_out_data_17; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_18 = pipe2_io_pipe_phv_out_data_18; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_19 = pipe2_io_pipe_phv_out_data_19; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_20 = pipe2_io_pipe_phv_out_data_20; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_21 = pipe2_io_pipe_phv_out_data_21; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_22 = pipe2_io_pipe_phv_out_data_22; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_23 = pipe2_io_pipe_phv_out_data_23; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_24 = pipe2_io_pipe_phv_out_data_24; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_25 = pipe2_io_pipe_phv_out_data_25; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_26 = pipe2_io_pipe_phv_out_data_26; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_27 = pipe2_io_pipe_phv_out_data_27; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_28 = pipe2_io_pipe_phv_out_data_28; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_29 = pipe2_io_pipe_phv_out_data_29; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_30 = pipe2_io_pipe_phv_out_data_30; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_31 = pipe2_io_pipe_phv_out_data_31; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_32 = pipe2_io_pipe_phv_out_data_32; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_33 = pipe2_io_pipe_phv_out_data_33; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_34 = pipe2_io_pipe_phv_out_data_34; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_35 = pipe2_io_pipe_phv_out_data_35; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_36 = pipe2_io_pipe_phv_out_data_36; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_37 = pipe2_io_pipe_phv_out_data_37; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_38 = pipe2_io_pipe_phv_out_data_38; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_39 = pipe2_io_pipe_phv_out_data_39; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_40 = pipe2_io_pipe_phv_out_data_40; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_41 = pipe2_io_pipe_phv_out_data_41; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_42 = pipe2_io_pipe_phv_out_data_42; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_43 = pipe2_io_pipe_phv_out_data_43; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_44 = pipe2_io_pipe_phv_out_data_44; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_45 = pipe2_io_pipe_phv_out_data_45; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_46 = pipe2_io_pipe_phv_out_data_46; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_47 = pipe2_io_pipe_phv_out_data_47; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_48 = pipe2_io_pipe_phv_out_data_48; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_49 = pipe2_io_pipe_phv_out_data_49; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_50 = pipe2_io_pipe_phv_out_data_50; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_51 = pipe2_io_pipe_phv_out_data_51; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_52 = pipe2_io_pipe_phv_out_data_52; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_53 = pipe2_io_pipe_phv_out_data_53; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_54 = pipe2_io_pipe_phv_out_data_54; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_55 = pipe2_io_pipe_phv_out_data_55; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_56 = pipe2_io_pipe_phv_out_data_56; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_57 = pipe2_io_pipe_phv_out_data_57; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_58 = pipe2_io_pipe_phv_out_data_58; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_59 = pipe2_io_pipe_phv_out_data_59; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_60 = pipe2_io_pipe_phv_out_data_60; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_61 = pipe2_io_pipe_phv_out_data_61; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_62 = pipe2_io_pipe_phv_out_data_62; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_63 = pipe2_io_pipe_phv_out_data_63; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_64 = pipe2_io_pipe_phv_out_data_64; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_65 = pipe2_io_pipe_phv_out_data_65; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_66 = pipe2_io_pipe_phv_out_data_66; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_67 = pipe2_io_pipe_phv_out_data_67; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_68 = pipe2_io_pipe_phv_out_data_68; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_69 = pipe2_io_pipe_phv_out_data_69; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_70 = pipe2_io_pipe_phv_out_data_70; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_71 = pipe2_io_pipe_phv_out_data_71; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_72 = pipe2_io_pipe_phv_out_data_72; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_73 = pipe2_io_pipe_phv_out_data_73; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_74 = pipe2_io_pipe_phv_out_data_74; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_75 = pipe2_io_pipe_phv_out_data_75; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_76 = pipe2_io_pipe_phv_out_data_76; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_77 = pipe2_io_pipe_phv_out_data_77; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_78 = pipe2_io_pipe_phv_out_data_78; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_79 = pipe2_io_pipe_phv_out_data_79; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_80 = pipe2_io_pipe_phv_out_data_80; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_81 = pipe2_io_pipe_phv_out_data_81; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_82 = pipe2_io_pipe_phv_out_data_82; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_83 = pipe2_io_pipe_phv_out_data_83; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_84 = pipe2_io_pipe_phv_out_data_84; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_85 = pipe2_io_pipe_phv_out_data_85; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_86 = pipe2_io_pipe_phv_out_data_86; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_87 = pipe2_io_pipe_phv_out_data_87; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_88 = pipe2_io_pipe_phv_out_data_88; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_89 = pipe2_io_pipe_phv_out_data_89; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_90 = pipe2_io_pipe_phv_out_data_90; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_91 = pipe2_io_pipe_phv_out_data_91; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_92 = pipe2_io_pipe_phv_out_data_92; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_93 = pipe2_io_pipe_phv_out_data_93; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_94 = pipe2_io_pipe_phv_out_data_94; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_95 = pipe2_io_pipe_phv_out_data_95; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_96 = pipe2_io_pipe_phv_out_data_96; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_97 = pipe2_io_pipe_phv_out_data_97; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_98 = pipe2_io_pipe_phv_out_data_98; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_99 = pipe2_io_pipe_phv_out_data_99; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_100 = pipe2_io_pipe_phv_out_data_100; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_101 = pipe2_io_pipe_phv_out_data_101; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_102 = pipe2_io_pipe_phv_out_data_102; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_103 = pipe2_io_pipe_phv_out_data_103; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_104 = pipe2_io_pipe_phv_out_data_104; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_105 = pipe2_io_pipe_phv_out_data_105; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_106 = pipe2_io_pipe_phv_out_data_106; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_107 = pipe2_io_pipe_phv_out_data_107; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_108 = pipe2_io_pipe_phv_out_data_108; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_109 = pipe2_io_pipe_phv_out_data_109; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_110 = pipe2_io_pipe_phv_out_data_110; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_111 = pipe2_io_pipe_phv_out_data_111; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_112 = pipe2_io_pipe_phv_out_data_112; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_113 = pipe2_io_pipe_phv_out_data_113; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_114 = pipe2_io_pipe_phv_out_data_114; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_115 = pipe2_io_pipe_phv_out_data_115; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_116 = pipe2_io_pipe_phv_out_data_116; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_117 = pipe2_io_pipe_phv_out_data_117; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_118 = pipe2_io_pipe_phv_out_data_118; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_119 = pipe2_io_pipe_phv_out_data_119; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_120 = pipe2_io_pipe_phv_out_data_120; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_121 = pipe2_io_pipe_phv_out_data_121; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_122 = pipe2_io_pipe_phv_out_data_122; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_123 = pipe2_io_pipe_phv_out_data_123; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_124 = pipe2_io_pipe_phv_out_data_124; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_125 = pipe2_io_pipe_phv_out_data_125; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_126 = pipe2_io_pipe_phv_out_data_126; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_127 = pipe2_io_pipe_phv_out_data_127; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_128 = pipe2_io_pipe_phv_out_data_128; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_129 = pipe2_io_pipe_phv_out_data_129; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_130 = pipe2_io_pipe_phv_out_data_130; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_131 = pipe2_io_pipe_phv_out_data_131; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_132 = pipe2_io_pipe_phv_out_data_132; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_133 = pipe2_io_pipe_phv_out_data_133; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_134 = pipe2_io_pipe_phv_out_data_134; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_135 = pipe2_io_pipe_phv_out_data_135; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_136 = pipe2_io_pipe_phv_out_data_136; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_137 = pipe2_io_pipe_phv_out_data_137; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_138 = pipe2_io_pipe_phv_out_data_138; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_139 = pipe2_io_pipe_phv_out_data_139; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_140 = pipe2_io_pipe_phv_out_data_140; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_141 = pipe2_io_pipe_phv_out_data_141; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_142 = pipe2_io_pipe_phv_out_data_142; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_143 = pipe2_io_pipe_phv_out_data_143; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_144 = pipe2_io_pipe_phv_out_data_144; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_145 = pipe2_io_pipe_phv_out_data_145; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_146 = pipe2_io_pipe_phv_out_data_146; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_147 = pipe2_io_pipe_phv_out_data_147; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_148 = pipe2_io_pipe_phv_out_data_148; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_149 = pipe2_io_pipe_phv_out_data_149; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_150 = pipe2_io_pipe_phv_out_data_150; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_151 = pipe2_io_pipe_phv_out_data_151; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_152 = pipe2_io_pipe_phv_out_data_152; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_153 = pipe2_io_pipe_phv_out_data_153; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_154 = pipe2_io_pipe_phv_out_data_154; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_155 = pipe2_io_pipe_phv_out_data_155; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_156 = pipe2_io_pipe_phv_out_data_156; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_157 = pipe2_io_pipe_phv_out_data_157; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_158 = pipe2_io_pipe_phv_out_data_158; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_159 = pipe2_io_pipe_phv_out_data_159; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_160 = pipe2_io_pipe_phv_out_data_160; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_161 = pipe2_io_pipe_phv_out_data_161; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_162 = pipe2_io_pipe_phv_out_data_162; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_163 = pipe2_io_pipe_phv_out_data_163; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_164 = pipe2_io_pipe_phv_out_data_164; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_165 = pipe2_io_pipe_phv_out_data_165; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_166 = pipe2_io_pipe_phv_out_data_166; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_167 = pipe2_io_pipe_phv_out_data_167; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_168 = pipe2_io_pipe_phv_out_data_168; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_169 = pipe2_io_pipe_phv_out_data_169; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_170 = pipe2_io_pipe_phv_out_data_170; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_171 = pipe2_io_pipe_phv_out_data_171; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_172 = pipe2_io_pipe_phv_out_data_172; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_173 = pipe2_io_pipe_phv_out_data_173; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_174 = pipe2_io_pipe_phv_out_data_174; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_175 = pipe2_io_pipe_phv_out_data_175; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_176 = pipe2_io_pipe_phv_out_data_176; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_177 = pipe2_io_pipe_phv_out_data_177; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_178 = pipe2_io_pipe_phv_out_data_178; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_179 = pipe2_io_pipe_phv_out_data_179; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_180 = pipe2_io_pipe_phv_out_data_180; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_181 = pipe2_io_pipe_phv_out_data_181; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_182 = pipe2_io_pipe_phv_out_data_182; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_183 = pipe2_io_pipe_phv_out_data_183; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_184 = pipe2_io_pipe_phv_out_data_184; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_185 = pipe2_io_pipe_phv_out_data_185; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_186 = pipe2_io_pipe_phv_out_data_186; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_187 = pipe2_io_pipe_phv_out_data_187; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_188 = pipe2_io_pipe_phv_out_data_188; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_189 = pipe2_io_pipe_phv_out_data_189; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_190 = pipe2_io_pipe_phv_out_data_190; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_191 = pipe2_io_pipe_phv_out_data_191; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_192 = pipe2_io_pipe_phv_out_data_192; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_193 = pipe2_io_pipe_phv_out_data_193; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_194 = pipe2_io_pipe_phv_out_data_194; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_195 = pipe2_io_pipe_phv_out_data_195; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_196 = pipe2_io_pipe_phv_out_data_196; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_197 = pipe2_io_pipe_phv_out_data_197; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_198 = pipe2_io_pipe_phv_out_data_198; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_199 = pipe2_io_pipe_phv_out_data_199; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_200 = pipe2_io_pipe_phv_out_data_200; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_201 = pipe2_io_pipe_phv_out_data_201; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_202 = pipe2_io_pipe_phv_out_data_202; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_203 = pipe2_io_pipe_phv_out_data_203; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_204 = pipe2_io_pipe_phv_out_data_204; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_205 = pipe2_io_pipe_phv_out_data_205; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_206 = pipe2_io_pipe_phv_out_data_206; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_207 = pipe2_io_pipe_phv_out_data_207; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_208 = pipe2_io_pipe_phv_out_data_208; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_209 = pipe2_io_pipe_phv_out_data_209; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_210 = pipe2_io_pipe_phv_out_data_210; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_211 = pipe2_io_pipe_phv_out_data_211; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_212 = pipe2_io_pipe_phv_out_data_212; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_213 = pipe2_io_pipe_phv_out_data_213; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_214 = pipe2_io_pipe_phv_out_data_214; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_215 = pipe2_io_pipe_phv_out_data_215; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_216 = pipe2_io_pipe_phv_out_data_216; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_217 = pipe2_io_pipe_phv_out_data_217; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_218 = pipe2_io_pipe_phv_out_data_218; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_219 = pipe2_io_pipe_phv_out_data_219; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_220 = pipe2_io_pipe_phv_out_data_220; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_221 = pipe2_io_pipe_phv_out_data_221; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_222 = pipe2_io_pipe_phv_out_data_222; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_223 = pipe2_io_pipe_phv_out_data_223; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_224 = pipe2_io_pipe_phv_out_data_224; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_225 = pipe2_io_pipe_phv_out_data_225; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_226 = pipe2_io_pipe_phv_out_data_226; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_227 = pipe2_io_pipe_phv_out_data_227; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_228 = pipe2_io_pipe_phv_out_data_228; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_229 = pipe2_io_pipe_phv_out_data_229; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_230 = pipe2_io_pipe_phv_out_data_230; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_231 = pipe2_io_pipe_phv_out_data_231; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_232 = pipe2_io_pipe_phv_out_data_232; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_233 = pipe2_io_pipe_phv_out_data_233; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_234 = pipe2_io_pipe_phv_out_data_234; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_235 = pipe2_io_pipe_phv_out_data_235; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_236 = pipe2_io_pipe_phv_out_data_236; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_237 = pipe2_io_pipe_phv_out_data_237; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_238 = pipe2_io_pipe_phv_out_data_238; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_239 = pipe2_io_pipe_phv_out_data_239; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_240 = pipe2_io_pipe_phv_out_data_240; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_241 = pipe2_io_pipe_phv_out_data_241; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_242 = pipe2_io_pipe_phv_out_data_242; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_243 = pipe2_io_pipe_phv_out_data_243; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_244 = pipe2_io_pipe_phv_out_data_244; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_245 = pipe2_io_pipe_phv_out_data_245; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_246 = pipe2_io_pipe_phv_out_data_246; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_247 = pipe2_io_pipe_phv_out_data_247; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_248 = pipe2_io_pipe_phv_out_data_248; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_249 = pipe2_io_pipe_phv_out_data_249; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_250 = pipe2_io_pipe_phv_out_data_250; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_251 = pipe2_io_pipe_phv_out_data_251; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_252 = pipe2_io_pipe_phv_out_data_252; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_253 = pipe2_io_pipe_phv_out_data_253; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_254 = pipe2_io_pipe_phv_out_data_254; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_255 = pipe2_io_pipe_phv_out_data_255; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_next_processor_id = pipe2_io_pipe_phv_out_next_processor_id; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_next_config_id = pipe2_io_pipe_phv_out_next_config_id; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_is_valid_processor = pipe2_io_pipe_phv_out_is_valid_processor; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_table_config_0_table_depth = table_config_0_table_depth; // @[matcher_pisa.scala 348:27]
  assign pipe3_io_table_config_0_table_width = table_config_0_table_width; // @[matcher_pisa.scala 348:27]
  assign pipe3_io_table_config_1_table_depth = table_config_1_table_depth; // @[matcher_pisa.scala 348:27]
  assign pipe3_io_table_config_1_table_width = table_config_1_table_width; // @[matcher_pisa.scala 348:27]
  assign pipe3_io_key_in = pipe2_io_key_out; // @[matcher_pisa.scala 349:26]
  assign pipe3_io_addr_in = pipe2_io_hash_val; // @[matcher_pisa.scala 350:26]
  assign pipe3_io_cs_in = pipe2_io_hash_val_cs; // @[matcher_pisa.scala 351:26]
  assign pipe3_io_w_en = io_mod_w_en; // @[matcher_pisa.scala 352:26]
  assign pipe3_io_w_sram_id = io_mod_w_sram_id; // @[matcher_pisa.scala 352:26]
  assign pipe3_io_w_addr = io_mod_w_addr; // @[matcher_pisa.scala 352:26]
  assign pipe3_io_w_data = io_mod_w_data; // @[matcher_pisa.scala 352:26]
  assign pipe4_clock = clock;
  assign pipe4_io_pipe_phv_in_data_0 = pipe3_io_pipe_phv_out_data_0; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_1 = pipe3_io_pipe_phv_out_data_1; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_2 = pipe3_io_pipe_phv_out_data_2; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_3 = pipe3_io_pipe_phv_out_data_3; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_4 = pipe3_io_pipe_phv_out_data_4; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_5 = pipe3_io_pipe_phv_out_data_5; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_6 = pipe3_io_pipe_phv_out_data_6; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_7 = pipe3_io_pipe_phv_out_data_7; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_8 = pipe3_io_pipe_phv_out_data_8; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_9 = pipe3_io_pipe_phv_out_data_9; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_10 = pipe3_io_pipe_phv_out_data_10; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_11 = pipe3_io_pipe_phv_out_data_11; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_12 = pipe3_io_pipe_phv_out_data_12; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_13 = pipe3_io_pipe_phv_out_data_13; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_14 = pipe3_io_pipe_phv_out_data_14; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_15 = pipe3_io_pipe_phv_out_data_15; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_16 = pipe3_io_pipe_phv_out_data_16; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_17 = pipe3_io_pipe_phv_out_data_17; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_18 = pipe3_io_pipe_phv_out_data_18; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_19 = pipe3_io_pipe_phv_out_data_19; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_20 = pipe3_io_pipe_phv_out_data_20; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_21 = pipe3_io_pipe_phv_out_data_21; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_22 = pipe3_io_pipe_phv_out_data_22; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_23 = pipe3_io_pipe_phv_out_data_23; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_24 = pipe3_io_pipe_phv_out_data_24; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_25 = pipe3_io_pipe_phv_out_data_25; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_26 = pipe3_io_pipe_phv_out_data_26; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_27 = pipe3_io_pipe_phv_out_data_27; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_28 = pipe3_io_pipe_phv_out_data_28; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_29 = pipe3_io_pipe_phv_out_data_29; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_30 = pipe3_io_pipe_phv_out_data_30; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_31 = pipe3_io_pipe_phv_out_data_31; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_32 = pipe3_io_pipe_phv_out_data_32; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_33 = pipe3_io_pipe_phv_out_data_33; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_34 = pipe3_io_pipe_phv_out_data_34; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_35 = pipe3_io_pipe_phv_out_data_35; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_36 = pipe3_io_pipe_phv_out_data_36; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_37 = pipe3_io_pipe_phv_out_data_37; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_38 = pipe3_io_pipe_phv_out_data_38; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_39 = pipe3_io_pipe_phv_out_data_39; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_40 = pipe3_io_pipe_phv_out_data_40; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_41 = pipe3_io_pipe_phv_out_data_41; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_42 = pipe3_io_pipe_phv_out_data_42; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_43 = pipe3_io_pipe_phv_out_data_43; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_44 = pipe3_io_pipe_phv_out_data_44; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_45 = pipe3_io_pipe_phv_out_data_45; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_46 = pipe3_io_pipe_phv_out_data_46; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_47 = pipe3_io_pipe_phv_out_data_47; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_48 = pipe3_io_pipe_phv_out_data_48; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_49 = pipe3_io_pipe_phv_out_data_49; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_50 = pipe3_io_pipe_phv_out_data_50; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_51 = pipe3_io_pipe_phv_out_data_51; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_52 = pipe3_io_pipe_phv_out_data_52; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_53 = pipe3_io_pipe_phv_out_data_53; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_54 = pipe3_io_pipe_phv_out_data_54; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_55 = pipe3_io_pipe_phv_out_data_55; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_56 = pipe3_io_pipe_phv_out_data_56; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_57 = pipe3_io_pipe_phv_out_data_57; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_58 = pipe3_io_pipe_phv_out_data_58; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_59 = pipe3_io_pipe_phv_out_data_59; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_60 = pipe3_io_pipe_phv_out_data_60; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_61 = pipe3_io_pipe_phv_out_data_61; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_62 = pipe3_io_pipe_phv_out_data_62; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_63 = pipe3_io_pipe_phv_out_data_63; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_64 = pipe3_io_pipe_phv_out_data_64; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_65 = pipe3_io_pipe_phv_out_data_65; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_66 = pipe3_io_pipe_phv_out_data_66; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_67 = pipe3_io_pipe_phv_out_data_67; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_68 = pipe3_io_pipe_phv_out_data_68; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_69 = pipe3_io_pipe_phv_out_data_69; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_70 = pipe3_io_pipe_phv_out_data_70; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_71 = pipe3_io_pipe_phv_out_data_71; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_72 = pipe3_io_pipe_phv_out_data_72; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_73 = pipe3_io_pipe_phv_out_data_73; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_74 = pipe3_io_pipe_phv_out_data_74; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_75 = pipe3_io_pipe_phv_out_data_75; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_76 = pipe3_io_pipe_phv_out_data_76; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_77 = pipe3_io_pipe_phv_out_data_77; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_78 = pipe3_io_pipe_phv_out_data_78; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_79 = pipe3_io_pipe_phv_out_data_79; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_80 = pipe3_io_pipe_phv_out_data_80; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_81 = pipe3_io_pipe_phv_out_data_81; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_82 = pipe3_io_pipe_phv_out_data_82; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_83 = pipe3_io_pipe_phv_out_data_83; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_84 = pipe3_io_pipe_phv_out_data_84; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_85 = pipe3_io_pipe_phv_out_data_85; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_86 = pipe3_io_pipe_phv_out_data_86; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_87 = pipe3_io_pipe_phv_out_data_87; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_88 = pipe3_io_pipe_phv_out_data_88; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_89 = pipe3_io_pipe_phv_out_data_89; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_90 = pipe3_io_pipe_phv_out_data_90; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_91 = pipe3_io_pipe_phv_out_data_91; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_92 = pipe3_io_pipe_phv_out_data_92; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_93 = pipe3_io_pipe_phv_out_data_93; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_94 = pipe3_io_pipe_phv_out_data_94; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_95 = pipe3_io_pipe_phv_out_data_95; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_96 = pipe3_io_pipe_phv_out_data_96; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_97 = pipe3_io_pipe_phv_out_data_97; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_98 = pipe3_io_pipe_phv_out_data_98; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_99 = pipe3_io_pipe_phv_out_data_99; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_100 = pipe3_io_pipe_phv_out_data_100; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_101 = pipe3_io_pipe_phv_out_data_101; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_102 = pipe3_io_pipe_phv_out_data_102; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_103 = pipe3_io_pipe_phv_out_data_103; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_104 = pipe3_io_pipe_phv_out_data_104; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_105 = pipe3_io_pipe_phv_out_data_105; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_106 = pipe3_io_pipe_phv_out_data_106; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_107 = pipe3_io_pipe_phv_out_data_107; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_108 = pipe3_io_pipe_phv_out_data_108; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_109 = pipe3_io_pipe_phv_out_data_109; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_110 = pipe3_io_pipe_phv_out_data_110; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_111 = pipe3_io_pipe_phv_out_data_111; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_112 = pipe3_io_pipe_phv_out_data_112; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_113 = pipe3_io_pipe_phv_out_data_113; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_114 = pipe3_io_pipe_phv_out_data_114; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_115 = pipe3_io_pipe_phv_out_data_115; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_116 = pipe3_io_pipe_phv_out_data_116; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_117 = pipe3_io_pipe_phv_out_data_117; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_118 = pipe3_io_pipe_phv_out_data_118; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_119 = pipe3_io_pipe_phv_out_data_119; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_120 = pipe3_io_pipe_phv_out_data_120; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_121 = pipe3_io_pipe_phv_out_data_121; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_122 = pipe3_io_pipe_phv_out_data_122; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_123 = pipe3_io_pipe_phv_out_data_123; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_124 = pipe3_io_pipe_phv_out_data_124; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_125 = pipe3_io_pipe_phv_out_data_125; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_126 = pipe3_io_pipe_phv_out_data_126; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_127 = pipe3_io_pipe_phv_out_data_127; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_128 = pipe3_io_pipe_phv_out_data_128; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_129 = pipe3_io_pipe_phv_out_data_129; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_130 = pipe3_io_pipe_phv_out_data_130; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_131 = pipe3_io_pipe_phv_out_data_131; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_132 = pipe3_io_pipe_phv_out_data_132; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_133 = pipe3_io_pipe_phv_out_data_133; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_134 = pipe3_io_pipe_phv_out_data_134; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_135 = pipe3_io_pipe_phv_out_data_135; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_136 = pipe3_io_pipe_phv_out_data_136; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_137 = pipe3_io_pipe_phv_out_data_137; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_138 = pipe3_io_pipe_phv_out_data_138; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_139 = pipe3_io_pipe_phv_out_data_139; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_140 = pipe3_io_pipe_phv_out_data_140; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_141 = pipe3_io_pipe_phv_out_data_141; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_142 = pipe3_io_pipe_phv_out_data_142; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_143 = pipe3_io_pipe_phv_out_data_143; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_144 = pipe3_io_pipe_phv_out_data_144; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_145 = pipe3_io_pipe_phv_out_data_145; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_146 = pipe3_io_pipe_phv_out_data_146; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_147 = pipe3_io_pipe_phv_out_data_147; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_148 = pipe3_io_pipe_phv_out_data_148; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_149 = pipe3_io_pipe_phv_out_data_149; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_150 = pipe3_io_pipe_phv_out_data_150; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_151 = pipe3_io_pipe_phv_out_data_151; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_152 = pipe3_io_pipe_phv_out_data_152; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_153 = pipe3_io_pipe_phv_out_data_153; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_154 = pipe3_io_pipe_phv_out_data_154; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_155 = pipe3_io_pipe_phv_out_data_155; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_156 = pipe3_io_pipe_phv_out_data_156; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_157 = pipe3_io_pipe_phv_out_data_157; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_158 = pipe3_io_pipe_phv_out_data_158; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_159 = pipe3_io_pipe_phv_out_data_159; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_160 = pipe3_io_pipe_phv_out_data_160; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_161 = pipe3_io_pipe_phv_out_data_161; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_162 = pipe3_io_pipe_phv_out_data_162; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_163 = pipe3_io_pipe_phv_out_data_163; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_164 = pipe3_io_pipe_phv_out_data_164; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_165 = pipe3_io_pipe_phv_out_data_165; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_166 = pipe3_io_pipe_phv_out_data_166; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_167 = pipe3_io_pipe_phv_out_data_167; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_168 = pipe3_io_pipe_phv_out_data_168; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_169 = pipe3_io_pipe_phv_out_data_169; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_170 = pipe3_io_pipe_phv_out_data_170; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_171 = pipe3_io_pipe_phv_out_data_171; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_172 = pipe3_io_pipe_phv_out_data_172; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_173 = pipe3_io_pipe_phv_out_data_173; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_174 = pipe3_io_pipe_phv_out_data_174; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_175 = pipe3_io_pipe_phv_out_data_175; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_176 = pipe3_io_pipe_phv_out_data_176; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_177 = pipe3_io_pipe_phv_out_data_177; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_178 = pipe3_io_pipe_phv_out_data_178; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_179 = pipe3_io_pipe_phv_out_data_179; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_180 = pipe3_io_pipe_phv_out_data_180; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_181 = pipe3_io_pipe_phv_out_data_181; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_182 = pipe3_io_pipe_phv_out_data_182; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_183 = pipe3_io_pipe_phv_out_data_183; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_184 = pipe3_io_pipe_phv_out_data_184; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_185 = pipe3_io_pipe_phv_out_data_185; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_186 = pipe3_io_pipe_phv_out_data_186; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_187 = pipe3_io_pipe_phv_out_data_187; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_188 = pipe3_io_pipe_phv_out_data_188; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_189 = pipe3_io_pipe_phv_out_data_189; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_190 = pipe3_io_pipe_phv_out_data_190; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_191 = pipe3_io_pipe_phv_out_data_191; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_192 = pipe3_io_pipe_phv_out_data_192; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_193 = pipe3_io_pipe_phv_out_data_193; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_194 = pipe3_io_pipe_phv_out_data_194; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_195 = pipe3_io_pipe_phv_out_data_195; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_196 = pipe3_io_pipe_phv_out_data_196; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_197 = pipe3_io_pipe_phv_out_data_197; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_198 = pipe3_io_pipe_phv_out_data_198; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_199 = pipe3_io_pipe_phv_out_data_199; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_200 = pipe3_io_pipe_phv_out_data_200; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_201 = pipe3_io_pipe_phv_out_data_201; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_202 = pipe3_io_pipe_phv_out_data_202; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_203 = pipe3_io_pipe_phv_out_data_203; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_204 = pipe3_io_pipe_phv_out_data_204; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_205 = pipe3_io_pipe_phv_out_data_205; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_206 = pipe3_io_pipe_phv_out_data_206; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_207 = pipe3_io_pipe_phv_out_data_207; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_208 = pipe3_io_pipe_phv_out_data_208; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_209 = pipe3_io_pipe_phv_out_data_209; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_210 = pipe3_io_pipe_phv_out_data_210; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_211 = pipe3_io_pipe_phv_out_data_211; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_212 = pipe3_io_pipe_phv_out_data_212; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_213 = pipe3_io_pipe_phv_out_data_213; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_214 = pipe3_io_pipe_phv_out_data_214; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_215 = pipe3_io_pipe_phv_out_data_215; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_216 = pipe3_io_pipe_phv_out_data_216; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_217 = pipe3_io_pipe_phv_out_data_217; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_218 = pipe3_io_pipe_phv_out_data_218; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_219 = pipe3_io_pipe_phv_out_data_219; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_220 = pipe3_io_pipe_phv_out_data_220; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_221 = pipe3_io_pipe_phv_out_data_221; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_222 = pipe3_io_pipe_phv_out_data_222; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_223 = pipe3_io_pipe_phv_out_data_223; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_224 = pipe3_io_pipe_phv_out_data_224; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_225 = pipe3_io_pipe_phv_out_data_225; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_226 = pipe3_io_pipe_phv_out_data_226; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_227 = pipe3_io_pipe_phv_out_data_227; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_228 = pipe3_io_pipe_phv_out_data_228; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_229 = pipe3_io_pipe_phv_out_data_229; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_230 = pipe3_io_pipe_phv_out_data_230; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_231 = pipe3_io_pipe_phv_out_data_231; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_232 = pipe3_io_pipe_phv_out_data_232; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_233 = pipe3_io_pipe_phv_out_data_233; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_234 = pipe3_io_pipe_phv_out_data_234; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_235 = pipe3_io_pipe_phv_out_data_235; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_236 = pipe3_io_pipe_phv_out_data_236; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_237 = pipe3_io_pipe_phv_out_data_237; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_238 = pipe3_io_pipe_phv_out_data_238; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_239 = pipe3_io_pipe_phv_out_data_239; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_240 = pipe3_io_pipe_phv_out_data_240; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_241 = pipe3_io_pipe_phv_out_data_241; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_242 = pipe3_io_pipe_phv_out_data_242; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_243 = pipe3_io_pipe_phv_out_data_243; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_244 = pipe3_io_pipe_phv_out_data_244; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_245 = pipe3_io_pipe_phv_out_data_245; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_246 = pipe3_io_pipe_phv_out_data_246; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_247 = pipe3_io_pipe_phv_out_data_247; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_248 = pipe3_io_pipe_phv_out_data_248; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_249 = pipe3_io_pipe_phv_out_data_249; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_250 = pipe3_io_pipe_phv_out_data_250; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_251 = pipe3_io_pipe_phv_out_data_251; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_252 = pipe3_io_pipe_phv_out_data_252; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_253 = pipe3_io_pipe_phv_out_data_253; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_254 = pipe3_io_pipe_phv_out_data_254; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_255 = pipe3_io_pipe_phv_out_data_255; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_next_processor_id = pipe3_io_pipe_phv_out_next_processor_id; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_next_config_id = pipe3_io_pipe_phv_out_next_config_id; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_is_valid_processor = pipe3_io_pipe_phv_out_is_valid_processor; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_key_config_0_field_config_0 = key_config_0_field_config_0; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_0_field_config_1 = key_config_0_field_config_1; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_0_field_config_2 = key_config_0_field_config_2; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_0_field_config_3 = key_config_0_field_config_3; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_0_field_config_4 = key_config_0_field_config_4; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_0_field_config_5 = key_config_0_field_config_5; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_0_field_mask_0_0 = key_config_0_field_mask_0_0; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_0_field_mask_0_1 = key_config_0_field_mask_0_1; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_0_field_mask_0_2 = key_config_0_field_mask_0_2; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_0_field_mask_0_3 = key_config_0_field_mask_0_3; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_0_field_mask_1_0 = key_config_0_field_mask_1_0; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_0_field_mask_1_1 = key_config_0_field_mask_1_1; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_0_field_mask_1_2 = key_config_0_field_mask_1_2; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_0_field_mask_1_3 = key_config_0_field_mask_1_3; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_0_field_mask_2_0 = key_config_0_field_mask_2_0; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_0_field_mask_2_1 = key_config_0_field_mask_2_1; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_0_field_mask_2_2 = key_config_0_field_mask_2_2; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_0_field_mask_2_3 = key_config_0_field_mask_2_3; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_0_field_mask_3_0 = key_config_0_field_mask_3_0; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_0_field_mask_3_1 = key_config_0_field_mask_3_1; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_0_field_mask_3_2 = key_config_0_field_mask_3_2; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_0_field_mask_3_3 = key_config_0_field_mask_3_3; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_0_field_mask_4_0 = key_config_0_field_mask_4_0; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_0_field_mask_4_1 = key_config_0_field_mask_4_1; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_0_field_mask_4_2 = key_config_0_field_mask_4_2; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_0_field_mask_4_3 = key_config_0_field_mask_4_3; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_0_field_mask_5_0 = key_config_0_field_mask_5_0; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_0_field_mask_5_1 = key_config_0_field_mask_5_1; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_0_field_mask_5_2 = key_config_0_field_mask_5_2; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_0_field_mask_5_3 = key_config_0_field_mask_5_3; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_1_field_config_0 = key_config_1_field_config_0; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_1_field_config_1 = key_config_1_field_config_1; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_1_field_config_2 = key_config_1_field_config_2; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_1_field_config_3 = key_config_1_field_config_3; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_1_field_config_4 = key_config_1_field_config_4; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_1_field_config_5 = key_config_1_field_config_5; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_1_field_mask_0_0 = key_config_1_field_mask_0_0; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_1_field_mask_0_1 = key_config_1_field_mask_0_1; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_1_field_mask_0_2 = key_config_1_field_mask_0_2; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_1_field_mask_0_3 = key_config_1_field_mask_0_3; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_1_field_mask_1_0 = key_config_1_field_mask_1_0; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_1_field_mask_1_1 = key_config_1_field_mask_1_1; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_1_field_mask_1_2 = key_config_1_field_mask_1_2; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_1_field_mask_1_3 = key_config_1_field_mask_1_3; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_1_field_mask_2_0 = key_config_1_field_mask_2_0; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_1_field_mask_2_1 = key_config_1_field_mask_2_1; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_1_field_mask_2_2 = key_config_1_field_mask_2_2; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_1_field_mask_2_3 = key_config_1_field_mask_2_3; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_1_field_mask_3_0 = key_config_1_field_mask_3_0; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_1_field_mask_3_1 = key_config_1_field_mask_3_1; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_1_field_mask_3_2 = key_config_1_field_mask_3_2; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_1_field_mask_3_3 = key_config_1_field_mask_3_3; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_1_field_mask_4_0 = key_config_1_field_mask_4_0; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_1_field_mask_4_1 = key_config_1_field_mask_4_1; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_1_field_mask_4_2 = key_config_1_field_mask_4_2; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_1_field_mask_4_3 = key_config_1_field_mask_4_3; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_1_field_mask_5_0 = key_config_1_field_mask_5_0; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_1_field_mask_5_1 = key_config_1_field_mask_5_1; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_1_field_mask_5_2 = key_config_1_field_mask_5_2; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_1_field_mask_5_3 = key_config_1_field_mask_5_3; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_in = pipe3_io_key_out; // @[matcher_pisa.scala 355:26]
  assign pipe4_io_data_in = pipe3_io_data_out; // @[matcher_pisa.scala 356:26]
  always @(posedge clock) begin
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (~io_mod_config_id & 3'h0 == io_mod_key_mod_group_index) begin // @[matcher_pisa.scala 74:83]
          key_config_0_field_config_0 <= io_mod_key_mod_group_config; // @[matcher_pisa.scala 74:83]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (~io_mod_config_id & 3'h1 == io_mod_key_mod_group_index) begin // @[matcher_pisa.scala 74:83]
          key_config_0_field_config_1 <= io_mod_key_mod_group_config; // @[matcher_pisa.scala 74:83]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (~io_mod_config_id & 3'h2 == io_mod_key_mod_group_index) begin // @[matcher_pisa.scala 74:83]
          key_config_0_field_config_2 <= io_mod_key_mod_group_config; // @[matcher_pisa.scala 74:83]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (~io_mod_config_id & 3'h3 == io_mod_key_mod_group_index) begin // @[matcher_pisa.scala 74:83]
          key_config_0_field_config_3 <= io_mod_key_mod_group_config; // @[matcher_pisa.scala 74:83]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (~io_mod_config_id & 3'h4 == io_mod_key_mod_group_index) begin // @[matcher_pisa.scala 74:83]
          key_config_0_field_config_4 <= io_mod_key_mod_group_config; // @[matcher_pisa.scala 74:83]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (~io_mod_config_id & 3'h5 == io_mod_key_mod_group_index) begin // @[matcher_pisa.scala 74:83]
          key_config_0_field_config_5 <= io_mod_key_mod_group_config; // @[matcher_pisa.scala 74:83]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_339) begin // @[matcher_pisa.scala 76:81]
          key_config_0_field_mask_0_0 <= io_mod_key_mod_group_mask_0; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_339) begin // @[matcher_pisa.scala 76:81]
          key_config_0_field_mask_0_1 <= io_mod_key_mod_group_mask_1; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_339) begin // @[matcher_pisa.scala 76:81]
          key_config_0_field_mask_0_2 <= io_mod_key_mod_group_mask_2; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_339) begin // @[matcher_pisa.scala 76:81]
          key_config_0_field_mask_0_3 <= io_mod_key_mod_group_mask_3; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_341) begin // @[matcher_pisa.scala 76:81]
          key_config_0_field_mask_1_0 <= io_mod_key_mod_group_mask_0; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_341) begin // @[matcher_pisa.scala 76:81]
          key_config_0_field_mask_1_1 <= io_mod_key_mod_group_mask_1; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_341) begin // @[matcher_pisa.scala 76:81]
          key_config_0_field_mask_1_2 <= io_mod_key_mod_group_mask_2; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_341) begin // @[matcher_pisa.scala 76:81]
          key_config_0_field_mask_1_3 <= io_mod_key_mod_group_mask_3; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_343) begin // @[matcher_pisa.scala 76:81]
          key_config_0_field_mask_2_0 <= io_mod_key_mod_group_mask_0; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_343) begin // @[matcher_pisa.scala 76:81]
          key_config_0_field_mask_2_1 <= io_mod_key_mod_group_mask_1; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_343) begin // @[matcher_pisa.scala 76:81]
          key_config_0_field_mask_2_2 <= io_mod_key_mod_group_mask_2; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_343) begin // @[matcher_pisa.scala 76:81]
          key_config_0_field_mask_2_3 <= io_mod_key_mod_group_mask_3; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_345) begin // @[matcher_pisa.scala 76:81]
          key_config_0_field_mask_3_0 <= io_mod_key_mod_group_mask_0; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_345) begin // @[matcher_pisa.scala 76:81]
          key_config_0_field_mask_3_1 <= io_mod_key_mod_group_mask_1; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_345) begin // @[matcher_pisa.scala 76:81]
          key_config_0_field_mask_3_2 <= io_mod_key_mod_group_mask_2; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_345) begin // @[matcher_pisa.scala 76:81]
          key_config_0_field_mask_3_3 <= io_mod_key_mod_group_mask_3; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_347) begin // @[matcher_pisa.scala 76:81]
          key_config_0_field_mask_4_0 <= io_mod_key_mod_group_mask_0; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_347) begin // @[matcher_pisa.scala 76:81]
          key_config_0_field_mask_4_1 <= io_mod_key_mod_group_mask_1; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_347) begin // @[matcher_pisa.scala 76:81]
          key_config_0_field_mask_4_2 <= io_mod_key_mod_group_mask_2; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_347) begin // @[matcher_pisa.scala 76:81]
          key_config_0_field_mask_4_3 <= io_mod_key_mod_group_mask_3; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_349) begin // @[matcher_pisa.scala 76:81]
          key_config_0_field_mask_5_0 <= io_mod_key_mod_group_mask_0; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_349) begin // @[matcher_pisa.scala 76:81]
          key_config_0_field_mask_5_1 <= io_mod_key_mod_group_mask_1; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_349) begin // @[matcher_pisa.scala 76:81]
          key_config_0_field_mask_5_2 <= io_mod_key_mod_group_mask_2; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_349) begin // @[matcher_pisa.scala 76:81]
          key_config_0_field_mask_5_3 <= io_mod_key_mod_group_mask_3; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_339) begin // @[matcher_pisa.scala 75:79]
          key_config_0_field_id_0_0 <= io_mod_key_mod_group_id_0; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_339) begin // @[matcher_pisa.scala 75:79]
          key_config_0_field_id_0_1 <= io_mod_key_mod_group_id_1; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_339) begin // @[matcher_pisa.scala 75:79]
          key_config_0_field_id_0_2 <= io_mod_key_mod_group_id_2; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_339) begin // @[matcher_pisa.scala 75:79]
          key_config_0_field_id_0_3 <= io_mod_key_mod_group_id_3; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_341) begin // @[matcher_pisa.scala 75:79]
          key_config_0_field_id_1_0 <= io_mod_key_mod_group_id_0; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_341) begin // @[matcher_pisa.scala 75:79]
          key_config_0_field_id_1_1 <= io_mod_key_mod_group_id_1; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_341) begin // @[matcher_pisa.scala 75:79]
          key_config_0_field_id_1_2 <= io_mod_key_mod_group_id_2; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_341) begin // @[matcher_pisa.scala 75:79]
          key_config_0_field_id_1_3 <= io_mod_key_mod_group_id_3; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_343) begin // @[matcher_pisa.scala 75:79]
          key_config_0_field_id_2_0 <= io_mod_key_mod_group_id_0; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_343) begin // @[matcher_pisa.scala 75:79]
          key_config_0_field_id_2_1 <= io_mod_key_mod_group_id_1; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_343) begin // @[matcher_pisa.scala 75:79]
          key_config_0_field_id_2_2 <= io_mod_key_mod_group_id_2; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_343) begin // @[matcher_pisa.scala 75:79]
          key_config_0_field_id_2_3 <= io_mod_key_mod_group_id_3; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_345) begin // @[matcher_pisa.scala 75:79]
          key_config_0_field_id_3_0 <= io_mod_key_mod_group_id_0; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_345) begin // @[matcher_pisa.scala 75:79]
          key_config_0_field_id_3_1 <= io_mod_key_mod_group_id_1; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_345) begin // @[matcher_pisa.scala 75:79]
          key_config_0_field_id_3_2 <= io_mod_key_mod_group_id_2; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_345) begin // @[matcher_pisa.scala 75:79]
          key_config_0_field_id_3_3 <= io_mod_key_mod_group_id_3; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_347) begin // @[matcher_pisa.scala 75:79]
          key_config_0_field_id_4_0 <= io_mod_key_mod_group_id_0; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_347) begin // @[matcher_pisa.scala 75:79]
          key_config_0_field_id_4_1 <= io_mod_key_mod_group_id_1; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_347) begin // @[matcher_pisa.scala 75:79]
          key_config_0_field_id_4_2 <= io_mod_key_mod_group_id_2; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_347) begin // @[matcher_pisa.scala 75:79]
          key_config_0_field_id_4_3 <= io_mod_key_mod_group_id_3; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_349) begin // @[matcher_pisa.scala 75:79]
          key_config_0_field_id_5_0 <= io_mod_key_mod_group_id_0; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_349) begin // @[matcher_pisa.scala 75:79]
          key_config_0_field_id_5_1 <= io_mod_key_mod_group_id_1; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_349) begin // @[matcher_pisa.scala 75:79]
          key_config_0_field_id_5_2 <= io_mod_key_mod_group_id_2; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_349) begin // @[matcher_pisa.scala 75:79]
          key_config_0_field_id_5_3 <= io_mod_key_mod_group_id_3; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & 3'h0 == io_mod_key_mod_group_index) begin // @[matcher_pisa.scala 74:83]
          key_config_1_field_config_0 <= io_mod_key_mod_group_config; // @[matcher_pisa.scala 74:83]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & 3'h1 == io_mod_key_mod_group_index) begin // @[matcher_pisa.scala 74:83]
          key_config_1_field_config_1 <= io_mod_key_mod_group_config; // @[matcher_pisa.scala 74:83]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & 3'h2 == io_mod_key_mod_group_index) begin // @[matcher_pisa.scala 74:83]
          key_config_1_field_config_2 <= io_mod_key_mod_group_config; // @[matcher_pisa.scala 74:83]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & 3'h3 == io_mod_key_mod_group_index) begin // @[matcher_pisa.scala 74:83]
          key_config_1_field_config_3 <= io_mod_key_mod_group_config; // @[matcher_pisa.scala 74:83]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & 3'h4 == io_mod_key_mod_group_index) begin // @[matcher_pisa.scala 74:83]
          key_config_1_field_config_4 <= io_mod_key_mod_group_config; // @[matcher_pisa.scala 74:83]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & 3'h5 == io_mod_key_mod_group_index) begin // @[matcher_pisa.scala 74:83]
          key_config_1_field_config_5 <= io_mod_key_mod_group_config; // @[matcher_pisa.scala 74:83]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_339) begin // @[matcher_pisa.scala 76:81]
          key_config_1_field_mask_0_0 <= io_mod_key_mod_group_mask_0; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_339) begin // @[matcher_pisa.scala 76:81]
          key_config_1_field_mask_0_1 <= io_mod_key_mod_group_mask_1; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_339) begin // @[matcher_pisa.scala 76:81]
          key_config_1_field_mask_0_2 <= io_mod_key_mod_group_mask_2; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_339) begin // @[matcher_pisa.scala 76:81]
          key_config_1_field_mask_0_3 <= io_mod_key_mod_group_mask_3; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_341) begin // @[matcher_pisa.scala 76:81]
          key_config_1_field_mask_1_0 <= io_mod_key_mod_group_mask_0; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_341) begin // @[matcher_pisa.scala 76:81]
          key_config_1_field_mask_1_1 <= io_mod_key_mod_group_mask_1; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_341) begin // @[matcher_pisa.scala 76:81]
          key_config_1_field_mask_1_2 <= io_mod_key_mod_group_mask_2; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_341) begin // @[matcher_pisa.scala 76:81]
          key_config_1_field_mask_1_3 <= io_mod_key_mod_group_mask_3; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_343) begin // @[matcher_pisa.scala 76:81]
          key_config_1_field_mask_2_0 <= io_mod_key_mod_group_mask_0; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_343) begin // @[matcher_pisa.scala 76:81]
          key_config_1_field_mask_2_1 <= io_mod_key_mod_group_mask_1; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_343) begin // @[matcher_pisa.scala 76:81]
          key_config_1_field_mask_2_2 <= io_mod_key_mod_group_mask_2; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_343) begin // @[matcher_pisa.scala 76:81]
          key_config_1_field_mask_2_3 <= io_mod_key_mod_group_mask_3; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_345) begin // @[matcher_pisa.scala 76:81]
          key_config_1_field_mask_3_0 <= io_mod_key_mod_group_mask_0; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_345) begin // @[matcher_pisa.scala 76:81]
          key_config_1_field_mask_3_1 <= io_mod_key_mod_group_mask_1; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_345) begin // @[matcher_pisa.scala 76:81]
          key_config_1_field_mask_3_2 <= io_mod_key_mod_group_mask_2; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_345) begin // @[matcher_pisa.scala 76:81]
          key_config_1_field_mask_3_3 <= io_mod_key_mod_group_mask_3; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_347) begin // @[matcher_pisa.scala 76:81]
          key_config_1_field_mask_4_0 <= io_mod_key_mod_group_mask_0; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_347) begin // @[matcher_pisa.scala 76:81]
          key_config_1_field_mask_4_1 <= io_mod_key_mod_group_mask_1; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_347) begin // @[matcher_pisa.scala 76:81]
          key_config_1_field_mask_4_2 <= io_mod_key_mod_group_mask_2; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_347) begin // @[matcher_pisa.scala 76:81]
          key_config_1_field_mask_4_3 <= io_mod_key_mod_group_mask_3; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_349) begin // @[matcher_pisa.scala 76:81]
          key_config_1_field_mask_5_0 <= io_mod_key_mod_group_mask_0; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_349) begin // @[matcher_pisa.scala 76:81]
          key_config_1_field_mask_5_1 <= io_mod_key_mod_group_mask_1; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_349) begin // @[matcher_pisa.scala 76:81]
          key_config_1_field_mask_5_2 <= io_mod_key_mod_group_mask_2; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_349) begin // @[matcher_pisa.scala 76:81]
          key_config_1_field_mask_5_3 <= io_mod_key_mod_group_mask_3; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_339) begin // @[matcher_pisa.scala 75:79]
          key_config_1_field_id_0_0 <= io_mod_key_mod_group_id_0; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_339) begin // @[matcher_pisa.scala 75:79]
          key_config_1_field_id_0_1 <= io_mod_key_mod_group_id_1; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_339) begin // @[matcher_pisa.scala 75:79]
          key_config_1_field_id_0_2 <= io_mod_key_mod_group_id_2; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_339) begin // @[matcher_pisa.scala 75:79]
          key_config_1_field_id_0_3 <= io_mod_key_mod_group_id_3; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_341) begin // @[matcher_pisa.scala 75:79]
          key_config_1_field_id_1_0 <= io_mod_key_mod_group_id_0; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_341) begin // @[matcher_pisa.scala 75:79]
          key_config_1_field_id_1_1 <= io_mod_key_mod_group_id_1; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_341) begin // @[matcher_pisa.scala 75:79]
          key_config_1_field_id_1_2 <= io_mod_key_mod_group_id_2; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_341) begin // @[matcher_pisa.scala 75:79]
          key_config_1_field_id_1_3 <= io_mod_key_mod_group_id_3; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_343) begin // @[matcher_pisa.scala 75:79]
          key_config_1_field_id_2_0 <= io_mod_key_mod_group_id_0; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_343) begin // @[matcher_pisa.scala 75:79]
          key_config_1_field_id_2_1 <= io_mod_key_mod_group_id_1; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_343) begin // @[matcher_pisa.scala 75:79]
          key_config_1_field_id_2_2 <= io_mod_key_mod_group_id_2; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_343) begin // @[matcher_pisa.scala 75:79]
          key_config_1_field_id_2_3 <= io_mod_key_mod_group_id_3; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_345) begin // @[matcher_pisa.scala 75:79]
          key_config_1_field_id_3_0 <= io_mod_key_mod_group_id_0; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_345) begin // @[matcher_pisa.scala 75:79]
          key_config_1_field_id_3_1 <= io_mod_key_mod_group_id_1; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_345) begin // @[matcher_pisa.scala 75:79]
          key_config_1_field_id_3_2 <= io_mod_key_mod_group_id_2; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_345) begin // @[matcher_pisa.scala 75:79]
          key_config_1_field_id_3_3 <= io_mod_key_mod_group_id_3; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_347) begin // @[matcher_pisa.scala 75:79]
          key_config_1_field_id_4_0 <= io_mod_key_mod_group_id_0; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_347) begin // @[matcher_pisa.scala 75:79]
          key_config_1_field_id_4_1 <= io_mod_key_mod_group_id_1; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_347) begin // @[matcher_pisa.scala 75:79]
          key_config_1_field_id_4_2 <= io_mod_key_mod_group_id_2; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_347) begin // @[matcher_pisa.scala 75:79]
          key_config_1_field_id_4_3 <= io_mod_key_mod_group_id_3; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_349) begin // @[matcher_pisa.scala 75:79]
          key_config_1_field_id_5_0 <= io_mod_key_mod_group_id_0; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_349) begin // @[matcher_pisa.scala 75:79]
          key_config_1_field_id_5_1 <= io_mod_key_mod_group_id_1; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_349) begin // @[matcher_pisa.scala 75:79]
          key_config_1_field_id_5_2 <= io_mod_key_mod_group_id_2; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_349) begin // @[matcher_pisa.scala 75:79]
          key_config_1_field_id_5_3 <= io_mod_key_mod_group_id_3; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (~io_mod_config_id) begin // @[matcher_pisa.scala 79:40]
        table_config_0_table_depth <= io_mod_table_mod_table_depth; // @[matcher_pisa.scala 79:40]
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (~io_mod_config_id) begin // @[matcher_pisa.scala 79:40]
        table_config_0_table_width <= io_mod_table_mod_table_width; // @[matcher_pisa.scala 79:40]
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_config_id) begin // @[matcher_pisa.scala 79:40]
        table_config_1_table_depth <= io_mod_table_mod_table_depth; // @[matcher_pisa.scala 79:40]
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_config_id) begin // @[matcher_pisa.scala 79:40]
        table_config_1_table_width <= io_mod_table_mod_table_width; // @[matcher_pisa.scala 79:40]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  key_config_0_field_config_0 = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  key_config_0_field_config_1 = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  key_config_0_field_config_2 = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  key_config_0_field_config_3 = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  key_config_0_field_config_4 = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  key_config_0_field_config_5 = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  key_config_0_field_mask_0_0 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  key_config_0_field_mask_0_1 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  key_config_0_field_mask_0_2 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  key_config_0_field_mask_0_3 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  key_config_0_field_mask_1_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  key_config_0_field_mask_1_1 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  key_config_0_field_mask_1_2 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  key_config_0_field_mask_1_3 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  key_config_0_field_mask_2_0 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  key_config_0_field_mask_2_1 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  key_config_0_field_mask_2_2 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  key_config_0_field_mask_2_3 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  key_config_0_field_mask_3_0 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  key_config_0_field_mask_3_1 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  key_config_0_field_mask_3_2 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  key_config_0_field_mask_3_3 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  key_config_0_field_mask_4_0 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  key_config_0_field_mask_4_1 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  key_config_0_field_mask_4_2 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  key_config_0_field_mask_4_3 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  key_config_0_field_mask_5_0 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  key_config_0_field_mask_5_1 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  key_config_0_field_mask_5_2 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  key_config_0_field_mask_5_3 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  key_config_0_field_id_0_0 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  key_config_0_field_id_0_1 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  key_config_0_field_id_0_2 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  key_config_0_field_id_0_3 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  key_config_0_field_id_1_0 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  key_config_0_field_id_1_1 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  key_config_0_field_id_1_2 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  key_config_0_field_id_1_3 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  key_config_0_field_id_2_0 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  key_config_0_field_id_2_1 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  key_config_0_field_id_2_2 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  key_config_0_field_id_2_3 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  key_config_0_field_id_3_0 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  key_config_0_field_id_3_1 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  key_config_0_field_id_3_2 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  key_config_0_field_id_3_3 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  key_config_0_field_id_4_0 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  key_config_0_field_id_4_1 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  key_config_0_field_id_4_2 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  key_config_0_field_id_4_3 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  key_config_0_field_id_5_0 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  key_config_0_field_id_5_1 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  key_config_0_field_id_5_2 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  key_config_0_field_id_5_3 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  key_config_1_field_config_0 = _RAND_54[1:0];
  _RAND_55 = {1{`RANDOM}};
  key_config_1_field_config_1 = _RAND_55[1:0];
  _RAND_56 = {1{`RANDOM}};
  key_config_1_field_config_2 = _RAND_56[1:0];
  _RAND_57 = {1{`RANDOM}};
  key_config_1_field_config_3 = _RAND_57[1:0];
  _RAND_58 = {1{`RANDOM}};
  key_config_1_field_config_4 = _RAND_58[1:0];
  _RAND_59 = {1{`RANDOM}};
  key_config_1_field_config_5 = _RAND_59[1:0];
  _RAND_60 = {1{`RANDOM}};
  key_config_1_field_mask_0_0 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  key_config_1_field_mask_0_1 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  key_config_1_field_mask_0_2 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  key_config_1_field_mask_0_3 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  key_config_1_field_mask_1_0 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  key_config_1_field_mask_1_1 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  key_config_1_field_mask_1_2 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  key_config_1_field_mask_1_3 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  key_config_1_field_mask_2_0 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  key_config_1_field_mask_2_1 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  key_config_1_field_mask_2_2 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  key_config_1_field_mask_2_3 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  key_config_1_field_mask_3_0 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  key_config_1_field_mask_3_1 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  key_config_1_field_mask_3_2 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  key_config_1_field_mask_3_3 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  key_config_1_field_mask_4_0 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  key_config_1_field_mask_4_1 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  key_config_1_field_mask_4_2 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  key_config_1_field_mask_4_3 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  key_config_1_field_mask_5_0 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  key_config_1_field_mask_5_1 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  key_config_1_field_mask_5_2 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  key_config_1_field_mask_5_3 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  key_config_1_field_id_0_0 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  key_config_1_field_id_0_1 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  key_config_1_field_id_0_2 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  key_config_1_field_id_0_3 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  key_config_1_field_id_1_0 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  key_config_1_field_id_1_1 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  key_config_1_field_id_1_2 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  key_config_1_field_id_1_3 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  key_config_1_field_id_2_0 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  key_config_1_field_id_2_1 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  key_config_1_field_id_2_2 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  key_config_1_field_id_2_3 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  key_config_1_field_id_3_0 = _RAND_96[7:0];
  _RAND_97 = {1{`RANDOM}};
  key_config_1_field_id_3_1 = _RAND_97[7:0];
  _RAND_98 = {1{`RANDOM}};
  key_config_1_field_id_3_2 = _RAND_98[7:0];
  _RAND_99 = {1{`RANDOM}};
  key_config_1_field_id_3_3 = _RAND_99[7:0];
  _RAND_100 = {1{`RANDOM}};
  key_config_1_field_id_4_0 = _RAND_100[7:0];
  _RAND_101 = {1{`RANDOM}};
  key_config_1_field_id_4_1 = _RAND_101[7:0];
  _RAND_102 = {1{`RANDOM}};
  key_config_1_field_id_4_2 = _RAND_102[7:0];
  _RAND_103 = {1{`RANDOM}};
  key_config_1_field_id_4_3 = _RAND_103[7:0];
  _RAND_104 = {1{`RANDOM}};
  key_config_1_field_id_5_0 = _RAND_104[7:0];
  _RAND_105 = {1{`RANDOM}};
  key_config_1_field_id_5_1 = _RAND_105[7:0];
  _RAND_106 = {1{`RANDOM}};
  key_config_1_field_id_5_2 = _RAND_106[7:0];
  _RAND_107 = {1{`RANDOM}};
  key_config_1_field_id_5_3 = _RAND_107[7:0];
  _RAND_108 = {1{`RANDOM}};
  table_config_0_table_depth = _RAND_108[4:0];
  _RAND_109 = {1{`RANDOM}};
  table_config_0_table_width = _RAND_109[4:0];
  _RAND_110 = {1{`RANDOM}};
  table_config_1_table_depth = _RAND_110[4:0];
  _RAND_111 = {1{`RANDOM}};
  table_config_1_table_width = _RAND_111[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
