module PrimitiveWriteBack(
  input         clock,
  input  [7:0]  io_pipe_phv_in_data_0,
  input  [7:0]  io_pipe_phv_in_data_1,
  input  [7:0]  io_pipe_phv_in_data_2,
  input  [7:0]  io_pipe_phv_in_data_3,
  input  [7:0]  io_pipe_phv_in_data_4,
  input  [7:0]  io_pipe_phv_in_data_5,
  input  [7:0]  io_pipe_phv_in_data_6,
  input  [7:0]  io_pipe_phv_in_data_7,
  input  [7:0]  io_pipe_phv_in_data_8,
  input  [7:0]  io_pipe_phv_in_data_9,
  input  [7:0]  io_pipe_phv_in_data_10,
  input  [7:0]  io_pipe_phv_in_data_11,
  input  [7:0]  io_pipe_phv_in_data_12,
  input  [7:0]  io_pipe_phv_in_data_13,
  input  [7:0]  io_pipe_phv_in_data_14,
  input  [7:0]  io_pipe_phv_in_data_15,
  input  [7:0]  io_pipe_phv_in_data_16,
  input  [7:0]  io_pipe_phv_in_data_17,
  input  [7:0]  io_pipe_phv_in_data_18,
  input  [7:0]  io_pipe_phv_in_data_19,
  input  [7:0]  io_pipe_phv_in_data_20,
  input  [7:0]  io_pipe_phv_in_data_21,
  input  [7:0]  io_pipe_phv_in_data_22,
  input  [7:0]  io_pipe_phv_in_data_23,
  input  [7:0]  io_pipe_phv_in_data_24,
  input  [7:0]  io_pipe_phv_in_data_25,
  input  [7:0]  io_pipe_phv_in_data_26,
  input  [7:0]  io_pipe_phv_in_data_27,
  input  [7:0]  io_pipe_phv_in_data_28,
  input  [7:0]  io_pipe_phv_in_data_29,
  input  [7:0]  io_pipe_phv_in_data_30,
  input  [7:0]  io_pipe_phv_in_data_31,
  input  [7:0]  io_pipe_phv_in_data_32,
  input  [7:0]  io_pipe_phv_in_data_33,
  input  [7:0]  io_pipe_phv_in_data_34,
  input  [7:0]  io_pipe_phv_in_data_35,
  input  [7:0]  io_pipe_phv_in_data_36,
  input  [7:0]  io_pipe_phv_in_data_37,
  input  [7:0]  io_pipe_phv_in_data_38,
  input  [7:0]  io_pipe_phv_in_data_39,
  input  [7:0]  io_pipe_phv_in_data_40,
  input  [7:0]  io_pipe_phv_in_data_41,
  input  [7:0]  io_pipe_phv_in_data_42,
  input  [7:0]  io_pipe_phv_in_data_43,
  input  [7:0]  io_pipe_phv_in_data_44,
  input  [7:0]  io_pipe_phv_in_data_45,
  input  [7:0]  io_pipe_phv_in_data_46,
  input  [7:0]  io_pipe_phv_in_data_47,
  input  [7:0]  io_pipe_phv_in_data_48,
  input  [7:0]  io_pipe_phv_in_data_49,
  input  [7:0]  io_pipe_phv_in_data_50,
  input  [7:0]  io_pipe_phv_in_data_51,
  input  [7:0]  io_pipe_phv_in_data_52,
  input  [7:0]  io_pipe_phv_in_data_53,
  input  [7:0]  io_pipe_phv_in_data_54,
  input  [7:0]  io_pipe_phv_in_data_55,
  input  [7:0]  io_pipe_phv_in_data_56,
  input  [7:0]  io_pipe_phv_in_data_57,
  input  [7:0]  io_pipe_phv_in_data_58,
  input  [7:0]  io_pipe_phv_in_data_59,
  input  [7:0]  io_pipe_phv_in_data_60,
  input  [7:0]  io_pipe_phv_in_data_61,
  input  [7:0]  io_pipe_phv_in_data_62,
  input  [7:0]  io_pipe_phv_in_data_63,
  input  [7:0]  io_pipe_phv_in_data_64,
  input  [7:0]  io_pipe_phv_in_data_65,
  input  [7:0]  io_pipe_phv_in_data_66,
  input  [7:0]  io_pipe_phv_in_data_67,
  input  [7:0]  io_pipe_phv_in_data_68,
  input  [7:0]  io_pipe_phv_in_data_69,
  input  [7:0]  io_pipe_phv_in_data_70,
  input  [7:0]  io_pipe_phv_in_data_71,
  input  [7:0]  io_pipe_phv_in_data_72,
  input  [7:0]  io_pipe_phv_in_data_73,
  input  [7:0]  io_pipe_phv_in_data_74,
  input  [7:0]  io_pipe_phv_in_data_75,
  input  [7:0]  io_pipe_phv_in_data_76,
  input  [7:0]  io_pipe_phv_in_data_77,
  input  [7:0]  io_pipe_phv_in_data_78,
  input  [7:0]  io_pipe_phv_in_data_79,
  input  [7:0]  io_pipe_phv_in_data_80,
  input  [7:0]  io_pipe_phv_in_data_81,
  input  [7:0]  io_pipe_phv_in_data_82,
  input  [7:0]  io_pipe_phv_in_data_83,
  input  [7:0]  io_pipe_phv_in_data_84,
  input  [7:0]  io_pipe_phv_in_data_85,
  input  [7:0]  io_pipe_phv_in_data_86,
  input  [7:0]  io_pipe_phv_in_data_87,
  input  [7:0]  io_pipe_phv_in_data_88,
  input  [7:0]  io_pipe_phv_in_data_89,
  input  [7:0]  io_pipe_phv_in_data_90,
  input  [7:0]  io_pipe_phv_in_data_91,
  input  [7:0]  io_pipe_phv_in_data_92,
  input  [7:0]  io_pipe_phv_in_data_93,
  input  [7:0]  io_pipe_phv_in_data_94,
  input  [7:0]  io_pipe_phv_in_data_95,
  input  [7:0]  io_pipe_phv_in_data_96,
  input  [7:0]  io_pipe_phv_in_data_97,
  input  [7:0]  io_pipe_phv_in_data_98,
  input  [7:0]  io_pipe_phv_in_data_99,
  input  [7:0]  io_pipe_phv_in_data_100,
  input  [7:0]  io_pipe_phv_in_data_101,
  input  [7:0]  io_pipe_phv_in_data_102,
  input  [7:0]  io_pipe_phv_in_data_103,
  input  [7:0]  io_pipe_phv_in_data_104,
  input  [7:0]  io_pipe_phv_in_data_105,
  input  [7:0]  io_pipe_phv_in_data_106,
  input  [7:0]  io_pipe_phv_in_data_107,
  input  [7:0]  io_pipe_phv_in_data_108,
  input  [7:0]  io_pipe_phv_in_data_109,
  input  [7:0]  io_pipe_phv_in_data_110,
  input  [7:0]  io_pipe_phv_in_data_111,
  input  [7:0]  io_pipe_phv_in_data_112,
  input  [7:0]  io_pipe_phv_in_data_113,
  input  [7:0]  io_pipe_phv_in_data_114,
  input  [7:0]  io_pipe_phv_in_data_115,
  input  [7:0]  io_pipe_phv_in_data_116,
  input  [7:0]  io_pipe_phv_in_data_117,
  input  [7:0]  io_pipe_phv_in_data_118,
  input  [7:0]  io_pipe_phv_in_data_119,
  input  [7:0]  io_pipe_phv_in_data_120,
  input  [7:0]  io_pipe_phv_in_data_121,
  input  [7:0]  io_pipe_phv_in_data_122,
  input  [7:0]  io_pipe_phv_in_data_123,
  input  [7:0]  io_pipe_phv_in_data_124,
  input  [7:0]  io_pipe_phv_in_data_125,
  input  [7:0]  io_pipe_phv_in_data_126,
  input  [7:0]  io_pipe_phv_in_data_127,
  input  [7:0]  io_pipe_phv_in_data_128,
  input  [7:0]  io_pipe_phv_in_data_129,
  input  [7:0]  io_pipe_phv_in_data_130,
  input  [7:0]  io_pipe_phv_in_data_131,
  input  [7:0]  io_pipe_phv_in_data_132,
  input  [7:0]  io_pipe_phv_in_data_133,
  input  [7:0]  io_pipe_phv_in_data_134,
  input  [7:0]  io_pipe_phv_in_data_135,
  input  [7:0]  io_pipe_phv_in_data_136,
  input  [7:0]  io_pipe_phv_in_data_137,
  input  [7:0]  io_pipe_phv_in_data_138,
  input  [7:0]  io_pipe_phv_in_data_139,
  input  [7:0]  io_pipe_phv_in_data_140,
  input  [7:0]  io_pipe_phv_in_data_141,
  input  [7:0]  io_pipe_phv_in_data_142,
  input  [7:0]  io_pipe_phv_in_data_143,
  input  [7:0]  io_pipe_phv_in_data_144,
  input  [7:0]  io_pipe_phv_in_data_145,
  input  [7:0]  io_pipe_phv_in_data_146,
  input  [7:0]  io_pipe_phv_in_data_147,
  input  [7:0]  io_pipe_phv_in_data_148,
  input  [7:0]  io_pipe_phv_in_data_149,
  input  [7:0]  io_pipe_phv_in_data_150,
  input  [7:0]  io_pipe_phv_in_data_151,
  input  [7:0]  io_pipe_phv_in_data_152,
  input  [7:0]  io_pipe_phv_in_data_153,
  input  [7:0]  io_pipe_phv_in_data_154,
  input  [7:0]  io_pipe_phv_in_data_155,
  input  [7:0]  io_pipe_phv_in_data_156,
  input  [7:0]  io_pipe_phv_in_data_157,
  input  [7:0]  io_pipe_phv_in_data_158,
  input  [7:0]  io_pipe_phv_in_data_159,
  input  [7:0]  io_pipe_phv_in_data_160,
  input  [7:0]  io_pipe_phv_in_data_161,
  input  [7:0]  io_pipe_phv_in_data_162,
  input  [7:0]  io_pipe_phv_in_data_163,
  input  [7:0]  io_pipe_phv_in_data_164,
  input  [7:0]  io_pipe_phv_in_data_165,
  input  [7:0]  io_pipe_phv_in_data_166,
  input  [7:0]  io_pipe_phv_in_data_167,
  input  [7:0]  io_pipe_phv_in_data_168,
  input  [7:0]  io_pipe_phv_in_data_169,
  input  [7:0]  io_pipe_phv_in_data_170,
  input  [7:0]  io_pipe_phv_in_data_171,
  input  [7:0]  io_pipe_phv_in_data_172,
  input  [7:0]  io_pipe_phv_in_data_173,
  input  [7:0]  io_pipe_phv_in_data_174,
  input  [7:0]  io_pipe_phv_in_data_175,
  input  [7:0]  io_pipe_phv_in_data_176,
  input  [7:0]  io_pipe_phv_in_data_177,
  input  [7:0]  io_pipe_phv_in_data_178,
  input  [7:0]  io_pipe_phv_in_data_179,
  input  [7:0]  io_pipe_phv_in_data_180,
  input  [7:0]  io_pipe_phv_in_data_181,
  input  [7:0]  io_pipe_phv_in_data_182,
  input  [7:0]  io_pipe_phv_in_data_183,
  input  [7:0]  io_pipe_phv_in_data_184,
  input  [7:0]  io_pipe_phv_in_data_185,
  input  [7:0]  io_pipe_phv_in_data_186,
  input  [7:0]  io_pipe_phv_in_data_187,
  input  [7:0]  io_pipe_phv_in_data_188,
  input  [7:0]  io_pipe_phv_in_data_189,
  input  [7:0]  io_pipe_phv_in_data_190,
  input  [7:0]  io_pipe_phv_in_data_191,
  input  [7:0]  io_pipe_phv_in_data_192,
  input  [7:0]  io_pipe_phv_in_data_193,
  input  [7:0]  io_pipe_phv_in_data_194,
  input  [7:0]  io_pipe_phv_in_data_195,
  input  [7:0]  io_pipe_phv_in_data_196,
  input  [7:0]  io_pipe_phv_in_data_197,
  input  [7:0]  io_pipe_phv_in_data_198,
  input  [7:0]  io_pipe_phv_in_data_199,
  input  [7:0]  io_pipe_phv_in_data_200,
  input  [7:0]  io_pipe_phv_in_data_201,
  input  [7:0]  io_pipe_phv_in_data_202,
  input  [7:0]  io_pipe_phv_in_data_203,
  input  [7:0]  io_pipe_phv_in_data_204,
  input  [7:0]  io_pipe_phv_in_data_205,
  input  [7:0]  io_pipe_phv_in_data_206,
  input  [7:0]  io_pipe_phv_in_data_207,
  input  [7:0]  io_pipe_phv_in_data_208,
  input  [7:0]  io_pipe_phv_in_data_209,
  input  [7:0]  io_pipe_phv_in_data_210,
  input  [7:0]  io_pipe_phv_in_data_211,
  input  [7:0]  io_pipe_phv_in_data_212,
  input  [7:0]  io_pipe_phv_in_data_213,
  input  [7:0]  io_pipe_phv_in_data_214,
  input  [7:0]  io_pipe_phv_in_data_215,
  input  [7:0]  io_pipe_phv_in_data_216,
  input  [7:0]  io_pipe_phv_in_data_217,
  input  [7:0]  io_pipe_phv_in_data_218,
  input  [7:0]  io_pipe_phv_in_data_219,
  input  [7:0]  io_pipe_phv_in_data_220,
  input  [7:0]  io_pipe_phv_in_data_221,
  input  [7:0]  io_pipe_phv_in_data_222,
  input  [7:0]  io_pipe_phv_in_data_223,
  input  [7:0]  io_pipe_phv_in_data_224,
  input  [7:0]  io_pipe_phv_in_data_225,
  input  [7:0]  io_pipe_phv_in_data_226,
  input  [7:0]  io_pipe_phv_in_data_227,
  input  [7:0]  io_pipe_phv_in_data_228,
  input  [7:0]  io_pipe_phv_in_data_229,
  input  [7:0]  io_pipe_phv_in_data_230,
  input  [7:0]  io_pipe_phv_in_data_231,
  input  [7:0]  io_pipe_phv_in_data_232,
  input  [7:0]  io_pipe_phv_in_data_233,
  input  [7:0]  io_pipe_phv_in_data_234,
  input  [7:0]  io_pipe_phv_in_data_235,
  input  [7:0]  io_pipe_phv_in_data_236,
  input  [7:0]  io_pipe_phv_in_data_237,
  input  [7:0]  io_pipe_phv_in_data_238,
  input  [7:0]  io_pipe_phv_in_data_239,
  input  [7:0]  io_pipe_phv_in_data_240,
  input  [7:0]  io_pipe_phv_in_data_241,
  input  [7:0]  io_pipe_phv_in_data_242,
  input  [7:0]  io_pipe_phv_in_data_243,
  input  [7:0]  io_pipe_phv_in_data_244,
  input  [7:0]  io_pipe_phv_in_data_245,
  input  [7:0]  io_pipe_phv_in_data_246,
  input  [7:0]  io_pipe_phv_in_data_247,
  input  [7:0]  io_pipe_phv_in_data_248,
  input  [7:0]  io_pipe_phv_in_data_249,
  input  [7:0]  io_pipe_phv_in_data_250,
  input  [7:0]  io_pipe_phv_in_data_251,
  input  [7:0]  io_pipe_phv_in_data_252,
  input  [7:0]  io_pipe_phv_in_data_253,
  input  [7:0]  io_pipe_phv_in_data_254,
  input  [7:0]  io_pipe_phv_in_data_255,
  input         io_pipe_phv_in_is_valid_processor,
  output [7:0]  io_pipe_phv_out_data_0,
  output [7:0]  io_pipe_phv_out_data_1,
  output [7:0]  io_pipe_phv_out_data_2,
  output [7:0]  io_pipe_phv_out_data_3,
  output [7:0]  io_pipe_phv_out_data_4,
  output [7:0]  io_pipe_phv_out_data_5,
  output [7:0]  io_pipe_phv_out_data_6,
  output [7:0]  io_pipe_phv_out_data_7,
  output [7:0]  io_pipe_phv_out_data_8,
  output [7:0]  io_pipe_phv_out_data_9,
  output [7:0]  io_pipe_phv_out_data_10,
  output [7:0]  io_pipe_phv_out_data_11,
  output [7:0]  io_pipe_phv_out_data_12,
  output [7:0]  io_pipe_phv_out_data_13,
  output [7:0]  io_pipe_phv_out_data_14,
  output [7:0]  io_pipe_phv_out_data_15,
  output [7:0]  io_pipe_phv_out_data_16,
  output [7:0]  io_pipe_phv_out_data_17,
  output [7:0]  io_pipe_phv_out_data_18,
  output [7:0]  io_pipe_phv_out_data_19,
  output [7:0]  io_pipe_phv_out_data_20,
  output [7:0]  io_pipe_phv_out_data_21,
  output [7:0]  io_pipe_phv_out_data_22,
  output [7:0]  io_pipe_phv_out_data_23,
  output [7:0]  io_pipe_phv_out_data_24,
  output [7:0]  io_pipe_phv_out_data_25,
  output [7:0]  io_pipe_phv_out_data_26,
  output [7:0]  io_pipe_phv_out_data_27,
  output [7:0]  io_pipe_phv_out_data_28,
  output [7:0]  io_pipe_phv_out_data_29,
  output [7:0]  io_pipe_phv_out_data_30,
  output [7:0]  io_pipe_phv_out_data_31,
  output [7:0]  io_pipe_phv_out_data_32,
  output [7:0]  io_pipe_phv_out_data_33,
  output [7:0]  io_pipe_phv_out_data_34,
  output [7:0]  io_pipe_phv_out_data_35,
  output [7:0]  io_pipe_phv_out_data_36,
  output [7:0]  io_pipe_phv_out_data_37,
  output [7:0]  io_pipe_phv_out_data_38,
  output [7:0]  io_pipe_phv_out_data_39,
  output [7:0]  io_pipe_phv_out_data_40,
  output [7:0]  io_pipe_phv_out_data_41,
  output [7:0]  io_pipe_phv_out_data_42,
  output [7:0]  io_pipe_phv_out_data_43,
  output [7:0]  io_pipe_phv_out_data_44,
  output [7:0]  io_pipe_phv_out_data_45,
  output [7:0]  io_pipe_phv_out_data_46,
  output [7:0]  io_pipe_phv_out_data_47,
  output [7:0]  io_pipe_phv_out_data_48,
  output [7:0]  io_pipe_phv_out_data_49,
  output [7:0]  io_pipe_phv_out_data_50,
  output [7:0]  io_pipe_phv_out_data_51,
  output [7:0]  io_pipe_phv_out_data_52,
  output [7:0]  io_pipe_phv_out_data_53,
  output [7:0]  io_pipe_phv_out_data_54,
  output [7:0]  io_pipe_phv_out_data_55,
  output [7:0]  io_pipe_phv_out_data_56,
  output [7:0]  io_pipe_phv_out_data_57,
  output [7:0]  io_pipe_phv_out_data_58,
  output [7:0]  io_pipe_phv_out_data_59,
  output [7:0]  io_pipe_phv_out_data_60,
  output [7:0]  io_pipe_phv_out_data_61,
  output [7:0]  io_pipe_phv_out_data_62,
  output [7:0]  io_pipe_phv_out_data_63,
  output [7:0]  io_pipe_phv_out_data_64,
  output [7:0]  io_pipe_phv_out_data_65,
  output [7:0]  io_pipe_phv_out_data_66,
  output [7:0]  io_pipe_phv_out_data_67,
  output [7:0]  io_pipe_phv_out_data_68,
  output [7:0]  io_pipe_phv_out_data_69,
  output [7:0]  io_pipe_phv_out_data_70,
  output [7:0]  io_pipe_phv_out_data_71,
  output [7:0]  io_pipe_phv_out_data_72,
  output [7:0]  io_pipe_phv_out_data_73,
  output [7:0]  io_pipe_phv_out_data_74,
  output [7:0]  io_pipe_phv_out_data_75,
  output [7:0]  io_pipe_phv_out_data_76,
  output [7:0]  io_pipe_phv_out_data_77,
  output [7:0]  io_pipe_phv_out_data_78,
  output [7:0]  io_pipe_phv_out_data_79,
  output [7:0]  io_pipe_phv_out_data_80,
  output [7:0]  io_pipe_phv_out_data_81,
  output [7:0]  io_pipe_phv_out_data_82,
  output [7:0]  io_pipe_phv_out_data_83,
  output [7:0]  io_pipe_phv_out_data_84,
  output [7:0]  io_pipe_phv_out_data_85,
  output [7:0]  io_pipe_phv_out_data_86,
  output [7:0]  io_pipe_phv_out_data_87,
  output [7:0]  io_pipe_phv_out_data_88,
  output [7:0]  io_pipe_phv_out_data_89,
  output [7:0]  io_pipe_phv_out_data_90,
  output [7:0]  io_pipe_phv_out_data_91,
  output [7:0]  io_pipe_phv_out_data_92,
  output [7:0]  io_pipe_phv_out_data_93,
  output [7:0]  io_pipe_phv_out_data_94,
  output [7:0]  io_pipe_phv_out_data_95,
  output [7:0]  io_pipe_phv_out_data_96,
  output [7:0]  io_pipe_phv_out_data_97,
  output [7:0]  io_pipe_phv_out_data_98,
  output [7:0]  io_pipe_phv_out_data_99,
  output [7:0]  io_pipe_phv_out_data_100,
  output [7:0]  io_pipe_phv_out_data_101,
  output [7:0]  io_pipe_phv_out_data_102,
  output [7:0]  io_pipe_phv_out_data_103,
  output [7:0]  io_pipe_phv_out_data_104,
  output [7:0]  io_pipe_phv_out_data_105,
  output [7:0]  io_pipe_phv_out_data_106,
  output [7:0]  io_pipe_phv_out_data_107,
  output [7:0]  io_pipe_phv_out_data_108,
  output [7:0]  io_pipe_phv_out_data_109,
  output [7:0]  io_pipe_phv_out_data_110,
  output [7:0]  io_pipe_phv_out_data_111,
  output [7:0]  io_pipe_phv_out_data_112,
  output [7:0]  io_pipe_phv_out_data_113,
  output [7:0]  io_pipe_phv_out_data_114,
  output [7:0]  io_pipe_phv_out_data_115,
  output [7:0]  io_pipe_phv_out_data_116,
  output [7:0]  io_pipe_phv_out_data_117,
  output [7:0]  io_pipe_phv_out_data_118,
  output [7:0]  io_pipe_phv_out_data_119,
  output [7:0]  io_pipe_phv_out_data_120,
  output [7:0]  io_pipe_phv_out_data_121,
  output [7:0]  io_pipe_phv_out_data_122,
  output [7:0]  io_pipe_phv_out_data_123,
  output [7:0]  io_pipe_phv_out_data_124,
  output [7:0]  io_pipe_phv_out_data_125,
  output [7:0]  io_pipe_phv_out_data_126,
  output [7:0]  io_pipe_phv_out_data_127,
  output [7:0]  io_pipe_phv_out_data_128,
  output [7:0]  io_pipe_phv_out_data_129,
  output [7:0]  io_pipe_phv_out_data_130,
  output [7:0]  io_pipe_phv_out_data_131,
  output [7:0]  io_pipe_phv_out_data_132,
  output [7:0]  io_pipe_phv_out_data_133,
  output [7:0]  io_pipe_phv_out_data_134,
  output [7:0]  io_pipe_phv_out_data_135,
  output [7:0]  io_pipe_phv_out_data_136,
  output [7:0]  io_pipe_phv_out_data_137,
  output [7:0]  io_pipe_phv_out_data_138,
  output [7:0]  io_pipe_phv_out_data_139,
  output [7:0]  io_pipe_phv_out_data_140,
  output [7:0]  io_pipe_phv_out_data_141,
  output [7:0]  io_pipe_phv_out_data_142,
  output [7:0]  io_pipe_phv_out_data_143,
  output [7:0]  io_pipe_phv_out_data_144,
  output [7:0]  io_pipe_phv_out_data_145,
  output [7:0]  io_pipe_phv_out_data_146,
  output [7:0]  io_pipe_phv_out_data_147,
  output [7:0]  io_pipe_phv_out_data_148,
  output [7:0]  io_pipe_phv_out_data_149,
  output [7:0]  io_pipe_phv_out_data_150,
  output [7:0]  io_pipe_phv_out_data_151,
  output [7:0]  io_pipe_phv_out_data_152,
  output [7:0]  io_pipe_phv_out_data_153,
  output [7:0]  io_pipe_phv_out_data_154,
  output [7:0]  io_pipe_phv_out_data_155,
  output [7:0]  io_pipe_phv_out_data_156,
  output [7:0]  io_pipe_phv_out_data_157,
  output [7:0]  io_pipe_phv_out_data_158,
  output [7:0]  io_pipe_phv_out_data_159,
  output [7:0]  io_pipe_phv_out_data_160,
  output [7:0]  io_pipe_phv_out_data_161,
  output [7:0]  io_pipe_phv_out_data_162,
  output [7:0]  io_pipe_phv_out_data_163,
  output [7:0]  io_pipe_phv_out_data_164,
  output [7:0]  io_pipe_phv_out_data_165,
  output [7:0]  io_pipe_phv_out_data_166,
  output [7:0]  io_pipe_phv_out_data_167,
  output [7:0]  io_pipe_phv_out_data_168,
  output [7:0]  io_pipe_phv_out_data_169,
  output [7:0]  io_pipe_phv_out_data_170,
  output [7:0]  io_pipe_phv_out_data_171,
  output [7:0]  io_pipe_phv_out_data_172,
  output [7:0]  io_pipe_phv_out_data_173,
  output [7:0]  io_pipe_phv_out_data_174,
  output [7:0]  io_pipe_phv_out_data_175,
  output [7:0]  io_pipe_phv_out_data_176,
  output [7:0]  io_pipe_phv_out_data_177,
  output [7:0]  io_pipe_phv_out_data_178,
  output [7:0]  io_pipe_phv_out_data_179,
  output [7:0]  io_pipe_phv_out_data_180,
  output [7:0]  io_pipe_phv_out_data_181,
  output [7:0]  io_pipe_phv_out_data_182,
  output [7:0]  io_pipe_phv_out_data_183,
  output [7:0]  io_pipe_phv_out_data_184,
  output [7:0]  io_pipe_phv_out_data_185,
  output [7:0]  io_pipe_phv_out_data_186,
  output [7:0]  io_pipe_phv_out_data_187,
  output [7:0]  io_pipe_phv_out_data_188,
  output [7:0]  io_pipe_phv_out_data_189,
  output [7:0]  io_pipe_phv_out_data_190,
  output [7:0]  io_pipe_phv_out_data_191,
  output [7:0]  io_pipe_phv_out_data_192,
  output [7:0]  io_pipe_phv_out_data_193,
  output [7:0]  io_pipe_phv_out_data_194,
  output [7:0]  io_pipe_phv_out_data_195,
  output [7:0]  io_pipe_phv_out_data_196,
  output [7:0]  io_pipe_phv_out_data_197,
  output [7:0]  io_pipe_phv_out_data_198,
  output [7:0]  io_pipe_phv_out_data_199,
  output [7:0]  io_pipe_phv_out_data_200,
  output [7:0]  io_pipe_phv_out_data_201,
  output [7:0]  io_pipe_phv_out_data_202,
  output [7:0]  io_pipe_phv_out_data_203,
  output [7:0]  io_pipe_phv_out_data_204,
  output [7:0]  io_pipe_phv_out_data_205,
  output [7:0]  io_pipe_phv_out_data_206,
  output [7:0]  io_pipe_phv_out_data_207,
  output [7:0]  io_pipe_phv_out_data_208,
  output [7:0]  io_pipe_phv_out_data_209,
  output [7:0]  io_pipe_phv_out_data_210,
  output [7:0]  io_pipe_phv_out_data_211,
  output [7:0]  io_pipe_phv_out_data_212,
  output [7:0]  io_pipe_phv_out_data_213,
  output [7:0]  io_pipe_phv_out_data_214,
  output [7:0]  io_pipe_phv_out_data_215,
  output [7:0]  io_pipe_phv_out_data_216,
  output [7:0]  io_pipe_phv_out_data_217,
  output [7:0]  io_pipe_phv_out_data_218,
  output [7:0]  io_pipe_phv_out_data_219,
  output [7:0]  io_pipe_phv_out_data_220,
  output [7:0]  io_pipe_phv_out_data_221,
  output [7:0]  io_pipe_phv_out_data_222,
  output [7:0]  io_pipe_phv_out_data_223,
  output [7:0]  io_pipe_phv_out_data_224,
  output [7:0]  io_pipe_phv_out_data_225,
  output [7:0]  io_pipe_phv_out_data_226,
  output [7:0]  io_pipe_phv_out_data_227,
  output [7:0]  io_pipe_phv_out_data_228,
  output [7:0]  io_pipe_phv_out_data_229,
  output [7:0]  io_pipe_phv_out_data_230,
  output [7:0]  io_pipe_phv_out_data_231,
  output [7:0]  io_pipe_phv_out_data_232,
  output [7:0]  io_pipe_phv_out_data_233,
  output [7:0]  io_pipe_phv_out_data_234,
  output [7:0]  io_pipe_phv_out_data_235,
  output [7:0]  io_pipe_phv_out_data_236,
  output [7:0]  io_pipe_phv_out_data_237,
  output [7:0]  io_pipe_phv_out_data_238,
  output [7:0]  io_pipe_phv_out_data_239,
  output [7:0]  io_pipe_phv_out_data_240,
  output [7:0]  io_pipe_phv_out_data_241,
  output [7:0]  io_pipe_phv_out_data_242,
  output [7:0]  io_pipe_phv_out_data_243,
  output [7:0]  io_pipe_phv_out_data_244,
  output [7:0]  io_pipe_phv_out_data_245,
  output [7:0]  io_pipe_phv_out_data_246,
  output [7:0]  io_pipe_phv_out_data_247,
  output [7:0]  io_pipe_phv_out_data_248,
  output [7:0]  io_pipe_phv_out_data_249,
  output [7:0]  io_pipe_phv_out_data_250,
  output [7:0]  io_pipe_phv_out_data_251,
  output [7:0]  io_pipe_phv_out_data_252,
  output [7:0]  io_pipe_phv_out_data_253,
  output [7:0]  io_pipe_phv_out_data_254,
  output [7:0]  io_pipe_phv_out_data_255,
  input  [31:0] io_vliw_in_0,
  input  [31:0] io_vliw_in_1,
  input  [31:0] io_vliw_in_2,
  input  [31:0] io_vliw_in_3,
  input  [31:0] io_field_in_0,
  input  [31:0] io_field_in_1,
  input  [31:0] io_field_in_2,
  input  [31:0] io_field_in_3,
  input  [3:0]  io_mask_in_0,
  input  [3:0]  io_mask_in_1,
  input  [3:0]  io_mask_in_2,
  input  [3:0]  io_mask_in_3,
  input  [5:0]  io_dst_offset_in_0,
  input  [5:0]  io_dst_offset_in_1,
  input  [5:0]  io_dst_offset_in_2,
  input  [5:0]  io_dst_offset_in_3
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] phv_data_0; // @[executor.scala 448:22]
  reg [7:0] phv_data_1; // @[executor.scala 448:22]
  reg [7:0] phv_data_2; // @[executor.scala 448:22]
  reg [7:0] phv_data_3; // @[executor.scala 448:22]
  reg [7:0] phv_data_4; // @[executor.scala 448:22]
  reg [7:0] phv_data_5; // @[executor.scala 448:22]
  reg [7:0] phv_data_6; // @[executor.scala 448:22]
  reg [7:0] phv_data_7; // @[executor.scala 448:22]
  reg [7:0] phv_data_8; // @[executor.scala 448:22]
  reg [7:0] phv_data_9; // @[executor.scala 448:22]
  reg [7:0] phv_data_10; // @[executor.scala 448:22]
  reg [7:0] phv_data_11; // @[executor.scala 448:22]
  reg [7:0] phv_data_12; // @[executor.scala 448:22]
  reg [7:0] phv_data_13; // @[executor.scala 448:22]
  reg [7:0] phv_data_14; // @[executor.scala 448:22]
  reg [7:0] phv_data_15; // @[executor.scala 448:22]
  reg [7:0] phv_data_16; // @[executor.scala 448:22]
  reg [7:0] phv_data_17; // @[executor.scala 448:22]
  reg [7:0] phv_data_18; // @[executor.scala 448:22]
  reg [7:0] phv_data_19; // @[executor.scala 448:22]
  reg [7:0] phv_data_20; // @[executor.scala 448:22]
  reg [7:0] phv_data_21; // @[executor.scala 448:22]
  reg [7:0] phv_data_22; // @[executor.scala 448:22]
  reg [7:0] phv_data_23; // @[executor.scala 448:22]
  reg [7:0] phv_data_24; // @[executor.scala 448:22]
  reg [7:0] phv_data_25; // @[executor.scala 448:22]
  reg [7:0] phv_data_26; // @[executor.scala 448:22]
  reg [7:0] phv_data_27; // @[executor.scala 448:22]
  reg [7:0] phv_data_28; // @[executor.scala 448:22]
  reg [7:0] phv_data_29; // @[executor.scala 448:22]
  reg [7:0] phv_data_30; // @[executor.scala 448:22]
  reg [7:0] phv_data_31; // @[executor.scala 448:22]
  reg [7:0] phv_data_32; // @[executor.scala 448:22]
  reg [7:0] phv_data_33; // @[executor.scala 448:22]
  reg [7:0] phv_data_34; // @[executor.scala 448:22]
  reg [7:0] phv_data_35; // @[executor.scala 448:22]
  reg [7:0] phv_data_36; // @[executor.scala 448:22]
  reg [7:0] phv_data_37; // @[executor.scala 448:22]
  reg [7:0] phv_data_38; // @[executor.scala 448:22]
  reg [7:0] phv_data_39; // @[executor.scala 448:22]
  reg [7:0] phv_data_40; // @[executor.scala 448:22]
  reg [7:0] phv_data_41; // @[executor.scala 448:22]
  reg [7:0] phv_data_42; // @[executor.scala 448:22]
  reg [7:0] phv_data_43; // @[executor.scala 448:22]
  reg [7:0] phv_data_44; // @[executor.scala 448:22]
  reg [7:0] phv_data_45; // @[executor.scala 448:22]
  reg [7:0] phv_data_46; // @[executor.scala 448:22]
  reg [7:0] phv_data_47; // @[executor.scala 448:22]
  reg [7:0] phv_data_48; // @[executor.scala 448:22]
  reg [7:0] phv_data_49; // @[executor.scala 448:22]
  reg [7:0] phv_data_50; // @[executor.scala 448:22]
  reg [7:0] phv_data_51; // @[executor.scala 448:22]
  reg [7:0] phv_data_52; // @[executor.scala 448:22]
  reg [7:0] phv_data_53; // @[executor.scala 448:22]
  reg [7:0] phv_data_54; // @[executor.scala 448:22]
  reg [7:0] phv_data_55; // @[executor.scala 448:22]
  reg [7:0] phv_data_56; // @[executor.scala 448:22]
  reg [7:0] phv_data_57; // @[executor.scala 448:22]
  reg [7:0] phv_data_58; // @[executor.scala 448:22]
  reg [7:0] phv_data_59; // @[executor.scala 448:22]
  reg [7:0] phv_data_60; // @[executor.scala 448:22]
  reg [7:0] phv_data_61; // @[executor.scala 448:22]
  reg [7:0] phv_data_62; // @[executor.scala 448:22]
  reg [7:0] phv_data_63; // @[executor.scala 448:22]
  reg [7:0] phv_data_64; // @[executor.scala 448:22]
  reg [7:0] phv_data_65; // @[executor.scala 448:22]
  reg [7:0] phv_data_66; // @[executor.scala 448:22]
  reg [7:0] phv_data_67; // @[executor.scala 448:22]
  reg [7:0] phv_data_68; // @[executor.scala 448:22]
  reg [7:0] phv_data_69; // @[executor.scala 448:22]
  reg [7:0] phv_data_70; // @[executor.scala 448:22]
  reg [7:0] phv_data_71; // @[executor.scala 448:22]
  reg [7:0] phv_data_72; // @[executor.scala 448:22]
  reg [7:0] phv_data_73; // @[executor.scala 448:22]
  reg [7:0] phv_data_74; // @[executor.scala 448:22]
  reg [7:0] phv_data_75; // @[executor.scala 448:22]
  reg [7:0] phv_data_76; // @[executor.scala 448:22]
  reg [7:0] phv_data_77; // @[executor.scala 448:22]
  reg [7:0] phv_data_78; // @[executor.scala 448:22]
  reg [7:0] phv_data_79; // @[executor.scala 448:22]
  reg [7:0] phv_data_80; // @[executor.scala 448:22]
  reg [7:0] phv_data_81; // @[executor.scala 448:22]
  reg [7:0] phv_data_82; // @[executor.scala 448:22]
  reg [7:0] phv_data_83; // @[executor.scala 448:22]
  reg [7:0] phv_data_84; // @[executor.scala 448:22]
  reg [7:0] phv_data_85; // @[executor.scala 448:22]
  reg [7:0] phv_data_86; // @[executor.scala 448:22]
  reg [7:0] phv_data_87; // @[executor.scala 448:22]
  reg [7:0] phv_data_88; // @[executor.scala 448:22]
  reg [7:0] phv_data_89; // @[executor.scala 448:22]
  reg [7:0] phv_data_90; // @[executor.scala 448:22]
  reg [7:0] phv_data_91; // @[executor.scala 448:22]
  reg [7:0] phv_data_92; // @[executor.scala 448:22]
  reg [7:0] phv_data_93; // @[executor.scala 448:22]
  reg [7:0] phv_data_94; // @[executor.scala 448:22]
  reg [7:0] phv_data_95; // @[executor.scala 448:22]
  reg [7:0] phv_data_96; // @[executor.scala 448:22]
  reg [7:0] phv_data_97; // @[executor.scala 448:22]
  reg [7:0] phv_data_98; // @[executor.scala 448:22]
  reg [7:0] phv_data_99; // @[executor.scala 448:22]
  reg [7:0] phv_data_100; // @[executor.scala 448:22]
  reg [7:0] phv_data_101; // @[executor.scala 448:22]
  reg [7:0] phv_data_102; // @[executor.scala 448:22]
  reg [7:0] phv_data_103; // @[executor.scala 448:22]
  reg [7:0] phv_data_104; // @[executor.scala 448:22]
  reg [7:0] phv_data_105; // @[executor.scala 448:22]
  reg [7:0] phv_data_106; // @[executor.scala 448:22]
  reg [7:0] phv_data_107; // @[executor.scala 448:22]
  reg [7:0] phv_data_108; // @[executor.scala 448:22]
  reg [7:0] phv_data_109; // @[executor.scala 448:22]
  reg [7:0] phv_data_110; // @[executor.scala 448:22]
  reg [7:0] phv_data_111; // @[executor.scala 448:22]
  reg [7:0] phv_data_112; // @[executor.scala 448:22]
  reg [7:0] phv_data_113; // @[executor.scala 448:22]
  reg [7:0] phv_data_114; // @[executor.scala 448:22]
  reg [7:0] phv_data_115; // @[executor.scala 448:22]
  reg [7:0] phv_data_116; // @[executor.scala 448:22]
  reg [7:0] phv_data_117; // @[executor.scala 448:22]
  reg [7:0] phv_data_118; // @[executor.scala 448:22]
  reg [7:0] phv_data_119; // @[executor.scala 448:22]
  reg [7:0] phv_data_120; // @[executor.scala 448:22]
  reg [7:0] phv_data_121; // @[executor.scala 448:22]
  reg [7:0] phv_data_122; // @[executor.scala 448:22]
  reg [7:0] phv_data_123; // @[executor.scala 448:22]
  reg [7:0] phv_data_124; // @[executor.scala 448:22]
  reg [7:0] phv_data_125; // @[executor.scala 448:22]
  reg [7:0] phv_data_126; // @[executor.scala 448:22]
  reg [7:0] phv_data_127; // @[executor.scala 448:22]
  reg [7:0] phv_data_128; // @[executor.scala 448:22]
  reg [7:0] phv_data_129; // @[executor.scala 448:22]
  reg [7:0] phv_data_130; // @[executor.scala 448:22]
  reg [7:0] phv_data_131; // @[executor.scala 448:22]
  reg [7:0] phv_data_132; // @[executor.scala 448:22]
  reg [7:0] phv_data_133; // @[executor.scala 448:22]
  reg [7:0] phv_data_134; // @[executor.scala 448:22]
  reg [7:0] phv_data_135; // @[executor.scala 448:22]
  reg [7:0] phv_data_136; // @[executor.scala 448:22]
  reg [7:0] phv_data_137; // @[executor.scala 448:22]
  reg [7:0] phv_data_138; // @[executor.scala 448:22]
  reg [7:0] phv_data_139; // @[executor.scala 448:22]
  reg [7:0] phv_data_140; // @[executor.scala 448:22]
  reg [7:0] phv_data_141; // @[executor.scala 448:22]
  reg [7:0] phv_data_142; // @[executor.scala 448:22]
  reg [7:0] phv_data_143; // @[executor.scala 448:22]
  reg [7:0] phv_data_144; // @[executor.scala 448:22]
  reg [7:0] phv_data_145; // @[executor.scala 448:22]
  reg [7:0] phv_data_146; // @[executor.scala 448:22]
  reg [7:0] phv_data_147; // @[executor.scala 448:22]
  reg [7:0] phv_data_148; // @[executor.scala 448:22]
  reg [7:0] phv_data_149; // @[executor.scala 448:22]
  reg [7:0] phv_data_150; // @[executor.scala 448:22]
  reg [7:0] phv_data_151; // @[executor.scala 448:22]
  reg [7:0] phv_data_152; // @[executor.scala 448:22]
  reg [7:0] phv_data_153; // @[executor.scala 448:22]
  reg [7:0] phv_data_154; // @[executor.scala 448:22]
  reg [7:0] phv_data_155; // @[executor.scala 448:22]
  reg [7:0] phv_data_156; // @[executor.scala 448:22]
  reg [7:0] phv_data_157; // @[executor.scala 448:22]
  reg [7:0] phv_data_158; // @[executor.scala 448:22]
  reg [7:0] phv_data_159; // @[executor.scala 448:22]
  reg [7:0] phv_data_160; // @[executor.scala 448:22]
  reg [7:0] phv_data_161; // @[executor.scala 448:22]
  reg [7:0] phv_data_162; // @[executor.scala 448:22]
  reg [7:0] phv_data_163; // @[executor.scala 448:22]
  reg [7:0] phv_data_164; // @[executor.scala 448:22]
  reg [7:0] phv_data_165; // @[executor.scala 448:22]
  reg [7:0] phv_data_166; // @[executor.scala 448:22]
  reg [7:0] phv_data_167; // @[executor.scala 448:22]
  reg [7:0] phv_data_168; // @[executor.scala 448:22]
  reg [7:0] phv_data_169; // @[executor.scala 448:22]
  reg [7:0] phv_data_170; // @[executor.scala 448:22]
  reg [7:0] phv_data_171; // @[executor.scala 448:22]
  reg [7:0] phv_data_172; // @[executor.scala 448:22]
  reg [7:0] phv_data_173; // @[executor.scala 448:22]
  reg [7:0] phv_data_174; // @[executor.scala 448:22]
  reg [7:0] phv_data_175; // @[executor.scala 448:22]
  reg [7:0] phv_data_176; // @[executor.scala 448:22]
  reg [7:0] phv_data_177; // @[executor.scala 448:22]
  reg [7:0] phv_data_178; // @[executor.scala 448:22]
  reg [7:0] phv_data_179; // @[executor.scala 448:22]
  reg [7:0] phv_data_180; // @[executor.scala 448:22]
  reg [7:0] phv_data_181; // @[executor.scala 448:22]
  reg [7:0] phv_data_182; // @[executor.scala 448:22]
  reg [7:0] phv_data_183; // @[executor.scala 448:22]
  reg [7:0] phv_data_184; // @[executor.scala 448:22]
  reg [7:0] phv_data_185; // @[executor.scala 448:22]
  reg [7:0] phv_data_186; // @[executor.scala 448:22]
  reg [7:0] phv_data_187; // @[executor.scala 448:22]
  reg [7:0] phv_data_188; // @[executor.scala 448:22]
  reg [7:0] phv_data_189; // @[executor.scala 448:22]
  reg [7:0] phv_data_190; // @[executor.scala 448:22]
  reg [7:0] phv_data_191; // @[executor.scala 448:22]
  reg [7:0] phv_data_192; // @[executor.scala 448:22]
  reg [7:0] phv_data_193; // @[executor.scala 448:22]
  reg [7:0] phv_data_194; // @[executor.scala 448:22]
  reg [7:0] phv_data_195; // @[executor.scala 448:22]
  reg [7:0] phv_data_196; // @[executor.scala 448:22]
  reg [7:0] phv_data_197; // @[executor.scala 448:22]
  reg [7:0] phv_data_198; // @[executor.scala 448:22]
  reg [7:0] phv_data_199; // @[executor.scala 448:22]
  reg [7:0] phv_data_200; // @[executor.scala 448:22]
  reg [7:0] phv_data_201; // @[executor.scala 448:22]
  reg [7:0] phv_data_202; // @[executor.scala 448:22]
  reg [7:0] phv_data_203; // @[executor.scala 448:22]
  reg [7:0] phv_data_204; // @[executor.scala 448:22]
  reg [7:0] phv_data_205; // @[executor.scala 448:22]
  reg [7:0] phv_data_206; // @[executor.scala 448:22]
  reg [7:0] phv_data_207; // @[executor.scala 448:22]
  reg [7:0] phv_data_208; // @[executor.scala 448:22]
  reg [7:0] phv_data_209; // @[executor.scala 448:22]
  reg [7:0] phv_data_210; // @[executor.scala 448:22]
  reg [7:0] phv_data_211; // @[executor.scala 448:22]
  reg [7:0] phv_data_212; // @[executor.scala 448:22]
  reg [7:0] phv_data_213; // @[executor.scala 448:22]
  reg [7:0] phv_data_214; // @[executor.scala 448:22]
  reg [7:0] phv_data_215; // @[executor.scala 448:22]
  reg [7:0] phv_data_216; // @[executor.scala 448:22]
  reg [7:0] phv_data_217; // @[executor.scala 448:22]
  reg [7:0] phv_data_218; // @[executor.scala 448:22]
  reg [7:0] phv_data_219; // @[executor.scala 448:22]
  reg [7:0] phv_data_220; // @[executor.scala 448:22]
  reg [7:0] phv_data_221; // @[executor.scala 448:22]
  reg [7:0] phv_data_222; // @[executor.scala 448:22]
  reg [7:0] phv_data_223; // @[executor.scala 448:22]
  reg [7:0] phv_data_224; // @[executor.scala 448:22]
  reg [7:0] phv_data_225; // @[executor.scala 448:22]
  reg [7:0] phv_data_226; // @[executor.scala 448:22]
  reg [7:0] phv_data_227; // @[executor.scala 448:22]
  reg [7:0] phv_data_228; // @[executor.scala 448:22]
  reg [7:0] phv_data_229; // @[executor.scala 448:22]
  reg [7:0] phv_data_230; // @[executor.scala 448:22]
  reg [7:0] phv_data_231; // @[executor.scala 448:22]
  reg [7:0] phv_data_232; // @[executor.scala 448:22]
  reg [7:0] phv_data_233; // @[executor.scala 448:22]
  reg [7:0] phv_data_234; // @[executor.scala 448:22]
  reg [7:0] phv_data_235; // @[executor.scala 448:22]
  reg [7:0] phv_data_236; // @[executor.scala 448:22]
  reg [7:0] phv_data_237; // @[executor.scala 448:22]
  reg [7:0] phv_data_238; // @[executor.scala 448:22]
  reg [7:0] phv_data_239; // @[executor.scala 448:22]
  reg [7:0] phv_data_240; // @[executor.scala 448:22]
  reg [7:0] phv_data_241; // @[executor.scala 448:22]
  reg [7:0] phv_data_242; // @[executor.scala 448:22]
  reg [7:0] phv_data_243; // @[executor.scala 448:22]
  reg [7:0] phv_data_244; // @[executor.scala 448:22]
  reg [7:0] phv_data_245; // @[executor.scala 448:22]
  reg [7:0] phv_data_246; // @[executor.scala 448:22]
  reg [7:0] phv_data_247; // @[executor.scala 448:22]
  reg [7:0] phv_data_248; // @[executor.scala 448:22]
  reg [7:0] phv_data_249; // @[executor.scala 448:22]
  reg [7:0] phv_data_250; // @[executor.scala 448:22]
  reg [7:0] phv_data_251; // @[executor.scala 448:22]
  reg [7:0] phv_data_252; // @[executor.scala 448:22]
  reg [7:0] phv_data_253; // @[executor.scala 448:22]
  reg [7:0] phv_data_254; // @[executor.scala 448:22]
  reg [7:0] phv_data_255; // @[executor.scala 448:22]
  reg  phv_is_valid_processor; // @[executor.scala 448:22]
  reg [31:0] vliw_0; // @[executor.scala 452:23]
  reg [31:0] vliw_1; // @[executor.scala 452:23]
  reg [31:0] vliw_2; // @[executor.scala 452:23]
  reg [31:0] vliw_3; // @[executor.scala 452:23]
  reg [31:0] field_0; // @[executor.scala 454:24]
  reg [31:0] field_1; // @[executor.scala 454:24]
  reg [31:0] field_2; // @[executor.scala 454:24]
  reg [31:0] field_3; // @[executor.scala 454:24]
  reg [3:0] mask_0; // @[executor.scala 456:23]
  reg [3:0] mask_1; // @[executor.scala 456:23]
  reg [3:0] mask_2; // @[executor.scala 456:23]
  reg [3:0] mask_3; // @[executor.scala 456:23]
  reg [5:0] dst_offset_0; // @[executor.scala 458:29]
  reg [5:0] dst_offset_1; // @[executor.scala 458:29]
  reg [5:0] dst_offset_2; // @[executor.scala 458:29]
  reg [5:0] dst_offset_3; // @[executor.scala 458:29]
  wire [3:0] opcode = vliw_0[31:28]; // @[primitive.scala 9:44]
  wire [7:0] _GEN_4362 = {{2'd0}, dst_offset_0}; // @[executor.scala 473:49]
  wire [7:0] byte_ = field_0[7:0]; // @[executor.scala 475:56]
  wire [7:0] _GEN_0 = mask_0[0] ? byte_ : phv_data_3; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] byte_1 = field_0[15:8]; // @[executor.scala 475:56]
  wire [7:0] _GEN_1 = mask_0[1] ? byte_1 : phv_data_2; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] byte_2 = field_0[23:16]; // @[executor.scala 475:56]
  wire [7:0] _GEN_2 = mask_0[2] ? byte_2 : phv_data_1; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] byte_3 = field_0[31:24]; // @[executor.scala 475:56]
  wire [7:0] _GEN_3 = mask_0[3] ? byte_3 : phv_data_0; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_4 = _GEN_4362 == 8'h0 ? _GEN_0 : phv_data_3; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_5 = _GEN_4362 == 8'h0 ? _GEN_1 : phv_data_2; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_6 = _GEN_4362 == 8'h0 ? _GEN_2 : phv_data_1; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_7 = _GEN_4362 == 8'h0 ? _GEN_3 : phv_data_0; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_8 = mask_0[0] ? byte_ : phv_data_7; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_9 = mask_0[1] ? byte_1 : phv_data_6; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_10 = mask_0[2] ? byte_2 : phv_data_5; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_11 = mask_0[3] ? byte_3 : phv_data_4; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_12 = _GEN_4362 == 8'h1 ? _GEN_8 : phv_data_7; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_13 = _GEN_4362 == 8'h1 ? _GEN_9 : phv_data_6; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_14 = _GEN_4362 == 8'h1 ? _GEN_10 : phv_data_5; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_15 = _GEN_4362 == 8'h1 ? _GEN_11 : phv_data_4; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_16 = mask_0[0] ? byte_ : phv_data_11; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_17 = mask_0[1] ? byte_1 : phv_data_10; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_18 = mask_0[2] ? byte_2 : phv_data_9; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_19 = mask_0[3] ? byte_3 : phv_data_8; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_20 = _GEN_4362 == 8'h2 ? _GEN_16 : phv_data_11; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_21 = _GEN_4362 == 8'h2 ? _GEN_17 : phv_data_10; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_22 = _GEN_4362 == 8'h2 ? _GEN_18 : phv_data_9; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_23 = _GEN_4362 == 8'h2 ? _GEN_19 : phv_data_8; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_24 = mask_0[0] ? byte_ : phv_data_15; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_25 = mask_0[1] ? byte_1 : phv_data_14; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_26 = mask_0[2] ? byte_2 : phv_data_13; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_27 = mask_0[3] ? byte_3 : phv_data_12; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_28 = _GEN_4362 == 8'h3 ? _GEN_24 : phv_data_15; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_29 = _GEN_4362 == 8'h3 ? _GEN_25 : phv_data_14; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_30 = _GEN_4362 == 8'h3 ? _GEN_26 : phv_data_13; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_31 = _GEN_4362 == 8'h3 ? _GEN_27 : phv_data_12; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_32 = mask_0[0] ? byte_ : phv_data_19; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_33 = mask_0[1] ? byte_1 : phv_data_18; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_34 = mask_0[2] ? byte_2 : phv_data_17; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_35 = mask_0[3] ? byte_3 : phv_data_16; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_36 = _GEN_4362 == 8'h4 ? _GEN_32 : phv_data_19; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_37 = _GEN_4362 == 8'h4 ? _GEN_33 : phv_data_18; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_38 = _GEN_4362 == 8'h4 ? _GEN_34 : phv_data_17; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_39 = _GEN_4362 == 8'h4 ? _GEN_35 : phv_data_16; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_40 = mask_0[0] ? byte_ : phv_data_23; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_41 = mask_0[1] ? byte_1 : phv_data_22; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_42 = mask_0[2] ? byte_2 : phv_data_21; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_43 = mask_0[3] ? byte_3 : phv_data_20; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_44 = _GEN_4362 == 8'h5 ? _GEN_40 : phv_data_23; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_45 = _GEN_4362 == 8'h5 ? _GEN_41 : phv_data_22; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_46 = _GEN_4362 == 8'h5 ? _GEN_42 : phv_data_21; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_47 = _GEN_4362 == 8'h5 ? _GEN_43 : phv_data_20; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_48 = mask_0[0] ? byte_ : phv_data_27; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_49 = mask_0[1] ? byte_1 : phv_data_26; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_50 = mask_0[2] ? byte_2 : phv_data_25; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_51 = mask_0[3] ? byte_3 : phv_data_24; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_52 = _GEN_4362 == 8'h6 ? _GEN_48 : phv_data_27; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_53 = _GEN_4362 == 8'h6 ? _GEN_49 : phv_data_26; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_54 = _GEN_4362 == 8'h6 ? _GEN_50 : phv_data_25; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_55 = _GEN_4362 == 8'h6 ? _GEN_51 : phv_data_24; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_56 = mask_0[0] ? byte_ : phv_data_31; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_57 = mask_0[1] ? byte_1 : phv_data_30; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_58 = mask_0[2] ? byte_2 : phv_data_29; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_59 = mask_0[3] ? byte_3 : phv_data_28; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_60 = _GEN_4362 == 8'h7 ? _GEN_56 : phv_data_31; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_61 = _GEN_4362 == 8'h7 ? _GEN_57 : phv_data_30; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_62 = _GEN_4362 == 8'h7 ? _GEN_58 : phv_data_29; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_63 = _GEN_4362 == 8'h7 ? _GEN_59 : phv_data_28; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_64 = mask_0[0] ? byte_ : phv_data_35; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_65 = mask_0[1] ? byte_1 : phv_data_34; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_66 = mask_0[2] ? byte_2 : phv_data_33; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_67 = mask_0[3] ? byte_3 : phv_data_32; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_68 = _GEN_4362 == 8'h8 ? _GEN_64 : phv_data_35; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_69 = _GEN_4362 == 8'h8 ? _GEN_65 : phv_data_34; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_70 = _GEN_4362 == 8'h8 ? _GEN_66 : phv_data_33; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_71 = _GEN_4362 == 8'h8 ? _GEN_67 : phv_data_32; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_72 = mask_0[0] ? byte_ : phv_data_39; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_73 = mask_0[1] ? byte_1 : phv_data_38; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_74 = mask_0[2] ? byte_2 : phv_data_37; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_75 = mask_0[3] ? byte_3 : phv_data_36; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_76 = _GEN_4362 == 8'h9 ? _GEN_72 : phv_data_39; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_77 = _GEN_4362 == 8'h9 ? _GEN_73 : phv_data_38; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_78 = _GEN_4362 == 8'h9 ? _GEN_74 : phv_data_37; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_79 = _GEN_4362 == 8'h9 ? _GEN_75 : phv_data_36; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_80 = mask_0[0] ? byte_ : phv_data_43; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_81 = mask_0[1] ? byte_1 : phv_data_42; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_82 = mask_0[2] ? byte_2 : phv_data_41; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_83 = mask_0[3] ? byte_3 : phv_data_40; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_84 = _GEN_4362 == 8'ha ? _GEN_80 : phv_data_43; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_85 = _GEN_4362 == 8'ha ? _GEN_81 : phv_data_42; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_86 = _GEN_4362 == 8'ha ? _GEN_82 : phv_data_41; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_87 = _GEN_4362 == 8'ha ? _GEN_83 : phv_data_40; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_88 = mask_0[0] ? byte_ : phv_data_47; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_89 = mask_0[1] ? byte_1 : phv_data_46; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_90 = mask_0[2] ? byte_2 : phv_data_45; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_91 = mask_0[3] ? byte_3 : phv_data_44; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_92 = _GEN_4362 == 8'hb ? _GEN_88 : phv_data_47; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_93 = _GEN_4362 == 8'hb ? _GEN_89 : phv_data_46; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_94 = _GEN_4362 == 8'hb ? _GEN_90 : phv_data_45; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_95 = _GEN_4362 == 8'hb ? _GEN_91 : phv_data_44; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_96 = mask_0[0] ? byte_ : phv_data_51; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_97 = mask_0[1] ? byte_1 : phv_data_50; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_98 = mask_0[2] ? byte_2 : phv_data_49; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_99 = mask_0[3] ? byte_3 : phv_data_48; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_100 = _GEN_4362 == 8'hc ? _GEN_96 : phv_data_51; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_101 = _GEN_4362 == 8'hc ? _GEN_97 : phv_data_50; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_102 = _GEN_4362 == 8'hc ? _GEN_98 : phv_data_49; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_103 = _GEN_4362 == 8'hc ? _GEN_99 : phv_data_48; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_104 = mask_0[0] ? byte_ : phv_data_55; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_105 = mask_0[1] ? byte_1 : phv_data_54; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_106 = mask_0[2] ? byte_2 : phv_data_53; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_107 = mask_0[3] ? byte_3 : phv_data_52; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_108 = _GEN_4362 == 8'hd ? _GEN_104 : phv_data_55; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_109 = _GEN_4362 == 8'hd ? _GEN_105 : phv_data_54; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_110 = _GEN_4362 == 8'hd ? _GEN_106 : phv_data_53; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_111 = _GEN_4362 == 8'hd ? _GEN_107 : phv_data_52; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_112 = mask_0[0] ? byte_ : phv_data_59; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_113 = mask_0[1] ? byte_1 : phv_data_58; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_114 = mask_0[2] ? byte_2 : phv_data_57; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_115 = mask_0[3] ? byte_3 : phv_data_56; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_116 = _GEN_4362 == 8'he ? _GEN_112 : phv_data_59; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_117 = _GEN_4362 == 8'he ? _GEN_113 : phv_data_58; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_118 = _GEN_4362 == 8'he ? _GEN_114 : phv_data_57; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_119 = _GEN_4362 == 8'he ? _GEN_115 : phv_data_56; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_120 = mask_0[0] ? byte_ : phv_data_63; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_121 = mask_0[1] ? byte_1 : phv_data_62; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_122 = mask_0[2] ? byte_2 : phv_data_61; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_123 = mask_0[3] ? byte_3 : phv_data_60; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_124 = _GEN_4362 == 8'hf ? _GEN_120 : phv_data_63; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_125 = _GEN_4362 == 8'hf ? _GEN_121 : phv_data_62; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_126 = _GEN_4362 == 8'hf ? _GEN_122 : phv_data_61; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_127 = _GEN_4362 == 8'hf ? _GEN_123 : phv_data_60; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_128 = mask_0[0] ? byte_ : phv_data_67; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_129 = mask_0[1] ? byte_1 : phv_data_66; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_130 = mask_0[2] ? byte_2 : phv_data_65; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_131 = mask_0[3] ? byte_3 : phv_data_64; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_132 = _GEN_4362 == 8'h10 ? _GEN_128 : phv_data_67; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_133 = _GEN_4362 == 8'h10 ? _GEN_129 : phv_data_66; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_134 = _GEN_4362 == 8'h10 ? _GEN_130 : phv_data_65; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_135 = _GEN_4362 == 8'h10 ? _GEN_131 : phv_data_64; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_136 = mask_0[0] ? byte_ : phv_data_71; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_137 = mask_0[1] ? byte_1 : phv_data_70; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_138 = mask_0[2] ? byte_2 : phv_data_69; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_139 = mask_0[3] ? byte_3 : phv_data_68; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_140 = _GEN_4362 == 8'h11 ? _GEN_136 : phv_data_71; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_141 = _GEN_4362 == 8'h11 ? _GEN_137 : phv_data_70; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_142 = _GEN_4362 == 8'h11 ? _GEN_138 : phv_data_69; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_143 = _GEN_4362 == 8'h11 ? _GEN_139 : phv_data_68; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_144 = mask_0[0] ? byte_ : phv_data_75; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_145 = mask_0[1] ? byte_1 : phv_data_74; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_146 = mask_0[2] ? byte_2 : phv_data_73; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_147 = mask_0[3] ? byte_3 : phv_data_72; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_148 = _GEN_4362 == 8'h12 ? _GEN_144 : phv_data_75; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_149 = _GEN_4362 == 8'h12 ? _GEN_145 : phv_data_74; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_150 = _GEN_4362 == 8'h12 ? _GEN_146 : phv_data_73; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_151 = _GEN_4362 == 8'h12 ? _GEN_147 : phv_data_72; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_152 = mask_0[0] ? byte_ : phv_data_79; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_153 = mask_0[1] ? byte_1 : phv_data_78; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_154 = mask_0[2] ? byte_2 : phv_data_77; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_155 = mask_0[3] ? byte_3 : phv_data_76; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_156 = _GEN_4362 == 8'h13 ? _GEN_152 : phv_data_79; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_157 = _GEN_4362 == 8'h13 ? _GEN_153 : phv_data_78; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_158 = _GEN_4362 == 8'h13 ? _GEN_154 : phv_data_77; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_159 = _GEN_4362 == 8'h13 ? _GEN_155 : phv_data_76; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_160 = mask_0[0] ? byte_ : phv_data_83; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_161 = mask_0[1] ? byte_1 : phv_data_82; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_162 = mask_0[2] ? byte_2 : phv_data_81; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_163 = mask_0[3] ? byte_3 : phv_data_80; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_164 = _GEN_4362 == 8'h14 ? _GEN_160 : phv_data_83; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_165 = _GEN_4362 == 8'h14 ? _GEN_161 : phv_data_82; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_166 = _GEN_4362 == 8'h14 ? _GEN_162 : phv_data_81; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_167 = _GEN_4362 == 8'h14 ? _GEN_163 : phv_data_80; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_168 = mask_0[0] ? byte_ : phv_data_87; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_169 = mask_0[1] ? byte_1 : phv_data_86; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_170 = mask_0[2] ? byte_2 : phv_data_85; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_171 = mask_0[3] ? byte_3 : phv_data_84; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_172 = _GEN_4362 == 8'h15 ? _GEN_168 : phv_data_87; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_173 = _GEN_4362 == 8'h15 ? _GEN_169 : phv_data_86; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_174 = _GEN_4362 == 8'h15 ? _GEN_170 : phv_data_85; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_175 = _GEN_4362 == 8'h15 ? _GEN_171 : phv_data_84; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_176 = mask_0[0] ? byte_ : phv_data_91; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_177 = mask_0[1] ? byte_1 : phv_data_90; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_178 = mask_0[2] ? byte_2 : phv_data_89; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_179 = mask_0[3] ? byte_3 : phv_data_88; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_180 = _GEN_4362 == 8'h16 ? _GEN_176 : phv_data_91; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_181 = _GEN_4362 == 8'h16 ? _GEN_177 : phv_data_90; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_182 = _GEN_4362 == 8'h16 ? _GEN_178 : phv_data_89; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_183 = _GEN_4362 == 8'h16 ? _GEN_179 : phv_data_88; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_184 = mask_0[0] ? byte_ : phv_data_95; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_185 = mask_0[1] ? byte_1 : phv_data_94; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_186 = mask_0[2] ? byte_2 : phv_data_93; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_187 = mask_0[3] ? byte_3 : phv_data_92; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_188 = _GEN_4362 == 8'h17 ? _GEN_184 : phv_data_95; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_189 = _GEN_4362 == 8'h17 ? _GEN_185 : phv_data_94; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_190 = _GEN_4362 == 8'h17 ? _GEN_186 : phv_data_93; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_191 = _GEN_4362 == 8'h17 ? _GEN_187 : phv_data_92; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_192 = mask_0[0] ? byte_ : phv_data_99; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_193 = mask_0[1] ? byte_1 : phv_data_98; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_194 = mask_0[2] ? byte_2 : phv_data_97; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_195 = mask_0[3] ? byte_3 : phv_data_96; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_196 = _GEN_4362 == 8'h18 ? _GEN_192 : phv_data_99; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_197 = _GEN_4362 == 8'h18 ? _GEN_193 : phv_data_98; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_198 = _GEN_4362 == 8'h18 ? _GEN_194 : phv_data_97; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_199 = _GEN_4362 == 8'h18 ? _GEN_195 : phv_data_96; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_200 = mask_0[0] ? byte_ : phv_data_103; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_201 = mask_0[1] ? byte_1 : phv_data_102; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_202 = mask_0[2] ? byte_2 : phv_data_101; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_203 = mask_0[3] ? byte_3 : phv_data_100; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_204 = _GEN_4362 == 8'h19 ? _GEN_200 : phv_data_103; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_205 = _GEN_4362 == 8'h19 ? _GEN_201 : phv_data_102; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_206 = _GEN_4362 == 8'h19 ? _GEN_202 : phv_data_101; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_207 = _GEN_4362 == 8'h19 ? _GEN_203 : phv_data_100; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_208 = mask_0[0] ? byte_ : phv_data_107; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_209 = mask_0[1] ? byte_1 : phv_data_106; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_210 = mask_0[2] ? byte_2 : phv_data_105; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_211 = mask_0[3] ? byte_3 : phv_data_104; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_212 = _GEN_4362 == 8'h1a ? _GEN_208 : phv_data_107; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_213 = _GEN_4362 == 8'h1a ? _GEN_209 : phv_data_106; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_214 = _GEN_4362 == 8'h1a ? _GEN_210 : phv_data_105; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_215 = _GEN_4362 == 8'h1a ? _GEN_211 : phv_data_104; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_216 = mask_0[0] ? byte_ : phv_data_111; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_217 = mask_0[1] ? byte_1 : phv_data_110; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_218 = mask_0[2] ? byte_2 : phv_data_109; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_219 = mask_0[3] ? byte_3 : phv_data_108; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_220 = _GEN_4362 == 8'h1b ? _GEN_216 : phv_data_111; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_221 = _GEN_4362 == 8'h1b ? _GEN_217 : phv_data_110; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_222 = _GEN_4362 == 8'h1b ? _GEN_218 : phv_data_109; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_223 = _GEN_4362 == 8'h1b ? _GEN_219 : phv_data_108; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_224 = mask_0[0] ? byte_ : phv_data_115; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_225 = mask_0[1] ? byte_1 : phv_data_114; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_226 = mask_0[2] ? byte_2 : phv_data_113; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_227 = mask_0[3] ? byte_3 : phv_data_112; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_228 = _GEN_4362 == 8'h1c ? _GEN_224 : phv_data_115; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_229 = _GEN_4362 == 8'h1c ? _GEN_225 : phv_data_114; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_230 = _GEN_4362 == 8'h1c ? _GEN_226 : phv_data_113; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_231 = _GEN_4362 == 8'h1c ? _GEN_227 : phv_data_112; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_232 = mask_0[0] ? byte_ : phv_data_119; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_233 = mask_0[1] ? byte_1 : phv_data_118; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_234 = mask_0[2] ? byte_2 : phv_data_117; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_235 = mask_0[3] ? byte_3 : phv_data_116; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_236 = _GEN_4362 == 8'h1d ? _GEN_232 : phv_data_119; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_237 = _GEN_4362 == 8'h1d ? _GEN_233 : phv_data_118; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_238 = _GEN_4362 == 8'h1d ? _GEN_234 : phv_data_117; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_239 = _GEN_4362 == 8'h1d ? _GEN_235 : phv_data_116; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_240 = mask_0[0] ? byte_ : phv_data_123; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_241 = mask_0[1] ? byte_1 : phv_data_122; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_242 = mask_0[2] ? byte_2 : phv_data_121; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_243 = mask_0[3] ? byte_3 : phv_data_120; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_244 = _GEN_4362 == 8'h1e ? _GEN_240 : phv_data_123; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_245 = _GEN_4362 == 8'h1e ? _GEN_241 : phv_data_122; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_246 = _GEN_4362 == 8'h1e ? _GEN_242 : phv_data_121; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_247 = _GEN_4362 == 8'h1e ? _GEN_243 : phv_data_120; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_248 = mask_0[0] ? byte_ : phv_data_127; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_249 = mask_0[1] ? byte_1 : phv_data_126; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_250 = mask_0[2] ? byte_2 : phv_data_125; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_251 = mask_0[3] ? byte_3 : phv_data_124; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_252 = _GEN_4362 == 8'h1f ? _GEN_248 : phv_data_127; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_253 = _GEN_4362 == 8'h1f ? _GEN_249 : phv_data_126; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_254 = _GEN_4362 == 8'h1f ? _GEN_250 : phv_data_125; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_255 = _GEN_4362 == 8'h1f ? _GEN_251 : phv_data_124; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_256 = mask_0[0] ? byte_ : phv_data_131; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_257 = mask_0[1] ? byte_1 : phv_data_130; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_258 = mask_0[2] ? byte_2 : phv_data_129; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_259 = mask_0[3] ? byte_3 : phv_data_128; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_260 = _GEN_4362 == 8'h20 ? _GEN_256 : phv_data_131; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_261 = _GEN_4362 == 8'h20 ? _GEN_257 : phv_data_130; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_262 = _GEN_4362 == 8'h20 ? _GEN_258 : phv_data_129; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_263 = _GEN_4362 == 8'h20 ? _GEN_259 : phv_data_128; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_264 = mask_0[0] ? byte_ : phv_data_135; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_265 = mask_0[1] ? byte_1 : phv_data_134; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_266 = mask_0[2] ? byte_2 : phv_data_133; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_267 = mask_0[3] ? byte_3 : phv_data_132; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_268 = _GEN_4362 == 8'h21 ? _GEN_264 : phv_data_135; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_269 = _GEN_4362 == 8'h21 ? _GEN_265 : phv_data_134; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_270 = _GEN_4362 == 8'h21 ? _GEN_266 : phv_data_133; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_271 = _GEN_4362 == 8'h21 ? _GEN_267 : phv_data_132; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_272 = mask_0[0] ? byte_ : phv_data_139; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_273 = mask_0[1] ? byte_1 : phv_data_138; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_274 = mask_0[2] ? byte_2 : phv_data_137; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_275 = mask_0[3] ? byte_3 : phv_data_136; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_276 = _GEN_4362 == 8'h22 ? _GEN_272 : phv_data_139; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_277 = _GEN_4362 == 8'h22 ? _GEN_273 : phv_data_138; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_278 = _GEN_4362 == 8'h22 ? _GEN_274 : phv_data_137; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_279 = _GEN_4362 == 8'h22 ? _GEN_275 : phv_data_136; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_280 = mask_0[0] ? byte_ : phv_data_143; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_281 = mask_0[1] ? byte_1 : phv_data_142; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_282 = mask_0[2] ? byte_2 : phv_data_141; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_283 = mask_0[3] ? byte_3 : phv_data_140; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_284 = _GEN_4362 == 8'h23 ? _GEN_280 : phv_data_143; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_285 = _GEN_4362 == 8'h23 ? _GEN_281 : phv_data_142; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_286 = _GEN_4362 == 8'h23 ? _GEN_282 : phv_data_141; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_287 = _GEN_4362 == 8'h23 ? _GEN_283 : phv_data_140; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_288 = mask_0[0] ? byte_ : phv_data_147; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_289 = mask_0[1] ? byte_1 : phv_data_146; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_290 = mask_0[2] ? byte_2 : phv_data_145; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_291 = mask_0[3] ? byte_3 : phv_data_144; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_292 = _GEN_4362 == 8'h24 ? _GEN_288 : phv_data_147; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_293 = _GEN_4362 == 8'h24 ? _GEN_289 : phv_data_146; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_294 = _GEN_4362 == 8'h24 ? _GEN_290 : phv_data_145; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_295 = _GEN_4362 == 8'h24 ? _GEN_291 : phv_data_144; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_296 = mask_0[0] ? byte_ : phv_data_151; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_297 = mask_0[1] ? byte_1 : phv_data_150; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_298 = mask_0[2] ? byte_2 : phv_data_149; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_299 = mask_0[3] ? byte_3 : phv_data_148; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_300 = _GEN_4362 == 8'h25 ? _GEN_296 : phv_data_151; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_301 = _GEN_4362 == 8'h25 ? _GEN_297 : phv_data_150; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_302 = _GEN_4362 == 8'h25 ? _GEN_298 : phv_data_149; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_303 = _GEN_4362 == 8'h25 ? _GEN_299 : phv_data_148; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_304 = mask_0[0] ? byte_ : phv_data_155; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_305 = mask_0[1] ? byte_1 : phv_data_154; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_306 = mask_0[2] ? byte_2 : phv_data_153; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_307 = mask_0[3] ? byte_3 : phv_data_152; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_308 = _GEN_4362 == 8'h26 ? _GEN_304 : phv_data_155; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_309 = _GEN_4362 == 8'h26 ? _GEN_305 : phv_data_154; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_310 = _GEN_4362 == 8'h26 ? _GEN_306 : phv_data_153; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_311 = _GEN_4362 == 8'h26 ? _GEN_307 : phv_data_152; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_312 = mask_0[0] ? byte_ : phv_data_159; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_313 = mask_0[1] ? byte_1 : phv_data_158; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_314 = mask_0[2] ? byte_2 : phv_data_157; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_315 = mask_0[3] ? byte_3 : phv_data_156; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_316 = _GEN_4362 == 8'h27 ? _GEN_312 : phv_data_159; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_317 = _GEN_4362 == 8'h27 ? _GEN_313 : phv_data_158; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_318 = _GEN_4362 == 8'h27 ? _GEN_314 : phv_data_157; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_319 = _GEN_4362 == 8'h27 ? _GEN_315 : phv_data_156; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_320 = mask_0[0] ? byte_ : phv_data_163; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_321 = mask_0[1] ? byte_1 : phv_data_162; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_322 = mask_0[2] ? byte_2 : phv_data_161; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_323 = mask_0[3] ? byte_3 : phv_data_160; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_324 = _GEN_4362 == 8'h28 ? _GEN_320 : phv_data_163; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_325 = _GEN_4362 == 8'h28 ? _GEN_321 : phv_data_162; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_326 = _GEN_4362 == 8'h28 ? _GEN_322 : phv_data_161; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_327 = _GEN_4362 == 8'h28 ? _GEN_323 : phv_data_160; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_328 = mask_0[0] ? byte_ : phv_data_167; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_329 = mask_0[1] ? byte_1 : phv_data_166; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_330 = mask_0[2] ? byte_2 : phv_data_165; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_331 = mask_0[3] ? byte_3 : phv_data_164; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_332 = _GEN_4362 == 8'h29 ? _GEN_328 : phv_data_167; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_333 = _GEN_4362 == 8'h29 ? _GEN_329 : phv_data_166; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_334 = _GEN_4362 == 8'h29 ? _GEN_330 : phv_data_165; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_335 = _GEN_4362 == 8'h29 ? _GEN_331 : phv_data_164; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_336 = mask_0[0] ? byte_ : phv_data_171; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_337 = mask_0[1] ? byte_1 : phv_data_170; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_338 = mask_0[2] ? byte_2 : phv_data_169; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_339 = mask_0[3] ? byte_3 : phv_data_168; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_340 = _GEN_4362 == 8'h2a ? _GEN_336 : phv_data_171; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_341 = _GEN_4362 == 8'h2a ? _GEN_337 : phv_data_170; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_342 = _GEN_4362 == 8'h2a ? _GEN_338 : phv_data_169; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_343 = _GEN_4362 == 8'h2a ? _GEN_339 : phv_data_168; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_344 = mask_0[0] ? byte_ : phv_data_175; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_345 = mask_0[1] ? byte_1 : phv_data_174; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_346 = mask_0[2] ? byte_2 : phv_data_173; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_347 = mask_0[3] ? byte_3 : phv_data_172; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_348 = _GEN_4362 == 8'h2b ? _GEN_344 : phv_data_175; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_349 = _GEN_4362 == 8'h2b ? _GEN_345 : phv_data_174; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_350 = _GEN_4362 == 8'h2b ? _GEN_346 : phv_data_173; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_351 = _GEN_4362 == 8'h2b ? _GEN_347 : phv_data_172; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_352 = mask_0[0] ? byte_ : phv_data_179; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_353 = mask_0[1] ? byte_1 : phv_data_178; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_354 = mask_0[2] ? byte_2 : phv_data_177; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_355 = mask_0[3] ? byte_3 : phv_data_176; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_356 = _GEN_4362 == 8'h2c ? _GEN_352 : phv_data_179; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_357 = _GEN_4362 == 8'h2c ? _GEN_353 : phv_data_178; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_358 = _GEN_4362 == 8'h2c ? _GEN_354 : phv_data_177; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_359 = _GEN_4362 == 8'h2c ? _GEN_355 : phv_data_176; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_360 = mask_0[0] ? byte_ : phv_data_183; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_361 = mask_0[1] ? byte_1 : phv_data_182; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_362 = mask_0[2] ? byte_2 : phv_data_181; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_363 = mask_0[3] ? byte_3 : phv_data_180; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_364 = _GEN_4362 == 8'h2d ? _GEN_360 : phv_data_183; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_365 = _GEN_4362 == 8'h2d ? _GEN_361 : phv_data_182; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_366 = _GEN_4362 == 8'h2d ? _GEN_362 : phv_data_181; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_367 = _GEN_4362 == 8'h2d ? _GEN_363 : phv_data_180; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_368 = mask_0[0] ? byte_ : phv_data_187; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_369 = mask_0[1] ? byte_1 : phv_data_186; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_370 = mask_0[2] ? byte_2 : phv_data_185; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_371 = mask_0[3] ? byte_3 : phv_data_184; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_372 = _GEN_4362 == 8'h2e ? _GEN_368 : phv_data_187; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_373 = _GEN_4362 == 8'h2e ? _GEN_369 : phv_data_186; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_374 = _GEN_4362 == 8'h2e ? _GEN_370 : phv_data_185; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_375 = _GEN_4362 == 8'h2e ? _GEN_371 : phv_data_184; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_376 = mask_0[0] ? byte_ : phv_data_191; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_377 = mask_0[1] ? byte_1 : phv_data_190; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_378 = mask_0[2] ? byte_2 : phv_data_189; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_379 = mask_0[3] ? byte_3 : phv_data_188; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_380 = _GEN_4362 == 8'h2f ? _GEN_376 : phv_data_191; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_381 = _GEN_4362 == 8'h2f ? _GEN_377 : phv_data_190; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_382 = _GEN_4362 == 8'h2f ? _GEN_378 : phv_data_189; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_383 = _GEN_4362 == 8'h2f ? _GEN_379 : phv_data_188; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_384 = mask_0[0] ? byte_ : phv_data_195; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_385 = mask_0[1] ? byte_1 : phv_data_194; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_386 = mask_0[2] ? byte_2 : phv_data_193; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_387 = mask_0[3] ? byte_3 : phv_data_192; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_388 = _GEN_4362 == 8'h30 ? _GEN_384 : phv_data_195; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_389 = _GEN_4362 == 8'h30 ? _GEN_385 : phv_data_194; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_390 = _GEN_4362 == 8'h30 ? _GEN_386 : phv_data_193; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_391 = _GEN_4362 == 8'h30 ? _GEN_387 : phv_data_192; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_392 = mask_0[0] ? byte_ : phv_data_199; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_393 = mask_0[1] ? byte_1 : phv_data_198; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_394 = mask_0[2] ? byte_2 : phv_data_197; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_395 = mask_0[3] ? byte_3 : phv_data_196; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_396 = _GEN_4362 == 8'h31 ? _GEN_392 : phv_data_199; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_397 = _GEN_4362 == 8'h31 ? _GEN_393 : phv_data_198; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_398 = _GEN_4362 == 8'h31 ? _GEN_394 : phv_data_197; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_399 = _GEN_4362 == 8'h31 ? _GEN_395 : phv_data_196; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_400 = mask_0[0] ? byte_ : phv_data_203; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_401 = mask_0[1] ? byte_1 : phv_data_202; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_402 = mask_0[2] ? byte_2 : phv_data_201; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_403 = mask_0[3] ? byte_3 : phv_data_200; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_404 = _GEN_4362 == 8'h32 ? _GEN_400 : phv_data_203; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_405 = _GEN_4362 == 8'h32 ? _GEN_401 : phv_data_202; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_406 = _GEN_4362 == 8'h32 ? _GEN_402 : phv_data_201; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_407 = _GEN_4362 == 8'h32 ? _GEN_403 : phv_data_200; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_408 = mask_0[0] ? byte_ : phv_data_207; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_409 = mask_0[1] ? byte_1 : phv_data_206; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_410 = mask_0[2] ? byte_2 : phv_data_205; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_411 = mask_0[3] ? byte_3 : phv_data_204; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_412 = _GEN_4362 == 8'h33 ? _GEN_408 : phv_data_207; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_413 = _GEN_4362 == 8'h33 ? _GEN_409 : phv_data_206; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_414 = _GEN_4362 == 8'h33 ? _GEN_410 : phv_data_205; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_415 = _GEN_4362 == 8'h33 ? _GEN_411 : phv_data_204; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_416 = mask_0[0] ? byte_ : phv_data_211; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_417 = mask_0[1] ? byte_1 : phv_data_210; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_418 = mask_0[2] ? byte_2 : phv_data_209; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_419 = mask_0[3] ? byte_3 : phv_data_208; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_420 = _GEN_4362 == 8'h34 ? _GEN_416 : phv_data_211; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_421 = _GEN_4362 == 8'h34 ? _GEN_417 : phv_data_210; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_422 = _GEN_4362 == 8'h34 ? _GEN_418 : phv_data_209; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_423 = _GEN_4362 == 8'h34 ? _GEN_419 : phv_data_208; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_424 = mask_0[0] ? byte_ : phv_data_215; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_425 = mask_0[1] ? byte_1 : phv_data_214; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_426 = mask_0[2] ? byte_2 : phv_data_213; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_427 = mask_0[3] ? byte_3 : phv_data_212; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_428 = _GEN_4362 == 8'h35 ? _GEN_424 : phv_data_215; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_429 = _GEN_4362 == 8'h35 ? _GEN_425 : phv_data_214; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_430 = _GEN_4362 == 8'h35 ? _GEN_426 : phv_data_213; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_431 = _GEN_4362 == 8'h35 ? _GEN_427 : phv_data_212; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_432 = mask_0[0] ? byte_ : phv_data_219; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_433 = mask_0[1] ? byte_1 : phv_data_218; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_434 = mask_0[2] ? byte_2 : phv_data_217; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_435 = mask_0[3] ? byte_3 : phv_data_216; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_436 = _GEN_4362 == 8'h36 ? _GEN_432 : phv_data_219; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_437 = _GEN_4362 == 8'h36 ? _GEN_433 : phv_data_218; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_438 = _GEN_4362 == 8'h36 ? _GEN_434 : phv_data_217; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_439 = _GEN_4362 == 8'h36 ? _GEN_435 : phv_data_216; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_440 = mask_0[0] ? byte_ : phv_data_223; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_441 = mask_0[1] ? byte_1 : phv_data_222; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_442 = mask_0[2] ? byte_2 : phv_data_221; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_443 = mask_0[3] ? byte_3 : phv_data_220; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_444 = _GEN_4362 == 8'h37 ? _GEN_440 : phv_data_223; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_445 = _GEN_4362 == 8'h37 ? _GEN_441 : phv_data_222; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_446 = _GEN_4362 == 8'h37 ? _GEN_442 : phv_data_221; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_447 = _GEN_4362 == 8'h37 ? _GEN_443 : phv_data_220; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_448 = mask_0[0] ? byte_ : phv_data_227; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_449 = mask_0[1] ? byte_1 : phv_data_226; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_450 = mask_0[2] ? byte_2 : phv_data_225; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_451 = mask_0[3] ? byte_3 : phv_data_224; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_452 = _GEN_4362 == 8'h38 ? _GEN_448 : phv_data_227; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_453 = _GEN_4362 == 8'h38 ? _GEN_449 : phv_data_226; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_454 = _GEN_4362 == 8'h38 ? _GEN_450 : phv_data_225; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_455 = _GEN_4362 == 8'h38 ? _GEN_451 : phv_data_224; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_456 = mask_0[0] ? byte_ : phv_data_231; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_457 = mask_0[1] ? byte_1 : phv_data_230; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_458 = mask_0[2] ? byte_2 : phv_data_229; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_459 = mask_0[3] ? byte_3 : phv_data_228; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_460 = _GEN_4362 == 8'h39 ? _GEN_456 : phv_data_231; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_461 = _GEN_4362 == 8'h39 ? _GEN_457 : phv_data_230; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_462 = _GEN_4362 == 8'h39 ? _GEN_458 : phv_data_229; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_463 = _GEN_4362 == 8'h39 ? _GEN_459 : phv_data_228; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_464 = mask_0[0] ? byte_ : phv_data_235; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_465 = mask_0[1] ? byte_1 : phv_data_234; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_466 = mask_0[2] ? byte_2 : phv_data_233; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_467 = mask_0[3] ? byte_3 : phv_data_232; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_468 = _GEN_4362 == 8'h3a ? _GEN_464 : phv_data_235; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_469 = _GEN_4362 == 8'h3a ? _GEN_465 : phv_data_234; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_470 = _GEN_4362 == 8'h3a ? _GEN_466 : phv_data_233; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_471 = _GEN_4362 == 8'h3a ? _GEN_467 : phv_data_232; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_472 = mask_0[0] ? byte_ : phv_data_239; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_473 = mask_0[1] ? byte_1 : phv_data_238; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_474 = mask_0[2] ? byte_2 : phv_data_237; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_475 = mask_0[3] ? byte_3 : phv_data_236; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_476 = _GEN_4362 == 8'h3b ? _GEN_472 : phv_data_239; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_477 = _GEN_4362 == 8'h3b ? _GEN_473 : phv_data_238; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_478 = _GEN_4362 == 8'h3b ? _GEN_474 : phv_data_237; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_479 = _GEN_4362 == 8'h3b ? _GEN_475 : phv_data_236; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_480 = mask_0[0] ? byte_ : phv_data_243; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_481 = mask_0[1] ? byte_1 : phv_data_242; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_482 = mask_0[2] ? byte_2 : phv_data_241; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_483 = mask_0[3] ? byte_3 : phv_data_240; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_484 = _GEN_4362 == 8'h3c ? _GEN_480 : phv_data_243; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_485 = _GEN_4362 == 8'h3c ? _GEN_481 : phv_data_242; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_486 = _GEN_4362 == 8'h3c ? _GEN_482 : phv_data_241; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_487 = _GEN_4362 == 8'h3c ? _GEN_483 : phv_data_240; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_488 = mask_0[0] ? byte_ : phv_data_247; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_489 = mask_0[1] ? byte_1 : phv_data_246; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_490 = mask_0[2] ? byte_2 : phv_data_245; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_491 = mask_0[3] ? byte_3 : phv_data_244; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_492 = _GEN_4362 == 8'h3d ? _GEN_488 : phv_data_247; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_493 = _GEN_4362 == 8'h3d ? _GEN_489 : phv_data_246; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_494 = _GEN_4362 == 8'h3d ? _GEN_490 : phv_data_245; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_495 = _GEN_4362 == 8'h3d ? _GEN_491 : phv_data_244; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_496 = mask_0[0] ? byte_ : phv_data_251; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_497 = mask_0[1] ? byte_1 : phv_data_250; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_498 = mask_0[2] ? byte_2 : phv_data_249; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_499 = mask_0[3] ? byte_3 : phv_data_248; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_500 = _GEN_4362 == 8'h3e ? _GEN_496 : phv_data_251; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_501 = _GEN_4362 == 8'h3e ? _GEN_497 : phv_data_250; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_502 = _GEN_4362 == 8'h3e ? _GEN_498 : phv_data_249; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_503 = _GEN_4362 == 8'h3e ? _GEN_499 : phv_data_248; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_504 = mask_0[0] ? byte_ : phv_data_255; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_505 = mask_0[1] ? byte_1 : phv_data_254; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_506 = mask_0[2] ? byte_2 : phv_data_253; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_507 = mask_0[3] ? byte_3 : phv_data_252; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_508 = _GEN_4362 == 8'h3f ? _GEN_504 : phv_data_255; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_509 = _GEN_4362 == 8'h3f ? _GEN_505 : phv_data_254; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_510 = _GEN_4362 == 8'h3f ? _GEN_506 : phv_data_253; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_511 = _GEN_4362 == 8'h3f ? _GEN_507 : phv_data_252; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_512 = opcode != 4'h0 ? _GEN_4 : phv_data_3; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_513 = opcode != 4'h0 ? _GEN_5 : phv_data_2; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_514 = opcode != 4'h0 ? _GEN_6 : phv_data_1; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_515 = opcode != 4'h0 ? _GEN_7 : phv_data_0; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_516 = opcode != 4'h0 ? _GEN_12 : phv_data_7; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_517 = opcode != 4'h0 ? _GEN_13 : phv_data_6; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_518 = opcode != 4'h0 ? _GEN_14 : phv_data_5; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_519 = opcode != 4'h0 ? _GEN_15 : phv_data_4; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_520 = opcode != 4'h0 ? _GEN_20 : phv_data_11; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_521 = opcode != 4'h0 ? _GEN_21 : phv_data_10; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_522 = opcode != 4'h0 ? _GEN_22 : phv_data_9; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_523 = opcode != 4'h0 ? _GEN_23 : phv_data_8; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_524 = opcode != 4'h0 ? _GEN_28 : phv_data_15; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_525 = opcode != 4'h0 ? _GEN_29 : phv_data_14; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_526 = opcode != 4'h0 ? _GEN_30 : phv_data_13; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_527 = opcode != 4'h0 ? _GEN_31 : phv_data_12; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_528 = opcode != 4'h0 ? _GEN_36 : phv_data_19; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_529 = opcode != 4'h0 ? _GEN_37 : phv_data_18; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_530 = opcode != 4'h0 ? _GEN_38 : phv_data_17; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_531 = opcode != 4'h0 ? _GEN_39 : phv_data_16; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_532 = opcode != 4'h0 ? _GEN_44 : phv_data_23; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_533 = opcode != 4'h0 ? _GEN_45 : phv_data_22; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_534 = opcode != 4'h0 ? _GEN_46 : phv_data_21; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_535 = opcode != 4'h0 ? _GEN_47 : phv_data_20; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_536 = opcode != 4'h0 ? _GEN_52 : phv_data_27; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_537 = opcode != 4'h0 ? _GEN_53 : phv_data_26; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_538 = opcode != 4'h0 ? _GEN_54 : phv_data_25; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_539 = opcode != 4'h0 ? _GEN_55 : phv_data_24; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_540 = opcode != 4'h0 ? _GEN_60 : phv_data_31; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_541 = opcode != 4'h0 ? _GEN_61 : phv_data_30; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_542 = opcode != 4'h0 ? _GEN_62 : phv_data_29; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_543 = opcode != 4'h0 ? _GEN_63 : phv_data_28; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_544 = opcode != 4'h0 ? _GEN_68 : phv_data_35; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_545 = opcode != 4'h0 ? _GEN_69 : phv_data_34; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_546 = opcode != 4'h0 ? _GEN_70 : phv_data_33; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_547 = opcode != 4'h0 ? _GEN_71 : phv_data_32; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_548 = opcode != 4'h0 ? _GEN_76 : phv_data_39; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_549 = opcode != 4'h0 ? _GEN_77 : phv_data_38; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_550 = opcode != 4'h0 ? _GEN_78 : phv_data_37; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_551 = opcode != 4'h0 ? _GEN_79 : phv_data_36; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_552 = opcode != 4'h0 ? _GEN_84 : phv_data_43; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_553 = opcode != 4'h0 ? _GEN_85 : phv_data_42; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_554 = opcode != 4'h0 ? _GEN_86 : phv_data_41; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_555 = opcode != 4'h0 ? _GEN_87 : phv_data_40; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_556 = opcode != 4'h0 ? _GEN_92 : phv_data_47; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_557 = opcode != 4'h0 ? _GEN_93 : phv_data_46; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_558 = opcode != 4'h0 ? _GEN_94 : phv_data_45; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_559 = opcode != 4'h0 ? _GEN_95 : phv_data_44; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_560 = opcode != 4'h0 ? _GEN_100 : phv_data_51; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_561 = opcode != 4'h0 ? _GEN_101 : phv_data_50; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_562 = opcode != 4'h0 ? _GEN_102 : phv_data_49; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_563 = opcode != 4'h0 ? _GEN_103 : phv_data_48; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_564 = opcode != 4'h0 ? _GEN_108 : phv_data_55; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_565 = opcode != 4'h0 ? _GEN_109 : phv_data_54; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_566 = opcode != 4'h0 ? _GEN_110 : phv_data_53; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_567 = opcode != 4'h0 ? _GEN_111 : phv_data_52; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_568 = opcode != 4'h0 ? _GEN_116 : phv_data_59; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_569 = opcode != 4'h0 ? _GEN_117 : phv_data_58; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_570 = opcode != 4'h0 ? _GEN_118 : phv_data_57; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_571 = opcode != 4'h0 ? _GEN_119 : phv_data_56; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_572 = opcode != 4'h0 ? _GEN_124 : phv_data_63; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_573 = opcode != 4'h0 ? _GEN_125 : phv_data_62; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_574 = opcode != 4'h0 ? _GEN_126 : phv_data_61; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_575 = opcode != 4'h0 ? _GEN_127 : phv_data_60; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_576 = opcode != 4'h0 ? _GEN_132 : phv_data_67; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_577 = opcode != 4'h0 ? _GEN_133 : phv_data_66; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_578 = opcode != 4'h0 ? _GEN_134 : phv_data_65; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_579 = opcode != 4'h0 ? _GEN_135 : phv_data_64; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_580 = opcode != 4'h0 ? _GEN_140 : phv_data_71; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_581 = opcode != 4'h0 ? _GEN_141 : phv_data_70; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_582 = opcode != 4'h0 ? _GEN_142 : phv_data_69; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_583 = opcode != 4'h0 ? _GEN_143 : phv_data_68; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_584 = opcode != 4'h0 ? _GEN_148 : phv_data_75; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_585 = opcode != 4'h0 ? _GEN_149 : phv_data_74; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_586 = opcode != 4'h0 ? _GEN_150 : phv_data_73; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_587 = opcode != 4'h0 ? _GEN_151 : phv_data_72; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_588 = opcode != 4'h0 ? _GEN_156 : phv_data_79; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_589 = opcode != 4'h0 ? _GEN_157 : phv_data_78; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_590 = opcode != 4'h0 ? _GEN_158 : phv_data_77; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_591 = opcode != 4'h0 ? _GEN_159 : phv_data_76; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_592 = opcode != 4'h0 ? _GEN_164 : phv_data_83; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_593 = opcode != 4'h0 ? _GEN_165 : phv_data_82; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_594 = opcode != 4'h0 ? _GEN_166 : phv_data_81; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_595 = opcode != 4'h0 ? _GEN_167 : phv_data_80; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_596 = opcode != 4'h0 ? _GEN_172 : phv_data_87; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_597 = opcode != 4'h0 ? _GEN_173 : phv_data_86; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_598 = opcode != 4'h0 ? _GEN_174 : phv_data_85; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_599 = opcode != 4'h0 ? _GEN_175 : phv_data_84; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_600 = opcode != 4'h0 ? _GEN_180 : phv_data_91; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_601 = opcode != 4'h0 ? _GEN_181 : phv_data_90; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_602 = opcode != 4'h0 ? _GEN_182 : phv_data_89; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_603 = opcode != 4'h0 ? _GEN_183 : phv_data_88; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_604 = opcode != 4'h0 ? _GEN_188 : phv_data_95; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_605 = opcode != 4'h0 ? _GEN_189 : phv_data_94; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_606 = opcode != 4'h0 ? _GEN_190 : phv_data_93; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_607 = opcode != 4'h0 ? _GEN_191 : phv_data_92; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_608 = opcode != 4'h0 ? _GEN_196 : phv_data_99; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_609 = opcode != 4'h0 ? _GEN_197 : phv_data_98; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_610 = opcode != 4'h0 ? _GEN_198 : phv_data_97; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_611 = opcode != 4'h0 ? _GEN_199 : phv_data_96; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_612 = opcode != 4'h0 ? _GEN_204 : phv_data_103; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_613 = opcode != 4'h0 ? _GEN_205 : phv_data_102; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_614 = opcode != 4'h0 ? _GEN_206 : phv_data_101; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_615 = opcode != 4'h0 ? _GEN_207 : phv_data_100; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_616 = opcode != 4'h0 ? _GEN_212 : phv_data_107; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_617 = opcode != 4'h0 ? _GEN_213 : phv_data_106; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_618 = opcode != 4'h0 ? _GEN_214 : phv_data_105; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_619 = opcode != 4'h0 ? _GEN_215 : phv_data_104; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_620 = opcode != 4'h0 ? _GEN_220 : phv_data_111; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_621 = opcode != 4'h0 ? _GEN_221 : phv_data_110; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_622 = opcode != 4'h0 ? _GEN_222 : phv_data_109; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_623 = opcode != 4'h0 ? _GEN_223 : phv_data_108; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_624 = opcode != 4'h0 ? _GEN_228 : phv_data_115; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_625 = opcode != 4'h0 ? _GEN_229 : phv_data_114; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_626 = opcode != 4'h0 ? _GEN_230 : phv_data_113; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_627 = opcode != 4'h0 ? _GEN_231 : phv_data_112; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_628 = opcode != 4'h0 ? _GEN_236 : phv_data_119; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_629 = opcode != 4'h0 ? _GEN_237 : phv_data_118; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_630 = opcode != 4'h0 ? _GEN_238 : phv_data_117; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_631 = opcode != 4'h0 ? _GEN_239 : phv_data_116; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_632 = opcode != 4'h0 ? _GEN_244 : phv_data_123; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_633 = opcode != 4'h0 ? _GEN_245 : phv_data_122; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_634 = opcode != 4'h0 ? _GEN_246 : phv_data_121; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_635 = opcode != 4'h0 ? _GEN_247 : phv_data_120; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_636 = opcode != 4'h0 ? _GEN_252 : phv_data_127; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_637 = opcode != 4'h0 ? _GEN_253 : phv_data_126; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_638 = opcode != 4'h0 ? _GEN_254 : phv_data_125; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_639 = opcode != 4'h0 ? _GEN_255 : phv_data_124; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_640 = opcode != 4'h0 ? _GEN_260 : phv_data_131; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_641 = opcode != 4'h0 ? _GEN_261 : phv_data_130; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_642 = opcode != 4'h0 ? _GEN_262 : phv_data_129; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_643 = opcode != 4'h0 ? _GEN_263 : phv_data_128; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_644 = opcode != 4'h0 ? _GEN_268 : phv_data_135; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_645 = opcode != 4'h0 ? _GEN_269 : phv_data_134; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_646 = opcode != 4'h0 ? _GEN_270 : phv_data_133; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_647 = opcode != 4'h0 ? _GEN_271 : phv_data_132; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_648 = opcode != 4'h0 ? _GEN_276 : phv_data_139; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_649 = opcode != 4'h0 ? _GEN_277 : phv_data_138; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_650 = opcode != 4'h0 ? _GEN_278 : phv_data_137; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_651 = opcode != 4'h0 ? _GEN_279 : phv_data_136; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_652 = opcode != 4'h0 ? _GEN_284 : phv_data_143; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_653 = opcode != 4'h0 ? _GEN_285 : phv_data_142; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_654 = opcode != 4'h0 ? _GEN_286 : phv_data_141; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_655 = opcode != 4'h0 ? _GEN_287 : phv_data_140; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_656 = opcode != 4'h0 ? _GEN_292 : phv_data_147; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_657 = opcode != 4'h0 ? _GEN_293 : phv_data_146; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_658 = opcode != 4'h0 ? _GEN_294 : phv_data_145; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_659 = opcode != 4'h0 ? _GEN_295 : phv_data_144; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_660 = opcode != 4'h0 ? _GEN_300 : phv_data_151; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_661 = opcode != 4'h0 ? _GEN_301 : phv_data_150; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_662 = opcode != 4'h0 ? _GEN_302 : phv_data_149; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_663 = opcode != 4'h0 ? _GEN_303 : phv_data_148; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_664 = opcode != 4'h0 ? _GEN_308 : phv_data_155; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_665 = opcode != 4'h0 ? _GEN_309 : phv_data_154; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_666 = opcode != 4'h0 ? _GEN_310 : phv_data_153; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_667 = opcode != 4'h0 ? _GEN_311 : phv_data_152; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_668 = opcode != 4'h0 ? _GEN_316 : phv_data_159; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_669 = opcode != 4'h0 ? _GEN_317 : phv_data_158; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_670 = opcode != 4'h0 ? _GEN_318 : phv_data_157; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_671 = opcode != 4'h0 ? _GEN_319 : phv_data_156; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_672 = opcode != 4'h0 ? _GEN_324 : phv_data_163; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_673 = opcode != 4'h0 ? _GEN_325 : phv_data_162; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_674 = opcode != 4'h0 ? _GEN_326 : phv_data_161; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_675 = opcode != 4'h0 ? _GEN_327 : phv_data_160; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_676 = opcode != 4'h0 ? _GEN_332 : phv_data_167; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_677 = opcode != 4'h0 ? _GEN_333 : phv_data_166; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_678 = opcode != 4'h0 ? _GEN_334 : phv_data_165; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_679 = opcode != 4'h0 ? _GEN_335 : phv_data_164; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_680 = opcode != 4'h0 ? _GEN_340 : phv_data_171; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_681 = opcode != 4'h0 ? _GEN_341 : phv_data_170; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_682 = opcode != 4'h0 ? _GEN_342 : phv_data_169; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_683 = opcode != 4'h0 ? _GEN_343 : phv_data_168; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_684 = opcode != 4'h0 ? _GEN_348 : phv_data_175; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_685 = opcode != 4'h0 ? _GEN_349 : phv_data_174; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_686 = opcode != 4'h0 ? _GEN_350 : phv_data_173; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_687 = opcode != 4'h0 ? _GEN_351 : phv_data_172; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_688 = opcode != 4'h0 ? _GEN_356 : phv_data_179; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_689 = opcode != 4'h0 ? _GEN_357 : phv_data_178; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_690 = opcode != 4'h0 ? _GEN_358 : phv_data_177; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_691 = opcode != 4'h0 ? _GEN_359 : phv_data_176; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_692 = opcode != 4'h0 ? _GEN_364 : phv_data_183; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_693 = opcode != 4'h0 ? _GEN_365 : phv_data_182; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_694 = opcode != 4'h0 ? _GEN_366 : phv_data_181; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_695 = opcode != 4'h0 ? _GEN_367 : phv_data_180; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_696 = opcode != 4'h0 ? _GEN_372 : phv_data_187; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_697 = opcode != 4'h0 ? _GEN_373 : phv_data_186; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_698 = opcode != 4'h0 ? _GEN_374 : phv_data_185; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_699 = opcode != 4'h0 ? _GEN_375 : phv_data_184; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_700 = opcode != 4'h0 ? _GEN_380 : phv_data_191; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_701 = opcode != 4'h0 ? _GEN_381 : phv_data_190; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_702 = opcode != 4'h0 ? _GEN_382 : phv_data_189; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_703 = opcode != 4'h0 ? _GEN_383 : phv_data_188; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_704 = opcode != 4'h0 ? _GEN_388 : phv_data_195; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_705 = opcode != 4'h0 ? _GEN_389 : phv_data_194; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_706 = opcode != 4'h0 ? _GEN_390 : phv_data_193; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_707 = opcode != 4'h0 ? _GEN_391 : phv_data_192; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_708 = opcode != 4'h0 ? _GEN_396 : phv_data_199; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_709 = opcode != 4'h0 ? _GEN_397 : phv_data_198; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_710 = opcode != 4'h0 ? _GEN_398 : phv_data_197; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_711 = opcode != 4'h0 ? _GEN_399 : phv_data_196; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_712 = opcode != 4'h0 ? _GEN_404 : phv_data_203; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_713 = opcode != 4'h0 ? _GEN_405 : phv_data_202; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_714 = opcode != 4'h0 ? _GEN_406 : phv_data_201; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_715 = opcode != 4'h0 ? _GEN_407 : phv_data_200; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_716 = opcode != 4'h0 ? _GEN_412 : phv_data_207; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_717 = opcode != 4'h0 ? _GEN_413 : phv_data_206; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_718 = opcode != 4'h0 ? _GEN_414 : phv_data_205; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_719 = opcode != 4'h0 ? _GEN_415 : phv_data_204; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_720 = opcode != 4'h0 ? _GEN_420 : phv_data_211; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_721 = opcode != 4'h0 ? _GEN_421 : phv_data_210; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_722 = opcode != 4'h0 ? _GEN_422 : phv_data_209; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_723 = opcode != 4'h0 ? _GEN_423 : phv_data_208; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_724 = opcode != 4'h0 ? _GEN_428 : phv_data_215; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_725 = opcode != 4'h0 ? _GEN_429 : phv_data_214; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_726 = opcode != 4'h0 ? _GEN_430 : phv_data_213; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_727 = opcode != 4'h0 ? _GEN_431 : phv_data_212; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_728 = opcode != 4'h0 ? _GEN_436 : phv_data_219; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_729 = opcode != 4'h0 ? _GEN_437 : phv_data_218; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_730 = opcode != 4'h0 ? _GEN_438 : phv_data_217; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_731 = opcode != 4'h0 ? _GEN_439 : phv_data_216; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_732 = opcode != 4'h0 ? _GEN_444 : phv_data_223; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_733 = opcode != 4'h0 ? _GEN_445 : phv_data_222; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_734 = opcode != 4'h0 ? _GEN_446 : phv_data_221; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_735 = opcode != 4'h0 ? _GEN_447 : phv_data_220; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_736 = opcode != 4'h0 ? _GEN_452 : phv_data_227; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_737 = opcode != 4'h0 ? _GEN_453 : phv_data_226; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_738 = opcode != 4'h0 ? _GEN_454 : phv_data_225; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_739 = opcode != 4'h0 ? _GEN_455 : phv_data_224; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_740 = opcode != 4'h0 ? _GEN_460 : phv_data_231; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_741 = opcode != 4'h0 ? _GEN_461 : phv_data_230; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_742 = opcode != 4'h0 ? _GEN_462 : phv_data_229; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_743 = opcode != 4'h0 ? _GEN_463 : phv_data_228; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_744 = opcode != 4'h0 ? _GEN_468 : phv_data_235; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_745 = opcode != 4'h0 ? _GEN_469 : phv_data_234; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_746 = opcode != 4'h0 ? _GEN_470 : phv_data_233; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_747 = opcode != 4'h0 ? _GEN_471 : phv_data_232; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_748 = opcode != 4'h0 ? _GEN_476 : phv_data_239; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_749 = opcode != 4'h0 ? _GEN_477 : phv_data_238; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_750 = opcode != 4'h0 ? _GEN_478 : phv_data_237; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_751 = opcode != 4'h0 ? _GEN_479 : phv_data_236; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_752 = opcode != 4'h0 ? _GEN_484 : phv_data_243; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_753 = opcode != 4'h0 ? _GEN_485 : phv_data_242; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_754 = opcode != 4'h0 ? _GEN_486 : phv_data_241; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_755 = opcode != 4'h0 ? _GEN_487 : phv_data_240; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_756 = opcode != 4'h0 ? _GEN_492 : phv_data_247; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_757 = opcode != 4'h0 ? _GEN_493 : phv_data_246; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_758 = opcode != 4'h0 ? _GEN_494 : phv_data_245; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_759 = opcode != 4'h0 ? _GEN_495 : phv_data_244; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_760 = opcode != 4'h0 ? _GEN_500 : phv_data_251; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_761 = opcode != 4'h0 ? _GEN_501 : phv_data_250; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_762 = opcode != 4'h0 ? _GEN_502 : phv_data_249; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_763 = opcode != 4'h0 ? _GEN_503 : phv_data_248; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_764 = opcode != 4'h0 ? _GEN_508 : phv_data_255; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_765 = opcode != 4'h0 ? _GEN_509 : phv_data_254; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_766 = opcode != 4'h0 ? _GEN_510 : phv_data_253; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_767 = opcode != 4'h0 ? _GEN_511 : phv_data_252; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_770 = opcode == 4'hf ? phv_data_3 : _GEN_512; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_771 = opcode == 4'hf ? phv_data_2 : _GEN_513; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_772 = opcode == 4'hf ? phv_data_1 : _GEN_514; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_773 = opcode == 4'hf ? phv_data_0 : _GEN_515; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_774 = opcode == 4'hf ? phv_data_7 : _GEN_516; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_775 = opcode == 4'hf ? phv_data_6 : _GEN_517; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_776 = opcode == 4'hf ? phv_data_5 : _GEN_518; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_777 = opcode == 4'hf ? phv_data_4 : _GEN_519; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_778 = opcode == 4'hf ? phv_data_11 : _GEN_520; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_779 = opcode == 4'hf ? phv_data_10 : _GEN_521; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_780 = opcode == 4'hf ? phv_data_9 : _GEN_522; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_781 = opcode == 4'hf ? phv_data_8 : _GEN_523; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_782 = opcode == 4'hf ? phv_data_15 : _GEN_524; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_783 = opcode == 4'hf ? phv_data_14 : _GEN_525; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_784 = opcode == 4'hf ? phv_data_13 : _GEN_526; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_785 = opcode == 4'hf ? phv_data_12 : _GEN_527; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_786 = opcode == 4'hf ? phv_data_19 : _GEN_528; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_787 = opcode == 4'hf ? phv_data_18 : _GEN_529; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_788 = opcode == 4'hf ? phv_data_17 : _GEN_530; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_789 = opcode == 4'hf ? phv_data_16 : _GEN_531; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_790 = opcode == 4'hf ? phv_data_23 : _GEN_532; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_791 = opcode == 4'hf ? phv_data_22 : _GEN_533; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_792 = opcode == 4'hf ? phv_data_21 : _GEN_534; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_793 = opcode == 4'hf ? phv_data_20 : _GEN_535; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_794 = opcode == 4'hf ? phv_data_27 : _GEN_536; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_795 = opcode == 4'hf ? phv_data_26 : _GEN_537; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_796 = opcode == 4'hf ? phv_data_25 : _GEN_538; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_797 = opcode == 4'hf ? phv_data_24 : _GEN_539; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_798 = opcode == 4'hf ? phv_data_31 : _GEN_540; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_799 = opcode == 4'hf ? phv_data_30 : _GEN_541; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_800 = opcode == 4'hf ? phv_data_29 : _GEN_542; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_801 = opcode == 4'hf ? phv_data_28 : _GEN_543; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_802 = opcode == 4'hf ? phv_data_35 : _GEN_544; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_803 = opcode == 4'hf ? phv_data_34 : _GEN_545; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_804 = opcode == 4'hf ? phv_data_33 : _GEN_546; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_805 = opcode == 4'hf ? phv_data_32 : _GEN_547; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_806 = opcode == 4'hf ? phv_data_39 : _GEN_548; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_807 = opcode == 4'hf ? phv_data_38 : _GEN_549; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_808 = opcode == 4'hf ? phv_data_37 : _GEN_550; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_809 = opcode == 4'hf ? phv_data_36 : _GEN_551; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_810 = opcode == 4'hf ? phv_data_43 : _GEN_552; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_811 = opcode == 4'hf ? phv_data_42 : _GEN_553; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_812 = opcode == 4'hf ? phv_data_41 : _GEN_554; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_813 = opcode == 4'hf ? phv_data_40 : _GEN_555; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_814 = opcode == 4'hf ? phv_data_47 : _GEN_556; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_815 = opcode == 4'hf ? phv_data_46 : _GEN_557; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_816 = opcode == 4'hf ? phv_data_45 : _GEN_558; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_817 = opcode == 4'hf ? phv_data_44 : _GEN_559; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_818 = opcode == 4'hf ? phv_data_51 : _GEN_560; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_819 = opcode == 4'hf ? phv_data_50 : _GEN_561; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_820 = opcode == 4'hf ? phv_data_49 : _GEN_562; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_821 = opcode == 4'hf ? phv_data_48 : _GEN_563; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_822 = opcode == 4'hf ? phv_data_55 : _GEN_564; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_823 = opcode == 4'hf ? phv_data_54 : _GEN_565; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_824 = opcode == 4'hf ? phv_data_53 : _GEN_566; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_825 = opcode == 4'hf ? phv_data_52 : _GEN_567; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_826 = opcode == 4'hf ? phv_data_59 : _GEN_568; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_827 = opcode == 4'hf ? phv_data_58 : _GEN_569; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_828 = opcode == 4'hf ? phv_data_57 : _GEN_570; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_829 = opcode == 4'hf ? phv_data_56 : _GEN_571; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_830 = opcode == 4'hf ? phv_data_63 : _GEN_572; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_831 = opcode == 4'hf ? phv_data_62 : _GEN_573; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_832 = opcode == 4'hf ? phv_data_61 : _GEN_574; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_833 = opcode == 4'hf ? phv_data_60 : _GEN_575; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_834 = opcode == 4'hf ? phv_data_67 : _GEN_576; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_835 = opcode == 4'hf ? phv_data_66 : _GEN_577; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_836 = opcode == 4'hf ? phv_data_65 : _GEN_578; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_837 = opcode == 4'hf ? phv_data_64 : _GEN_579; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_838 = opcode == 4'hf ? phv_data_71 : _GEN_580; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_839 = opcode == 4'hf ? phv_data_70 : _GEN_581; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_840 = opcode == 4'hf ? phv_data_69 : _GEN_582; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_841 = opcode == 4'hf ? phv_data_68 : _GEN_583; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_842 = opcode == 4'hf ? phv_data_75 : _GEN_584; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_843 = opcode == 4'hf ? phv_data_74 : _GEN_585; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_844 = opcode == 4'hf ? phv_data_73 : _GEN_586; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_845 = opcode == 4'hf ? phv_data_72 : _GEN_587; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_846 = opcode == 4'hf ? phv_data_79 : _GEN_588; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_847 = opcode == 4'hf ? phv_data_78 : _GEN_589; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_848 = opcode == 4'hf ? phv_data_77 : _GEN_590; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_849 = opcode == 4'hf ? phv_data_76 : _GEN_591; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_850 = opcode == 4'hf ? phv_data_83 : _GEN_592; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_851 = opcode == 4'hf ? phv_data_82 : _GEN_593; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_852 = opcode == 4'hf ? phv_data_81 : _GEN_594; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_853 = opcode == 4'hf ? phv_data_80 : _GEN_595; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_854 = opcode == 4'hf ? phv_data_87 : _GEN_596; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_855 = opcode == 4'hf ? phv_data_86 : _GEN_597; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_856 = opcode == 4'hf ? phv_data_85 : _GEN_598; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_857 = opcode == 4'hf ? phv_data_84 : _GEN_599; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_858 = opcode == 4'hf ? phv_data_91 : _GEN_600; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_859 = opcode == 4'hf ? phv_data_90 : _GEN_601; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_860 = opcode == 4'hf ? phv_data_89 : _GEN_602; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_861 = opcode == 4'hf ? phv_data_88 : _GEN_603; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_862 = opcode == 4'hf ? phv_data_95 : _GEN_604; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_863 = opcode == 4'hf ? phv_data_94 : _GEN_605; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_864 = opcode == 4'hf ? phv_data_93 : _GEN_606; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_865 = opcode == 4'hf ? phv_data_92 : _GEN_607; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_866 = opcode == 4'hf ? phv_data_99 : _GEN_608; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_867 = opcode == 4'hf ? phv_data_98 : _GEN_609; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_868 = opcode == 4'hf ? phv_data_97 : _GEN_610; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_869 = opcode == 4'hf ? phv_data_96 : _GEN_611; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_870 = opcode == 4'hf ? phv_data_103 : _GEN_612; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_871 = opcode == 4'hf ? phv_data_102 : _GEN_613; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_872 = opcode == 4'hf ? phv_data_101 : _GEN_614; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_873 = opcode == 4'hf ? phv_data_100 : _GEN_615; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_874 = opcode == 4'hf ? phv_data_107 : _GEN_616; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_875 = opcode == 4'hf ? phv_data_106 : _GEN_617; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_876 = opcode == 4'hf ? phv_data_105 : _GEN_618; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_877 = opcode == 4'hf ? phv_data_104 : _GEN_619; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_878 = opcode == 4'hf ? phv_data_111 : _GEN_620; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_879 = opcode == 4'hf ? phv_data_110 : _GEN_621; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_880 = opcode == 4'hf ? phv_data_109 : _GEN_622; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_881 = opcode == 4'hf ? phv_data_108 : _GEN_623; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_882 = opcode == 4'hf ? phv_data_115 : _GEN_624; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_883 = opcode == 4'hf ? phv_data_114 : _GEN_625; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_884 = opcode == 4'hf ? phv_data_113 : _GEN_626; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_885 = opcode == 4'hf ? phv_data_112 : _GEN_627; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_886 = opcode == 4'hf ? phv_data_119 : _GEN_628; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_887 = opcode == 4'hf ? phv_data_118 : _GEN_629; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_888 = opcode == 4'hf ? phv_data_117 : _GEN_630; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_889 = opcode == 4'hf ? phv_data_116 : _GEN_631; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_890 = opcode == 4'hf ? phv_data_123 : _GEN_632; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_891 = opcode == 4'hf ? phv_data_122 : _GEN_633; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_892 = opcode == 4'hf ? phv_data_121 : _GEN_634; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_893 = opcode == 4'hf ? phv_data_120 : _GEN_635; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_894 = opcode == 4'hf ? phv_data_127 : _GEN_636; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_895 = opcode == 4'hf ? phv_data_126 : _GEN_637; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_896 = opcode == 4'hf ? phv_data_125 : _GEN_638; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_897 = opcode == 4'hf ? phv_data_124 : _GEN_639; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_898 = opcode == 4'hf ? phv_data_131 : _GEN_640; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_899 = opcode == 4'hf ? phv_data_130 : _GEN_641; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_900 = opcode == 4'hf ? phv_data_129 : _GEN_642; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_901 = opcode == 4'hf ? phv_data_128 : _GEN_643; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_902 = opcode == 4'hf ? phv_data_135 : _GEN_644; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_903 = opcode == 4'hf ? phv_data_134 : _GEN_645; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_904 = opcode == 4'hf ? phv_data_133 : _GEN_646; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_905 = opcode == 4'hf ? phv_data_132 : _GEN_647; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_906 = opcode == 4'hf ? phv_data_139 : _GEN_648; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_907 = opcode == 4'hf ? phv_data_138 : _GEN_649; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_908 = opcode == 4'hf ? phv_data_137 : _GEN_650; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_909 = opcode == 4'hf ? phv_data_136 : _GEN_651; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_910 = opcode == 4'hf ? phv_data_143 : _GEN_652; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_911 = opcode == 4'hf ? phv_data_142 : _GEN_653; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_912 = opcode == 4'hf ? phv_data_141 : _GEN_654; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_913 = opcode == 4'hf ? phv_data_140 : _GEN_655; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_914 = opcode == 4'hf ? phv_data_147 : _GEN_656; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_915 = opcode == 4'hf ? phv_data_146 : _GEN_657; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_916 = opcode == 4'hf ? phv_data_145 : _GEN_658; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_917 = opcode == 4'hf ? phv_data_144 : _GEN_659; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_918 = opcode == 4'hf ? phv_data_151 : _GEN_660; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_919 = opcode == 4'hf ? phv_data_150 : _GEN_661; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_920 = opcode == 4'hf ? phv_data_149 : _GEN_662; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_921 = opcode == 4'hf ? phv_data_148 : _GEN_663; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_922 = opcode == 4'hf ? phv_data_155 : _GEN_664; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_923 = opcode == 4'hf ? phv_data_154 : _GEN_665; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_924 = opcode == 4'hf ? phv_data_153 : _GEN_666; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_925 = opcode == 4'hf ? phv_data_152 : _GEN_667; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_926 = opcode == 4'hf ? phv_data_159 : _GEN_668; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_927 = opcode == 4'hf ? phv_data_158 : _GEN_669; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_928 = opcode == 4'hf ? phv_data_157 : _GEN_670; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_929 = opcode == 4'hf ? phv_data_156 : _GEN_671; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_930 = opcode == 4'hf ? phv_data_163 : _GEN_672; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_931 = opcode == 4'hf ? phv_data_162 : _GEN_673; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_932 = opcode == 4'hf ? phv_data_161 : _GEN_674; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_933 = opcode == 4'hf ? phv_data_160 : _GEN_675; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_934 = opcode == 4'hf ? phv_data_167 : _GEN_676; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_935 = opcode == 4'hf ? phv_data_166 : _GEN_677; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_936 = opcode == 4'hf ? phv_data_165 : _GEN_678; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_937 = opcode == 4'hf ? phv_data_164 : _GEN_679; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_938 = opcode == 4'hf ? phv_data_171 : _GEN_680; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_939 = opcode == 4'hf ? phv_data_170 : _GEN_681; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_940 = opcode == 4'hf ? phv_data_169 : _GEN_682; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_941 = opcode == 4'hf ? phv_data_168 : _GEN_683; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_942 = opcode == 4'hf ? phv_data_175 : _GEN_684; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_943 = opcode == 4'hf ? phv_data_174 : _GEN_685; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_944 = opcode == 4'hf ? phv_data_173 : _GEN_686; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_945 = opcode == 4'hf ? phv_data_172 : _GEN_687; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_946 = opcode == 4'hf ? phv_data_179 : _GEN_688; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_947 = opcode == 4'hf ? phv_data_178 : _GEN_689; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_948 = opcode == 4'hf ? phv_data_177 : _GEN_690; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_949 = opcode == 4'hf ? phv_data_176 : _GEN_691; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_950 = opcode == 4'hf ? phv_data_183 : _GEN_692; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_951 = opcode == 4'hf ? phv_data_182 : _GEN_693; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_952 = opcode == 4'hf ? phv_data_181 : _GEN_694; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_953 = opcode == 4'hf ? phv_data_180 : _GEN_695; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_954 = opcode == 4'hf ? phv_data_187 : _GEN_696; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_955 = opcode == 4'hf ? phv_data_186 : _GEN_697; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_956 = opcode == 4'hf ? phv_data_185 : _GEN_698; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_957 = opcode == 4'hf ? phv_data_184 : _GEN_699; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_958 = opcode == 4'hf ? phv_data_191 : _GEN_700; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_959 = opcode == 4'hf ? phv_data_190 : _GEN_701; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_960 = opcode == 4'hf ? phv_data_189 : _GEN_702; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_961 = opcode == 4'hf ? phv_data_188 : _GEN_703; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_962 = opcode == 4'hf ? phv_data_195 : _GEN_704; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_963 = opcode == 4'hf ? phv_data_194 : _GEN_705; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_964 = opcode == 4'hf ? phv_data_193 : _GEN_706; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_965 = opcode == 4'hf ? phv_data_192 : _GEN_707; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_966 = opcode == 4'hf ? phv_data_199 : _GEN_708; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_967 = opcode == 4'hf ? phv_data_198 : _GEN_709; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_968 = opcode == 4'hf ? phv_data_197 : _GEN_710; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_969 = opcode == 4'hf ? phv_data_196 : _GEN_711; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_970 = opcode == 4'hf ? phv_data_203 : _GEN_712; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_971 = opcode == 4'hf ? phv_data_202 : _GEN_713; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_972 = opcode == 4'hf ? phv_data_201 : _GEN_714; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_973 = opcode == 4'hf ? phv_data_200 : _GEN_715; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_974 = opcode == 4'hf ? phv_data_207 : _GEN_716; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_975 = opcode == 4'hf ? phv_data_206 : _GEN_717; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_976 = opcode == 4'hf ? phv_data_205 : _GEN_718; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_977 = opcode == 4'hf ? phv_data_204 : _GEN_719; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_978 = opcode == 4'hf ? phv_data_211 : _GEN_720; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_979 = opcode == 4'hf ? phv_data_210 : _GEN_721; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_980 = opcode == 4'hf ? phv_data_209 : _GEN_722; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_981 = opcode == 4'hf ? phv_data_208 : _GEN_723; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_982 = opcode == 4'hf ? phv_data_215 : _GEN_724; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_983 = opcode == 4'hf ? phv_data_214 : _GEN_725; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_984 = opcode == 4'hf ? phv_data_213 : _GEN_726; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_985 = opcode == 4'hf ? phv_data_212 : _GEN_727; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_986 = opcode == 4'hf ? phv_data_219 : _GEN_728; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_987 = opcode == 4'hf ? phv_data_218 : _GEN_729; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_988 = opcode == 4'hf ? phv_data_217 : _GEN_730; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_989 = opcode == 4'hf ? phv_data_216 : _GEN_731; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_990 = opcode == 4'hf ? phv_data_223 : _GEN_732; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_991 = opcode == 4'hf ? phv_data_222 : _GEN_733; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_992 = opcode == 4'hf ? phv_data_221 : _GEN_734; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_993 = opcode == 4'hf ? phv_data_220 : _GEN_735; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_994 = opcode == 4'hf ? phv_data_227 : _GEN_736; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_995 = opcode == 4'hf ? phv_data_226 : _GEN_737; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_996 = opcode == 4'hf ? phv_data_225 : _GEN_738; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_997 = opcode == 4'hf ? phv_data_224 : _GEN_739; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_998 = opcode == 4'hf ? phv_data_231 : _GEN_740; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_999 = opcode == 4'hf ? phv_data_230 : _GEN_741; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1000 = opcode == 4'hf ? phv_data_229 : _GEN_742; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1001 = opcode == 4'hf ? phv_data_228 : _GEN_743; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1002 = opcode == 4'hf ? phv_data_235 : _GEN_744; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1003 = opcode == 4'hf ? phv_data_234 : _GEN_745; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1004 = opcode == 4'hf ? phv_data_233 : _GEN_746; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1005 = opcode == 4'hf ? phv_data_232 : _GEN_747; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1006 = opcode == 4'hf ? phv_data_239 : _GEN_748; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1007 = opcode == 4'hf ? phv_data_238 : _GEN_749; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1008 = opcode == 4'hf ? phv_data_237 : _GEN_750; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1009 = opcode == 4'hf ? phv_data_236 : _GEN_751; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1010 = opcode == 4'hf ? phv_data_243 : _GEN_752; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1011 = opcode == 4'hf ? phv_data_242 : _GEN_753; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1012 = opcode == 4'hf ? phv_data_241 : _GEN_754; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1013 = opcode == 4'hf ? phv_data_240 : _GEN_755; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1014 = opcode == 4'hf ? phv_data_247 : _GEN_756; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1015 = opcode == 4'hf ? phv_data_246 : _GEN_757; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1016 = opcode == 4'hf ? phv_data_245 : _GEN_758; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1017 = opcode == 4'hf ? phv_data_244 : _GEN_759; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1018 = opcode == 4'hf ? phv_data_251 : _GEN_760; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1019 = opcode == 4'hf ? phv_data_250 : _GEN_761; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1020 = opcode == 4'hf ? phv_data_249 : _GEN_762; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1021 = opcode == 4'hf ? phv_data_248 : _GEN_763; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1022 = opcode == 4'hf ? phv_data_255 : _GEN_764; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1023 = opcode == 4'hf ? phv_data_254 : _GEN_765; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1024 = opcode == 4'hf ? phv_data_253 : _GEN_766; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1025 = opcode == 4'hf ? phv_data_252 : _GEN_767; // @[executor.scala 466:52 executor.scala 450:25]
  wire [3:0] opcode_1 = vliw_1[31:28]; // @[primitive.scala 9:44]
  wire [7:0] _GEN_4426 = {{2'd0}, dst_offset_1}; // @[executor.scala 473:49]
  wire [7:0] byte_256 = field_1[7:0]; // @[executor.scala 475:56]
  wire [7:0] _GEN_1026 = mask_1[0] ? byte_256 : _GEN_770; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] byte_257 = field_1[15:8]; // @[executor.scala 475:56]
  wire [7:0] _GEN_1027 = mask_1[1] ? byte_257 : _GEN_771; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] byte_258 = field_1[23:16]; // @[executor.scala 475:56]
  wire [7:0] _GEN_1028 = mask_1[2] ? byte_258 : _GEN_772; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] byte_259 = field_1[31:24]; // @[executor.scala 475:56]
  wire [7:0] _GEN_1029 = mask_1[3] ? byte_259 : _GEN_773; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1030 = _GEN_4426 == 8'h0 ? _GEN_1026 : _GEN_770; // @[executor.scala 473:84]
  wire [7:0] _GEN_1031 = _GEN_4426 == 8'h0 ? _GEN_1027 : _GEN_771; // @[executor.scala 473:84]
  wire [7:0] _GEN_1032 = _GEN_4426 == 8'h0 ? _GEN_1028 : _GEN_772; // @[executor.scala 473:84]
  wire [7:0] _GEN_1033 = _GEN_4426 == 8'h0 ? _GEN_1029 : _GEN_773; // @[executor.scala 473:84]
  wire [7:0] _GEN_1034 = mask_1[0] ? byte_256 : _GEN_774; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1035 = mask_1[1] ? byte_257 : _GEN_775; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1036 = mask_1[2] ? byte_258 : _GEN_776; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1037 = mask_1[3] ? byte_259 : _GEN_777; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1038 = _GEN_4426 == 8'h1 ? _GEN_1034 : _GEN_774; // @[executor.scala 473:84]
  wire [7:0] _GEN_1039 = _GEN_4426 == 8'h1 ? _GEN_1035 : _GEN_775; // @[executor.scala 473:84]
  wire [7:0] _GEN_1040 = _GEN_4426 == 8'h1 ? _GEN_1036 : _GEN_776; // @[executor.scala 473:84]
  wire [7:0] _GEN_1041 = _GEN_4426 == 8'h1 ? _GEN_1037 : _GEN_777; // @[executor.scala 473:84]
  wire [7:0] _GEN_1042 = mask_1[0] ? byte_256 : _GEN_778; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1043 = mask_1[1] ? byte_257 : _GEN_779; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1044 = mask_1[2] ? byte_258 : _GEN_780; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1045 = mask_1[3] ? byte_259 : _GEN_781; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1046 = _GEN_4426 == 8'h2 ? _GEN_1042 : _GEN_778; // @[executor.scala 473:84]
  wire [7:0] _GEN_1047 = _GEN_4426 == 8'h2 ? _GEN_1043 : _GEN_779; // @[executor.scala 473:84]
  wire [7:0] _GEN_1048 = _GEN_4426 == 8'h2 ? _GEN_1044 : _GEN_780; // @[executor.scala 473:84]
  wire [7:0] _GEN_1049 = _GEN_4426 == 8'h2 ? _GEN_1045 : _GEN_781; // @[executor.scala 473:84]
  wire [7:0] _GEN_1050 = mask_1[0] ? byte_256 : _GEN_782; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1051 = mask_1[1] ? byte_257 : _GEN_783; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1052 = mask_1[2] ? byte_258 : _GEN_784; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1053 = mask_1[3] ? byte_259 : _GEN_785; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1054 = _GEN_4426 == 8'h3 ? _GEN_1050 : _GEN_782; // @[executor.scala 473:84]
  wire [7:0] _GEN_1055 = _GEN_4426 == 8'h3 ? _GEN_1051 : _GEN_783; // @[executor.scala 473:84]
  wire [7:0] _GEN_1056 = _GEN_4426 == 8'h3 ? _GEN_1052 : _GEN_784; // @[executor.scala 473:84]
  wire [7:0] _GEN_1057 = _GEN_4426 == 8'h3 ? _GEN_1053 : _GEN_785; // @[executor.scala 473:84]
  wire [7:0] _GEN_1058 = mask_1[0] ? byte_256 : _GEN_786; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1059 = mask_1[1] ? byte_257 : _GEN_787; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1060 = mask_1[2] ? byte_258 : _GEN_788; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1061 = mask_1[3] ? byte_259 : _GEN_789; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1062 = _GEN_4426 == 8'h4 ? _GEN_1058 : _GEN_786; // @[executor.scala 473:84]
  wire [7:0] _GEN_1063 = _GEN_4426 == 8'h4 ? _GEN_1059 : _GEN_787; // @[executor.scala 473:84]
  wire [7:0] _GEN_1064 = _GEN_4426 == 8'h4 ? _GEN_1060 : _GEN_788; // @[executor.scala 473:84]
  wire [7:0] _GEN_1065 = _GEN_4426 == 8'h4 ? _GEN_1061 : _GEN_789; // @[executor.scala 473:84]
  wire [7:0] _GEN_1066 = mask_1[0] ? byte_256 : _GEN_790; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1067 = mask_1[1] ? byte_257 : _GEN_791; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1068 = mask_1[2] ? byte_258 : _GEN_792; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1069 = mask_1[3] ? byte_259 : _GEN_793; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1070 = _GEN_4426 == 8'h5 ? _GEN_1066 : _GEN_790; // @[executor.scala 473:84]
  wire [7:0] _GEN_1071 = _GEN_4426 == 8'h5 ? _GEN_1067 : _GEN_791; // @[executor.scala 473:84]
  wire [7:0] _GEN_1072 = _GEN_4426 == 8'h5 ? _GEN_1068 : _GEN_792; // @[executor.scala 473:84]
  wire [7:0] _GEN_1073 = _GEN_4426 == 8'h5 ? _GEN_1069 : _GEN_793; // @[executor.scala 473:84]
  wire [7:0] _GEN_1074 = mask_1[0] ? byte_256 : _GEN_794; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1075 = mask_1[1] ? byte_257 : _GEN_795; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1076 = mask_1[2] ? byte_258 : _GEN_796; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1077 = mask_1[3] ? byte_259 : _GEN_797; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1078 = _GEN_4426 == 8'h6 ? _GEN_1074 : _GEN_794; // @[executor.scala 473:84]
  wire [7:0] _GEN_1079 = _GEN_4426 == 8'h6 ? _GEN_1075 : _GEN_795; // @[executor.scala 473:84]
  wire [7:0] _GEN_1080 = _GEN_4426 == 8'h6 ? _GEN_1076 : _GEN_796; // @[executor.scala 473:84]
  wire [7:0] _GEN_1081 = _GEN_4426 == 8'h6 ? _GEN_1077 : _GEN_797; // @[executor.scala 473:84]
  wire [7:0] _GEN_1082 = mask_1[0] ? byte_256 : _GEN_798; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1083 = mask_1[1] ? byte_257 : _GEN_799; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1084 = mask_1[2] ? byte_258 : _GEN_800; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1085 = mask_1[3] ? byte_259 : _GEN_801; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1086 = _GEN_4426 == 8'h7 ? _GEN_1082 : _GEN_798; // @[executor.scala 473:84]
  wire [7:0] _GEN_1087 = _GEN_4426 == 8'h7 ? _GEN_1083 : _GEN_799; // @[executor.scala 473:84]
  wire [7:0] _GEN_1088 = _GEN_4426 == 8'h7 ? _GEN_1084 : _GEN_800; // @[executor.scala 473:84]
  wire [7:0] _GEN_1089 = _GEN_4426 == 8'h7 ? _GEN_1085 : _GEN_801; // @[executor.scala 473:84]
  wire [7:0] _GEN_1090 = mask_1[0] ? byte_256 : _GEN_802; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1091 = mask_1[1] ? byte_257 : _GEN_803; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1092 = mask_1[2] ? byte_258 : _GEN_804; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1093 = mask_1[3] ? byte_259 : _GEN_805; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1094 = _GEN_4426 == 8'h8 ? _GEN_1090 : _GEN_802; // @[executor.scala 473:84]
  wire [7:0] _GEN_1095 = _GEN_4426 == 8'h8 ? _GEN_1091 : _GEN_803; // @[executor.scala 473:84]
  wire [7:0] _GEN_1096 = _GEN_4426 == 8'h8 ? _GEN_1092 : _GEN_804; // @[executor.scala 473:84]
  wire [7:0] _GEN_1097 = _GEN_4426 == 8'h8 ? _GEN_1093 : _GEN_805; // @[executor.scala 473:84]
  wire [7:0] _GEN_1098 = mask_1[0] ? byte_256 : _GEN_806; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1099 = mask_1[1] ? byte_257 : _GEN_807; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1100 = mask_1[2] ? byte_258 : _GEN_808; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1101 = mask_1[3] ? byte_259 : _GEN_809; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1102 = _GEN_4426 == 8'h9 ? _GEN_1098 : _GEN_806; // @[executor.scala 473:84]
  wire [7:0] _GEN_1103 = _GEN_4426 == 8'h9 ? _GEN_1099 : _GEN_807; // @[executor.scala 473:84]
  wire [7:0] _GEN_1104 = _GEN_4426 == 8'h9 ? _GEN_1100 : _GEN_808; // @[executor.scala 473:84]
  wire [7:0] _GEN_1105 = _GEN_4426 == 8'h9 ? _GEN_1101 : _GEN_809; // @[executor.scala 473:84]
  wire [7:0] _GEN_1106 = mask_1[0] ? byte_256 : _GEN_810; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1107 = mask_1[1] ? byte_257 : _GEN_811; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1108 = mask_1[2] ? byte_258 : _GEN_812; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1109 = mask_1[3] ? byte_259 : _GEN_813; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1110 = _GEN_4426 == 8'ha ? _GEN_1106 : _GEN_810; // @[executor.scala 473:84]
  wire [7:0] _GEN_1111 = _GEN_4426 == 8'ha ? _GEN_1107 : _GEN_811; // @[executor.scala 473:84]
  wire [7:0] _GEN_1112 = _GEN_4426 == 8'ha ? _GEN_1108 : _GEN_812; // @[executor.scala 473:84]
  wire [7:0] _GEN_1113 = _GEN_4426 == 8'ha ? _GEN_1109 : _GEN_813; // @[executor.scala 473:84]
  wire [7:0] _GEN_1114 = mask_1[0] ? byte_256 : _GEN_814; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1115 = mask_1[1] ? byte_257 : _GEN_815; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1116 = mask_1[2] ? byte_258 : _GEN_816; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1117 = mask_1[3] ? byte_259 : _GEN_817; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1118 = _GEN_4426 == 8'hb ? _GEN_1114 : _GEN_814; // @[executor.scala 473:84]
  wire [7:0] _GEN_1119 = _GEN_4426 == 8'hb ? _GEN_1115 : _GEN_815; // @[executor.scala 473:84]
  wire [7:0] _GEN_1120 = _GEN_4426 == 8'hb ? _GEN_1116 : _GEN_816; // @[executor.scala 473:84]
  wire [7:0] _GEN_1121 = _GEN_4426 == 8'hb ? _GEN_1117 : _GEN_817; // @[executor.scala 473:84]
  wire [7:0] _GEN_1122 = mask_1[0] ? byte_256 : _GEN_818; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1123 = mask_1[1] ? byte_257 : _GEN_819; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1124 = mask_1[2] ? byte_258 : _GEN_820; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1125 = mask_1[3] ? byte_259 : _GEN_821; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1126 = _GEN_4426 == 8'hc ? _GEN_1122 : _GEN_818; // @[executor.scala 473:84]
  wire [7:0] _GEN_1127 = _GEN_4426 == 8'hc ? _GEN_1123 : _GEN_819; // @[executor.scala 473:84]
  wire [7:0] _GEN_1128 = _GEN_4426 == 8'hc ? _GEN_1124 : _GEN_820; // @[executor.scala 473:84]
  wire [7:0] _GEN_1129 = _GEN_4426 == 8'hc ? _GEN_1125 : _GEN_821; // @[executor.scala 473:84]
  wire [7:0] _GEN_1130 = mask_1[0] ? byte_256 : _GEN_822; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1131 = mask_1[1] ? byte_257 : _GEN_823; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1132 = mask_1[2] ? byte_258 : _GEN_824; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1133 = mask_1[3] ? byte_259 : _GEN_825; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1134 = _GEN_4426 == 8'hd ? _GEN_1130 : _GEN_822; // @[executor.scala 473:84]
  wire [7:0] _GEN_1135 = _GEN_4426 == 8'hd ? _GEN_1131 : _GEN_823; // @[executor.scala 473:84]
  wire [7:0] _GEN_1136 = _GEN_4426 == 8'hd ? _GEN_1132 : _GEN_824; // @[executor.scala 473:84]
  wire [7:0] _GEN_1137 = _GEN_4426 == 8'hd ? _GEN_1133 : _GEN_825; // @[executor.scala 473:84]
  wire [7:0] _GEN_1138 = mask_1[0] ? byte_256 : _GEN_826; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1139 = mask_1[1] ? byte_257 : _GEN_827; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1140 = mask_1[2] ? byte_258 : _GEN_828; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1141 = mask_1[3] ? byte_259 : _GEN_829; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1142 = _GEN_4426 == 8'he ? _GEN_1138 : _GEN_826; // @[executor.scala 473:84]
  wire [7:0] _GEN_1143 = _GEN_4426 == 8'he ? _GEN_1139 : _GEN_827; // @[executor.scala 473:84]
  wire [7:0] _GEN_1144 = _GEN_4426 == 8'he ? _GEN_1140 : _GEN_828; // @[executor.scala 473:84]
  wire [7:0] _GEN_1145 = _GEN_4426 == 8'he ? _GEN_1141 : _GEN_829; // @[executor.scala 473:84]
  wire [7:0] _GEN_1146 = mask_1[0] ? byte_256 : _GEN_830; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1147 = mask_1[1] ? byte_257 : _GEN_831; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1148 = mask_1[2] ? byte_258 : _GEN_832; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1149 = mask_1[3] ? byte_259 : _GEN_833; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1150 = _GEN_4426 == 8'hf ? _GEN_1146 : _GEN_830; // @[executor.scala 473:84]
  wire [7:0] _GEN_1151 = _GEN_4426 == 8'hf ? _GEN_1147 : _GEN_831; // @[executor.scala 473:84]
  wire [7:0] _GEN_1152 = _GEN_4426 == 8'hf ? _GEN_1148 : _GEN_832; // @[executor.scala 473:84]
  wire [7:0] _GEN_1153 = _GEN_4426 == 8'hf ? _GEN_1149 : _GEN_833; // @[executor.scala 473:84]
  wire [7:0] _GEN_1154 = mask_1[0] ? byte_256 : _GEN_834; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1155 = mask_1[1] ? byte_257 : _GEN_835; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1156 = mask_1[2] ? byte_258 : _GEN_836; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1157 = mask_1[3] ? byte_259 : _GEN_837; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1158 = _GEN_4426 == 8'h10 ? _GEN_1154 : _GEN_834; // @[executor.scala 473:84]
  wire [7:0] _GEN_1159 = _GEN_4426 == 8'h10 ? _GEN_1155 : _GEN_835; // @[executor.scala 473:84]
  wire [7:0] _GEN_1160 = _GEN_4426 == 8'h10 ? _GEN_1156 : _GEN_836; // @[executor.scala 473:84]
  wire [7:0] _GEN_1161 = _GEN_4426 == 8'h10 ? _GEN_1157 : _GEN_837; // @[executor.scala 473:84]
  wire [7:0] _GEN_1162 = mask_1[0] ? byte_256 : _GEN_838; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1163 = mask_1[1] ? byte_257 : _GEN_839; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1164 = mask_1[2] ? byte_258 : _GEN_840; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1165 = mask_1[3] ? byte_259 : _GEN_841; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1166 = _GEN_4426 == 8'h11 ? _GEN_1162 : _GEN_838; // @[executor.scala 473:84]
  wire [7:0] _GEN_1167 = _GEN_4426 == 8'h11 ? _GEN_1163 : _GEN_839; // @[executor.scala 473:84]
  wire [7:0] _GEN_1168 = _GEN_4426 == 8'h11 ? _GEN_1164 : _GEN_840; // @[executor.scala 473:84]
  wire [7:0] _GEN_1169 = _GEN_4426 == 8'h11 ? _GEN_1165 : _GEN_841; // @[executor.scala 473:84]
  wire [7:0] _GEN_1170 = mask_1[0] ? byte_256 : _GEN_842; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1171 = mask_1[1] ? byte_257 : _GEN_843; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1172 = mask_1[2] ? byte_258 : _GEN_844; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1173 = mask_1[3] ? byte_259 : _GEN_845; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1174 = _GEN_4426 == 8'h12 ? _GEN_1170 : _GEN_842; // @[executor.scala 473:84]
  wire [7:0] _GEN_1175 = _GEN_4426 == 8'h12 ? _GEN_1171 : _GEN_843; // @[executor.scala 473:84]
  wire [7:0] _GEN_1176 = _GEN_4426 == 8'h12 ? _GEN_1172 : _GEN_844; // @[executor.scala 473:84]
  wire [7:0] _GEN_1177 = _GEN_4426 == 8'h12 ? _GEN_1173 : _GEN_845; // @[executor.scala 473:84]
  wire [7:0] _GEN_1178 = mask_1[0] ? byte_256 : _GEN_846; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1179 = mask_1[1] ? byte_257 : _GEN_847; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1180 = mask_1[2] ? byte_258 : _GEN_848; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1181 = mask_1[3] ? byte_259 : _GEN_849; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1182 = _GEN_4426 == 8'h13 ? _GEN_1178 : _GEN_846; // @[executor.scala 473:84]
  wire [7:0] _GEN_1183 = _GEN_4426 == 8'h13 ? _GEN_1179 : _GEN_847; // @[executor.scala 473:84]
  wire [7:0] _GEN_1184 = _GEN_4426 == 8'h13 ? _GEN_1180 : _GEN_848; // @[executor.scala 473:84]
  wire [7:0] _GEN_1185 = _GEN_4426 == 8'h13 ? _GEN_1181 : _GEN_849; // @[executor.scala 473:84]
  wire [7:0] _GEN_1186 = mask_1[0] ? byte_256 : _GEN_850; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1187 = mask_1[1] ? byte_257 : _GEN_851; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1188 = mask_1[2] ? byte_258 : _GEN_852; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1189 = mask_1[3] ? byte_259 : _GEN_853; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1190 = _GEN_4426 == 8'h14 ? _GEN_1186 : _GEN_850; // @[executor.scala 473:84]
  wire [7:0] _GEN_1191 = _GEN_4426 == 8'h14 ? _GEN_1187 : _GEN_851; // @[executor.scala 473:84]
  wire [7:0] _GEN_1192 = _GEN_4426 == 8'h14 ? _GEN_1188 : _GEN_852; // @[executor.scala 473:84]
  wire [7:0] _GEN_1193 = _GEN_4426 == 8'h14 ? _GEN_1189 : _GEN_853; // @[executor.scala 473:84]
  wire [7:0] _GEN_1194 = mask_1[0] ? byte_256 : _GEN_854; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1195 = mask_1[1] ? byte_257 : _GEN_855; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1196 = mask_1[2] ? byte_258 : _GEN_856; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1197 = mask_1[3] ? byte_259 : _GEN_857; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1198 = _GEN_4426 == 8'h15 ? _GEN_1194 : _GEN_854; // @[executor.scala 473:84]
  wire [7:0] _GEN_1199 = _GEN_4426 == 8'h15 ? _GEN_1195 : _GEN_855; // @[executor.scala 473:84]
  wire [7:0] _GEN_1200 = _GEN_4426 == 8'h15 ? _GEN_1196 : _GEN_856; // @[executor.scala 473:84]
  wire [7:0] _GEN_1201 = _GEN_4426 == 8'h15 ? _GEN_1197 : _GEN_857; // @[executor.scala 473:84]
  wire [7:0] _GEN_1202 = mask_1[0] ? byte_256 : _GEN_858; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1203 = mask_1[1] ? byte_257 : _GEN_859; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1204 = mask_1[2] ? byte_258 : _GEN_860; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1205 = mask_1[3] ? byte_259 : _GEN_861; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1206 = _GEN_4426 == 8'h16 ? _GEN_1202 : _GEN_858; // @[executor.scala 473:84]
  wire [7:0] _GEN_1207 = _GEN_4426 == 8'h16 ? _GEN_1203 : _GEN_859; // @[executor.scala 473:84]
  wire [7:0] _GEN_1208 = _GEN_4426 == 8'h16 ? _GEN_1204 : _GEN_860; // @[executor.scala 473:84]
  wire [7:0] _GEN_1209 = _GEN_4426 == 8'h16 ? _GEN_1205 : _GEN_861; // @[executor.scala 473:84]
  wire [7:0] _GEN_1210 = mask_1[0] ? byte_256 : _GEN_862; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1211 = mask_1[1] ? byte_257 : _GEN_863; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1212 = mask_1[2] ? byte_258 : _GEN_864; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1213 = mask_1[3] ? byte_259 : _GEN_865; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1214 = _GEN_4426 == 8'h17 ? _GEN_1210 : _GEN_862; // @[executor.scala 473:84]
  wire [7:0] _GEN_1215 = _GEN_4426 == 8'h17 ? _GEN_1211 : _GEN_863; // @[executor.scala 473:84]
  wire [7:0] _GEN_1216 = _GEN_4426 == 8'h17 ? _GEN_1212 : _GEN_864; // @[executor.scala 473:84]
  wire [7:0] _GEN_1217 = _GEN_4426 == 8'h17 ? _GEN_1213 : _GEN_865; // @[executor.scala 473:84]
  wire [7:0] _GEN_1218 = mask_1[0] ? byte_256 : _GEN_866; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1219 = mask_1[1] ? byte_257 : _GEN_867; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1220 = mask_1[2] ? byte_258 : _GEN_868; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1221 = mask_1[3] ? byte_259 : _GEN_869; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1222 = _GEN_4426 == 8'h18 ? _GEN_1218 : _GEN_866; // @[executor.scala 473:84]
  wire [7:0] _GEN_1223 = _GEN_4426 == 8'h18 ? _GEN_1219 : _GEN_867; // @[executor.scala 473:84]
  wire [7:0] _GEN_1224 = _GEN_4426 == 8'h18 ? _GEN_1220 : _GEN_868; // @[executor.scala 473:84]
  wire [7:0] _GEN_1225 = _GEN_4426 == 8'h18 ? _GEN_1221 : _GEN_869; // @[executor.scala 473:84]
  wire [7:0] _GEN_1226 = mask_1[0] ? byte_256 : _GEN_870; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1227 = mask_1[1] ? byte_257 : _GEN_871; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1228 = mask_1[2] ? byte_258 : _GEN_872; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1229 = mask_1[3] ? byte_259 : _GEN_873; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1230 = _GEN_4426 == 8'h19 ? _GEN_1226 : _GEN_870; // @[executor.scala 473:84]
  wire [7:0] _GEN_1231 = _GEN_4426 == 8'h19 ? _GEN_1227 : _GEN_871; // @[executor.scala 473:84]
  wire [7:0] _GEN_1232 = _GEN_4426 == 8'h19 ? _GEN_1228 : _GEN_872; // @[executor.scala 473:84]
  wire [7:0] _GEN_1233 = _GEN_4426 == 8'h19 ? _GEN_1229 : _GEN_873; // @[executor.scala 473:84]
  wire [7:0] _GEN_1234 = mask_1[0] ? byte_256 : _GEN_874; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1235 = mask_1[1] ? byte_257 : _GEN_875; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1236 = mask_1[2] ? byte_258 : _GEN_876; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1237 = mask_1[3] ? byte_259 : _GEN_877; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1238 = _GEN_4426 == 8'h1a ? _GEN_1234 : _GEN_874; // @[executor.scala 473:84]
  wire [7:0] _GEN_1239 = _GEN_4426 == 8'h1a ? _GEN_1235 : _GEN_875; // @[executor.scala 473:84]
  wire [7:0] _GEN_1240 = _GEN_4426 == 8'h1a ? _GEN_1236 : _GEN_876; // @[executor.scala 473:84]
  wire [7:0] _GEN_1241 = _GEN_4426 == 8'h1a ? _GEN_1237 : _GEN_877; // @[executor.scala 473:84]
  wire [7:0] _GEN_1242 = mask_1[0] ? byte_256 : _GEN_878; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1243 = mask_1[1] ? byte_257 : _GEN_879; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1244 = mask_1[2] ? byte_258 : _GEN_880; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1245 = mask_1[3] ? byte_259 : _GEN_881; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1246 = _GEN_4426 == 8'h1b ? _GEN_1242 : _GEN_878; // @[executor.scala 473:84]
  wire [7:0] _GEN_1247 = _GEN_4426 == 8'h1b ? _GEN_1243 : _GEN_879; // @[executor.scala 473:84]
  wire [7:0] _GEN_1248 = _GEN_4426 == 8'h1b ? _GEN_1244 : _GEN_880; // @[executor.scala 473:84]
  wire [7:0] _GEN_1249 = _GEN_4426 == 8'h1b ? _GEN_1245 : _GEN_881; // @[executor.scala 473:84]
  wire [7:0] _GEN_1250 = mask_1[0] ? byte_256 : _GEN_882; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1251 = mask_1[1] ? byte_257 : _GEN_883; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1252 = mask_1[2] ? byte_258 : _GEN_884; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1253 = mask_1[3] ? byte_259 : _GEN_885; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1254 = _GEN_4426 == 8'h1c ? _GEN_1250 : _GEN_882; // @[executor.scala 473:84]
  wire [7:0] _GEN_1255 = _GEN_4426 == 8'h1c ? _GEN_1251 : _GEN_883; // @[executor.scala 473:84]
  wire [7:0] _GEN_1256 = _GEN_4426 == 8'h1c ? _GEN_1252 : _GEN_884; // @[executor.scala 473:84]
  wire [7:0] _GEN_1257 = _GEN_4426 == 8'h1c ? _GEN_1253 : _GEN_885; // @[executor.scala 473:84]
  wire [7:0] _GEN_1258 = mask_1[0] ? byte_256 : _GEN_886; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1259 = mask_1[1] ? byte_257 : _GEN_887; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1260 = mask_1[2] ? byte_258 : _GEN_888; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1261 = mask_1[3] ? byte_259 : _GEN_889; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1262 = _GEN_4426 == 8'h1d ? _GEN_1258 : _GEN_886; // @[executor.scala 473:84]
  wire [7:0] _GEN_1263 = _GEN_4426 == 8'h1d ? _GEN_1259 : _GEN_887; // @[executor.scala 473:84]
  wire [7:0] _GEN_1264 = _GEN_4426 == 8'h1d ? _GEN_1260 : _GEN_888; // @[executor.scala 473:84]
  wire [7:0] _GEN_1265 = _GEN_4426 == 8'h1d ? _GEN_1261 : _GEN_889; // @[executor.scala 473:84]
  wire [7:0] _GEN_1266 = mask_1[0] ? byte_256 : _GEN_890; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1267 = mask_1[1] ? byte_257 : _GEN_891; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1268 = mask_1[2] ? byte_258 : _GEN_892; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1269 = mask_1[3] ? byte_259 : _GEN_893; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1270 = _GEN_4426 == 8'h1e ? _GEN_1266 : _GEN_890; // @[executor.scala 473:84]
  wire [7:0] _GEN_1271 = _GEN_4426 == 8'h1e ? _GEN_1267 : _GEN_891; // @[executor.scala 473:84]
  wire [7:0] _GEN_1272 = _GEN_4426 == 8'h1e ? _GEN_1268 : _GEN_892; // @[executor.scala 473:84]
  wire [7:0] _GEN_1273 = _GEN_4426 == 8'h1e ? _GEN_1269 : _GEN_893; // @[executor.scala 473:84]
  wire [7:0] _GEN_1274 = mask_1[0] ? byte_256 : _GEN_894; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1275 = mask_1[1] ? byte_257 : _GEN_895; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1276 = mask_1[2] ? byte_258 : _GEN_896; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1277 = mask_1[3] ? byte_259 : _GEN_897; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1278 = _GEN_4426 == 8'h1f ? _GEN_1274 : _GEN_894; // @[executor.scala 473:84]
  wire [7:0] _GEN_1279 = _GEN_4426 == 8'h1f ? _GEN_1275 : _GEN_895; // @[executor.scala 473:84]
  wire [7:0] _GEN_1280 = _GEN_4426 == 8'h1f ? _GEN_1276 : _GEN_896; // @[executor.scala 473:84]
  wire [7:0] _GEN_1281 = _GEN_4426 == 8'h1f ? _GEN_1277 : _GEN_897; // @[executor.scala 473:84]
  wire [7:0] _GEN_1282 = mask_1[0] ? byte_256 : _GEN_898; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1283 = mask_1[1] ? byte_257 : _GEN_899; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1284 = mask_1[2] ? byte_258 : _GEN_900; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1285 = mask_1[3] ? byte_259 : _GEN_901; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1286 = _GEN_4426 == 8'h20 ? _GEN_1282 : _GEN_898; // @[executor.scala 473:84]
  wire [7:0] _GEN_1287 = _GEN_4426 == 8'h20 ? _GEN_1283 : _GEN_899; // @[executor.scala 473:84]
  wire [7:0] _GEN_1288 = _GEN_4426 == 8'h20 ? _GEN_1284 : _GEN_900; // @[executor.scala 473:84]
  wire [7:0] _GEN_1289 = _GEN_4426 == 8'h20 ? _GEN_1285 : _GEN_901; // @[executor.scala 473:84]
  wire [7:0] _GEN_1290 = mask_1[0] ? byte_256 : _GEN_902; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1291 = mask_1[1] ? byte_257 : _GEN_903; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1292 = mask_1[2] ? byte_258 : _GEN_904; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1293 = mask_1[3] ? byte_259 : _GEN_905; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1294 = _GEN_4426 == 8'h21 ? _GEN_1290 : _GEN_902; // @[executor.scala 473:84]
  wire [7:0] _GEN_1295 = _GEN_4426 == 8'h21 ? _GEN_1291 : _GEN_903; // @[executor.scala 473:84]
  wire [7:0] _GEN_1296 = _GEN_4426 == 8'h21 ? _GEN_1292 : _GEN_904; // @[executor.scala 473:84]
  wire [7:0] _GEN_1297 = _GEN_4426 == 8'h21 ? _GEN_1293 : _GEN_905; // @[executor.scala 473:84]
  wire [7:0] _GEN_1298 = mask_1[0] ? byte_256 : _GEN_906; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1299 = mask_1[1] ? byte_257 : _GEN_907; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1300 = mask_1[2] ? byte_258 : _GEN_908; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1301 = mask_1[3] ? byte_259 : _GEN_909; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1302 = _GEN_4426 == 8'h22 ? _GEN_1298 : _GEN_906; // @[executor.scala 473:84]
  wire [7:0] _GEN_1303 = _GEN_4426 == 8'h22 ? _GEN_1299 : _GEN_907; // @[executor.scala 473:84]
  wire [7:0] _GEN_1304 = _GEN_4426 == 8'h22 ? _GEN_1300 : _GEN_908; // @[executor.scala 473:84]
  wire [7:0] _GEN_1305 = _GEN_4426 == 8'h22 ? _GEN_1301 : _GEN_909; // @[executor.scala 473:84]
  wire [7:0] _GEN_1306 = mask_1[0] ? byte_256 : _GEN_910; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1307 = mask_1[1] ? byte_257 : _GEN_911; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1308 = mask_1[2] ? byte_258 : _GEN_912; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1309 = mask_1[3] ? byte_259 : _GEN_913; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1310 = _GEN_4426 == 8'h23 ? _GEN_1306 : _GEN_910; // @[executor.scala 473:84]
  wire [7:0] _GEN_1311 = _GEN_4426 == 8'h23 ? _GEN_1307 : _GEN_911; // @[executor.scala 473:84]
  wire [7:0] _GEN_1312 = _GEN_4426 == 8'h23 ? _GEN_1308 : _GEN_912; // @[executor.scala 473:84]
  wire [7:0] _GEN_1313 = _GEN_4426 == 8'h23 ? _GEN_1309 : _GEN_913; // @[executor.scala 473:84]
  wire [7:0] _GEN_1314 = mask_1[0] ? byte_256 : _GEN_914; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1315 = mask_1[1] ? byte_257 : _GEN_915; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1316 = mask_1[2] ? byte_258 : _GEN_916; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1317 = mask_1[3] ? byte_259 : _GEN_917; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1318 = _GEN_4426 == 8'h24 ? _GEN_1314 : _GEN_914; // @[executor.scala 473:84]
  wire [7:0] _GEN_1319 = _GEN_4426 == 8'h24 ? _GEN_1315 : _GEN_915; // @[executor.scala 473:84]
  wire [7:0] _GEN_1320 = _GEN_4426 == 8'h24 ? _GEN_1316 : _GEN_916; // @[executor.scala 473:84]
  wire [7:0] _GEN_1321 = _GEN_4426 == 8'h24 ? _GEN_1317 : _GEN_917; // @[executor.scala 473:84]
  wire [7:0] _GEN_1322 = mask_1[0] ? byte_256 : _GEN_918; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1323 = mask_1[1] ? byte_257 : _GEN_919; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1324 = mask_1[2] ? byte_258 : _GEN_920; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1325 = mask_1[3] ? byte_259 : _GEN_921; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1326 = _GEN_4426 == 8'h25 ? _GEN_1322 : _GEN_918; // @[executor.scala 473:84]
  wire [7:0] _GEN_1327 = _GEN_4426 == 8'h25 ? _GEN_1323 : _GEN_919; // @[executor.scala 473:84]
  wire [7:0] _GEN_1328 = _GEN_4426 == 8'h25 ? _GEN_1324 : _GEN_920; // @[executor.scala 473:84]
  wire [7:0] _GEN_1329 = _GEN_4426 == 8'h25 ? _GEN_1325 : _GEN_921; // @[executor.scala 473:84]
  wire [7:0] _GEN_1330 = mask_1[0] ? byte_256 : _GEN_922; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1331 = mask_1[1] ? byte_257 : _GEN_923; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1332 = mask_1[2] ? byte_258 : _GEN_924; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1333 = mask_1[3] ? byte_259 : _GEN_925; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1334 = _GEN_4426 == 8'h26 ? _GEN_1330 : _GEN_922; // @[executor.scala 473:84]
  wire [7:0] _GEN_1335 = _GEN_4426 == 8'h26 ? _GEN_1331 : _GEN_923; // @[executor.scala 473:84]
  wire [7:0] _GEN_1336 = _GEN_4426 == 8'h26 ? _GEN_1332 : _GEN_924; // @[executor.scala 473:84]
  wire [7:0] _GEN_1337 = _GEN_4426 == 8'h26 ? _GEN_1333 : _GEN_925; // @[executor.scala 473:84]
  wire [7:0] _GEN_1338 = mask_1[0] ? byte_256 : _GEN_926; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1339 = mask_1[1] ? byte_257 : _GEN_927; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1340 = mask_1[2] ? byte_258 : _GEN_928; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1341 = mask_1[3] ? byte_259 : _GEN_929; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1342 = _GEN_4426 == 8'h27 ? _GEN_1338 : _GEN_926; // @[executor.scala 473:84]
  wire [7:0] _GEN_1343 = _GEN_4426 == 8'h27 ? _GEN_1339 : _GEN_927; // @[executor.scala 473:84]
  wire [7:0] _GEN_1344 = _GEN_4426 == 8'h27 ? _GEN_1340 : _GEN_928; // @[executor.scala 473:84]
  wire [7:0] _GEN_1345 = _GEN_4426 == 8'h27 ? _GEN_1341 : _GEN_929; // @[executor.scala 473:84]
  wire [7:0] _GEN_1346 = mask_1[0] ? byte_256 : _GEN_930; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1347 = mask_1[1] ? byte_257 : _GEN_931; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1348 = mask_1[2] ? byte_258 : _GEN_932; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1349 = mask_1[3] ? byte_259 : _GEN_933; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1350 = _GEN_4426 == 8'h28 ? _GEN_1346 : _GEN_930; // @[executor.scala 473:84]
  wire [7:0] _GEN_1351 = _GEN_4426 == 8'h28 ? _GEN_1347 : _GEN_931; // @[executor.scala 473:84]
  wire [7:0] _GEN_1352 = _GEN_4426 == 8'h28 ? _GEN_1348 : _GEN_932; // @[executor.scala 473:84]
  wire [7:0] _GEN_1353 = _GEN_4426 == 8'h28 ? _GEN_1349 : _GEN_933; // @[executor.scala 473:84]
  wire [7:0] _GEN_1354 = mask_1[0] ? byte_256 : _GEN_934; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1355 = mask_1[1] ? byte_257 : _GEN_935; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1356 = mask_1[2] ? byte_258 : _GEN_936; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1357 = mask_1[3] ? byte_259 : _GEN_937; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1358 = _GEN_4426 == 8'h29 ? _GEN_1354 : _GEN_934; // @[executor.scala 473:84]
  wire [7:0] _GEN_1359 = _GEN_4426 == 8'h29 ? _GEN_1355 : _GEN_935; // @[executor.scala 473:84]
  wire [7:0] _GEN_1360 = _GEN_4426 == 8'h29 ? _GEN_1356 : _GEN_936; // @[executor.scala 473:84]
  wire [7:0] _GEN_1361 = _GEN_4426 == 8'h29 ? _GEN_1357 : _GEN_937; // @[executor.scala 473:84]
  wire [7:0] _GEN_1362 = mask_1[0] ? byte_256 : _GEN_938; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1363 = mask_1[1] ? byte_257 : _GEN_939; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1364 = mask_1[2] ? byte_258 : _GEN_940; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1365 = mask_1[3] ? byte_259 : _GEN_941; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1366 = _GEN_4426 == 8'h2a ? _GEN_1362 : _GEN_938; // @[executor.scala 473:84]
  wire [7:0] _GEN_1367 = _GEN_4426 == 8'h2a ? _GEN_1363 : _GEN_939; // @[executor.scala 473:84]
  wire [7:0] _GEN_1368 = _GEN_4426 == 8'h2a ? _GEN_1364 : _GEN_940; // @[executor.scala 473:84]
  wire [7:0] _GEN_1369 = _GEN_4426 == 8'h2a ? _GEN_1365 : _GEN_941; // @[executor.scala 473:84]
  wire [7:0] _GEN_1370 = mask_1[0] ? byte_256 : _GEN_942; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1371 = mask_1[1] ? byte_257 : _GEN_943; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1372 = mask_1[2] ? byte_258 : _GEN_944; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1373 = mask_1[3] ? byte_259 : _GEN_945; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1374 = _GEN_4426 == 8'h2b ? _GEN_1370 : _GEN_942; // @[executor.scala 473:84]
  wire [7:0] _GEN_1375 = _GEN_4426 == 8'h2b ? _GEN_1371 : _GEN_943; // @[executor.scala 473:84]
  wire [7:0] _GEN_1376 = _GEN_4426 == 8'h2b ? _GEN_1372 : _GEN_944; // @[executor.scala 473:84]
  wire [7:0] _GEN_1377 = _GEN_4426 == 8'h2b ? _GEN_1373 : _GEN_945; // @[executor.scala 473:84]
  wire [7:0] _GEN_1378 = mask_1[0] ? byte_256 : _GEN_946; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1379 = mask_1[1] ? byte_257 : _GEN_947; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1380 = mask_1[2] ? byte_258 : _GEN_948; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1381 = mask_1[3] ? byte_259 : _GEN_949; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1382 = _GEN_4426 == 8'h2c ? _GEN_1378 : _GEN_946; // @[executor.scala 473:84]
  wire [7:0] _GEN_1383 = _GEN_4426 == 8'h2c ? _GEN_1379 : _GEN_947; // @[executor.scala 473:84]
  wire [7:0] _GEN_1384 = _GEN_4426 == 8'h2c ? _GEN_1380 : _GEN_948; // @[executor.scala 473:84]
  wire [7:0] _GEN_1385 = _GEN_4426 == 8'h2c ? _GEN_1381 : _GEN_949; // @[executor.scala 473:84]
  wire [7:0] _GEN_1386 = mask_1[0] ? byte_256 : _GEN_950; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1387 = mask_1[1] ? byte_257 : _GEN_951; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1388 = mask_1[2] ? byte_258 : _GEN_952; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1389 = mask_1[3] ? byte_259 : _GEN_953; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1390 = _GEN_4426 == 8'h2d ? _GEN_1386 : _GEN_950; // @[executor.scala 473:84]
  wire [7:0] _GEN_1391 = _GEN_4426 == 8'h2d ? _GEN_1387 : _GEN_951; // @[executor.scala 473:84]
  wire [7:0] _GEN_1392 = _GEN_4426 == 8'h2d ? _GEN_1388 : _GEN_952; // @[executor.scala 473:84]
  wire [7:0] _GEN_1393 = _GEN_4426 == 8'h2d ? _GEN_1389 : _GEN_953; // @[executor.scala 473:84]
  wire [7:0] _GEN_1394 = mask_1[0] ? byte_256 : _GEN_954; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1395 = mask_1[1] ? byte_257 : _GEN_955; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1396 = mask_1[2] ? byte_258 : _GEN_956; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1397 = mask_1[3] ? byte_259 : _GEN_957; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1398 = _GEN_4426 == 8'h2e ? _GEN_1394 : _GEN_954; // @[executor.scala 473:84]
  wire [7:0] _GEN_1399 = _GEN_4426 == 8'h2e ? _GEN_1395 : _GEN_955; // @[executor.scala 473:84]
  wire [7:0] _GEN_1400 = _GEN_4426 == 8'h2e ? _GEN_1396 : _GEN_956; // @[executor.scala 473:84]
  wire [7:0] _GEN_1401 = _GEN_4426 == 8'h2e ? _GEN_1397 : _GEN_957; // @[executor.scala 473:84]
  wire [7:0] _GEN_1402 = mask_1[0] ? byte_256 : _GEN_958; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1403 = mask_1[1] ? byte_257 : _GEN_959; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1404 = mask_1[2] ? byte_258 : _GEN_960; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1405 = mask_1[3] ? byte_259 : _GEN_961; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1406 = _GEN_4426 == 8'h2f ? _GEN_1402 : _GEN_958; // @[executor.scala 473:84]
  wire [7:0] _GEN_1407 = _GEN_4426 == 8'h2f ? _GEN_1403 : _GEN_959; // @[executor.scala 473:84]
  wire [7:0] _GEN_1408 = _GEN_4426 == 8'h2f ? _GEN_1404 : _GEN_960; // @[executor.scala 473:84]
  wire [7:0] _GEN_1409 = _GEN_4426 == 8'h2f ? _GEN_1405 : _GEN_961; // @[executor.scala 473:84]
  wire [7:0] _GEN_1410 = mask_1[0] ? byte_256 : _GEN_962; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1411 = mask_1[1] ? byte_257 : _GEN_963; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1412 = mask_1[2] ? byte_258 : _GEN_964; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1413 = mask_1[3] ? byte_259 : _GEN_965; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1414 = _GEN_4426 == 8'h30 ? _GEN_1410 : _GEN_962; // @[executor.scala 473:84]
  wire [7:0] _GEN_1415 = _GEN_4426 == 8'h30 ? _GEN_1411 : _GEN_963; // @[executor.scala 473:84]
  wire [7:0] _GEN_1416 = _GEN_4426 == 8'h30 ? _GEN_1412 : _GEN_964; // @[executor.scala 473:84]
  wire [7:0] _GEN_1417 = _GEN_4426 == 8'h30 ? _GEN_1413 : _GEN_965; // @[executor.scala 473:84]
  wire [7:0] _GEN_1418 = mask_1[0] ? byte_256 : _GEN_966; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1419 = mask_1[1] ? byte_257 : _GEN_967; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1420 = mask_1[2] ? byte_258 : _GEN_968; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1421 = mask_1[3] ? byte_259 : _GEN_969; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1422 = _GEN_4426 == 8'h31 ? _GEN_1418 : _GEN_966; // @[executor.scala 473:84]
  wire [7:0] _GEN_1423 = _GEN_4426 == 8'h31 ? _GEN_1419 : _GEN_967; // @[executor.scala 473:84]
  wire [7:0] _GEN_1424 = _GEN_4426 == 8'h31 ? _GEN_1420 : _GEN_968; // @[executor.scala 473:84]
  wire [7:0] _GEN_1425 = _GEN_4426 == 8'h31 ? _GEN_1421 : _GEN_969; // @[executor.scala 473:84]
  wire [7:0] _GEN_1426 = mask_1[0] ? byte_256 : _GEN_970; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1427 = mask_1[1] ? byte_257 : _GEN_971; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1428 = mask_1[2] ? byte_258 : _GEN_972; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1429 = mask_1[3] ? byte_259 : _GEN_973; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1430 = _GEN_4426 == 8'h32 ? _GEN_1426 : _GEN_970; // @[executor.scala 473:84]
  wire [7:0] _GEN_1431 = _GEN_4426 == 8'h32 ? _GEN_1427 : _GEN_971; // @[executor.scala 473:84]
  wire [7:0] _GEN_1432 = _GEN_4426 == 8'h32 ? _GEN_1428 : _GEN_972; // @[executor.scala 473:84]
  wire [7:0] _GEN_1433 = _GEN_4426 == 8'h32 ? _GEN_1429 : _GEN_973; // @[executor.scala 473:84]
  wire [7:0] _GEN_1434 = mask_1[0] ? byte_256 : _GEN_974; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1435 = mask_1[1] ? byte_257 : _GEN_975; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1436 = mask_1[2] ? byte_258 : _GEN_976; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1437 = mask_1[3] ? byte_259 : _GEN_977; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1438 = _GEN_4426 == 8'h33 ? _GEN_1434 : _GEN_974; // @[executor.scala 473:84]
  wire [7:0] _GEN_1439 = _GEN_4426 == 8'h33 ? _GEN_1435 : _GEN_975; // @[executor.scala 473:84]
  wire [7:0] _GEN_1440 = _GEN_4426 == 8'h33 ? _GEN_1436 : _GEN_976; // @[executor.scala 473:84]
  wire [7:0] _GEN_1441 = _GEN_4426 == 8'h33 ? _GEN_1437 : _GEN_977; // @[executor.scala 473:84]
  wire [7:0] _GEN_1442 = mask_1[0] ? byte_256 : _GEN_978; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1443 = mask_1[1] ? byte_257 : _GEN_979; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1444 = mask_1[2] ? byte_258 : _GEN_980; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1445 = mask_1[3] ? byte_259 : _GEN_981; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1446 = _GEN_4426 == 8'h34 ? _GEN_1442 : _GEN_978; // @[executor.scala 473:84]
  wire [7:0] _GEN_1447 = _GEN_4426 == 8'h34 ? _GEN_1443 : _GEN_979; // @[executor.scala 473:84]
  wire [7:0] _GEN_1448 = _GEN_4426 == 8'h34 ? _GEN_1444 : _GEN_980; // @[executor.scala 473:84]
  wire [7:0] _GEN_1449 = _GEN_4426 == 8'h34 ? _GEN_1445 : _GEN_981; // @[executor.scala 473:84]
  wire [7:0] _GEN_1450 = mask_1[0] ? byte_256 : _GEN_982; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1451 = mask_1[1] ? byte_257 : _GEN_983; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1452 = mask_1[2] ? byte_258 : _GEN_984; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1453 = mask_1[3] ? byte_259 : _GEN_985; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1454 = _GEN_4426 == 8'h35 ? _GEN_1450 : _GEN_982; // @[executor.scala 473:84]
  wire [7:0] _GEN_1455 = _GEN_4426 == 8'h35 ? _GEN_1451 : _GEN_983; // @[executor.scala 473:84]
  wire [7:0] _GEN_1456 = _GEN_4426 == 8'h35 ? _GEN_1452 : _GEN_984; // @[executor.scala 473:84]
  wire [7:0] _GEN_1457 = _GEN_4426 == 8'h35 ? _GEN_1453 : _GEN_985; // @[executor.scala 473:84]
  wire [7:0] _GEN_1458 = mask_1[0] ? byte_256 : _GEN_986; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1459 = mask_1[1] ? byte_257 : _GEN_987; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1460 = mask_1[2] ? byte_258 : _GEN_988; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1461 = mask_1[3] ? byte_259 : _GEN_989; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1462 = _GEN_4426 == 8'h36 ? _GEN_1458 : _GEN_986; // @[executor.scala 473:84]
  wire [7:0] _GEN_1463 = _GEN_4426 == 8'h36 ? _GEN_1459 : _GEN_987; // @[executor.scala 473:84]
  wire [7:0] _GEN_1464 = _GEN_4426 == 8'h36 ? _GEN_1460 : _GEN_988; // @[executor.scala 473:84]
  wire [7:0] _GEN_1465 = _GEN_4426 == 8'h36 ? _GEN_1461 : _GEN_989; // @[executor.scala 473:84]
  wire [7:0] _GEN_1466 = mask_1[0] ? byte_256 : _GEN_990; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1467 = mask_1[1] ? byte_257 : _GEN_991; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1468 = mask_1[2] ? byte_258 : _GEN_992; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1469 = mask_1[3] ? byte_259 : _GEN_993; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1470 = _GEN_4426 == 8'h37 ? _GEN_1466 : _GEN_990; // @[executor.scala 473:84]
  wire [7:0] _GEN_1471 = _GEN_4426 == 8'h37 ? _GEN_1467 : _GEN_991; // @[executor.scala 473:84]
  wire [7:0] _GEN_1472 = _GEN_4426 == 8'h37 ? _GEN_1468 : _GEN_992; // @[executor.scala 473:84]
  wire [7:0] _GEN_1473 = _GEN_4426 == 8'h37 ? _GEN_1469 : _GEN_993; // @[executor.scala 473:84]
  wire [7:0] _GEN_1474 = mask_1[0] ? byte_256 : _GEN_994; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1475 = mask_1[1] ? byte_257 : _GEN_995; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1476 = mask_1[2] ? byte_258 : _GEN_996; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1477 = mask_1[3] ? byte_259 : _GEN_997; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1478 = _GEN_4426 == 8'h38 ? _GEN_1474 : _GEN_994; // @[executor.scala 473:84]
  wire [7:0] _GEN_1479 = _GEN_4426 == 8'h38 ? _GEN_1475 : _GEN_995; // @[executor.scala 473:84]
  wire [7:0] _GEN_1480 = _GEN_4426 == 8'h38 ? _GEN_1476 : _GEN_996; // @[executor.scala 473:84]
  wire [7:0] _GEN_1481 = _GEN_4426 == 8'h38 ? _GEN_1477 : _GEN_997; // @[executor.scala 473:84]
  wire [7:0] _GEN_1482 = mask_1[0] ? byte_256 : _GEN_998; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1483 = mask_1[1] ? byte_257 : _GEN_999; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1484 = mask_1[2] ? byte_258 : _GEN_1000; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1485 = mask_1[3] ? byte_259 : _GEN_1001; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1486 = _GEN_4426 == 8'h39 ? _GEN_1482 : _GEN_998; // @[executor.scala 473:84]
  wire [7:0] _GEN_1487 = _GEN_4426 == 8'h39 ? _GEN_1483 : _GEN_999; // @[executor.scala 473:84]
  wire [7:0] _GEN_1488 = _GEN_4426 == 8'h39 ? _GEN_1484 : _GEN_1000; // @[executor.scala 473:84]
  wire [7:0] _GEN_1489 = _GEN_4426 == 8'h39 ? _GEN_1485 : _GEN_1001; // @[executor.scala 473:84]
  wire [7:0] _GEN_1490 = mask_1[0] ? byte_256 : _GEN_1002; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1491 = mask_1[1] ? byte_257 : _GEN_1003; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1492 = mask_1[2] ? byte_258 : _GEN_1004; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1493 = mask_1[3] ? byte_259 : _GEN_1005; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1494 = _GEN_4426 == 8'h3a ? _GEN_1490 : _GEN_1002; // @[executor.scala 473:84]
  wire [7:0] _GEN_1495 = _GEN_4426 == 8'h3a ? _GEN_1491 : _GEN_1003; // @[executor.scala 473:84]
  wire [7:0] _GEN_1496 = _GEN_4426 == 8'h3a ? _GEN_1492 : _GEN_1004; // @[executor.scala 473:84]
  wire [7:0] _GEN_1497 = _GEN_4426 == 8'h3a ? _GEN_1493 : _GEN_1005; // @[executor.scala 473:84]
  wire [7:0] _GEN_1498 = mask_1[0] ? byte_256 : _GEN_1006; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1499 = mask_1[1] ? byte_257 : _GEN_1007; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1500 = mask_1[2] ? byte_258 : _GEN_1008; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1501 = mask_1[3] ? byte_259 : _GEN_1009; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1502 = _GEN_4426 == 8'h3b ? _GEN_1498 : _GEN_1006; // @[executor.scala 473:84]
  wire [7:0] _GEN_1503 = _GEN_4426 == 8'h3b ? _GEN_1499 : _GEN_1007; // @[executor.scala 473:84]
  wire [7:0] _GEN_1504 = _GEN_4426 == 8'h3b ? _GEN_1500 : _GEN_1008; // @[executor.scala 473:84]
  wire [7:0] _GEN_1505 = _GEN_4426 == 8'h3b ? _GEN_1501 : _GEN_1009; // @[executor.scala 473:84]
  wire [7:0] _GEN_1506 = mask_1[0] ? byte_256 : _GEN_1010; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1507 = mask_1[1] ? byte_257 : _GEN_1011; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1508 = mask_1[2] ? byte_258 : _GEN_1012; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1509 = mask_1[3] ? byte_259 : _GEN_1013; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1510 = _GEN_4426 == 8'h3c ? _GEN_1506 : _GEN_1010; // @[executor.scala 473:84]
  wire [7:0] _GEN_1511 = _GEN_4426 == 8'h3c ? _GEN_1507 : _GEN_1011; // @[executor.scala 473:84]
  wire [7:0] _GEN_1512 = _GEN_4426 == 8'h3c ? _GEN_1508 : _GEN_1012; // @[executor.scala 473:84]
  wire [7:0] _GEN_1513 = _GEN_4426 == 8'h3c ? _GEN_1509 : _GEN_1013; // @[executor.scala 473:84]
  wire [7:0] _GEN_1514 = mask_1[0] ? byte_256 : _GEN_1014; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1515 = mask_1[1] ? byte_257 : _GEN_1015; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1516 = mask_1[2] ? byte_258 : _GEN_1016; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1517 = mask_1[3] ? byte_259 : _GEN_1017; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1518 = _GEN_4426 == 8'h3d ? _GEN_1514 : _GEN_1014; // @[executor.scala 473:84]
  wire [7:0] _GEN_1519 = _GEN_4426 == 8'h3d ? _GEN_1515 : _GEN_1015; // @[executor.scala 473:84]
  wire [7:0] _GEN_1520 = _GEN_4426 == 8'h3d ? _GEN_1516 : _GEN_1016; // @[executor.scala 473:84]
  wire [7:0] _GEN_1521 = _GEN_4426 == 8'h3d ? _GEN_1517 : _GEN_1017; // @[executor.scala 473:84]
  wire [7:0] _GEN_1522 = mask_1[0] ? byte_256 : _GEN_1018; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1523 = mask_1[1] ? byte_257 : _GEN_1019; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1524 = mask_1[2] ? byte_258 : _GEN_1020; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1525 = mask_1[3] ? byte_259 : _GEN_1021; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1526 = _GEN_4426 == 8'h3e ? _GEN_1522 : _GEN_1018; // @[executor.scala 473:84]
  wire [7:0] _GEN_1527 = _GEN_4426 == 8'h3e ? _GEN_1523 : _GEN_1019; // @[executor.scala 473:84]
  wire [7:0] _GEN_1528 = _GEN_4426 == 8'h3e ? _GEN_1524 : _GEN_1020; // @[executor.scala 473:84]
  wire [7:0] _GEN_1529 = _GEN_4426 == 8'h3e ? _GEN_1525 : _GEN_1021; // @[executor.scala 473:84]
  wire [7:0] _GEN_1530 = mask_1[0] ? byte_256 : _GEN_1022; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1531 = mask_1[1] ? byte_257 : _GEN_1023; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1532 = mask_1[2] ? byte_258 : _GEN_1024; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1533 = mask_1[3] ? byte_259 : _GEN_1025; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1534 = _GEN_4426 == 8'h3f ? _GEN_1530 : _GEN_1022; // @[executor.scala 473:84]
  wire [7:0] _GEN_1535 = _GEN_4426 == 8'h3f ? _GEN_1531 : _GEN_1023; // @[executor.scala 473:84]
  wire [7:0] _GEN_1536 = _GEN_4426 == 8'h3f ? _GEN_1532 : _GEN_1024; // @[executor.scala 473:84]
  wire [7:0] _GEN_1537 = _GEN_4426 == 8'h3f ? _GEN_1533 : _GEN_1025; // @[executor.scala 473:84]
  wire [7:0] _GEN_1538 = opcode_1 != 4'h0 ? _GEN_1030 : _GEN_770; // @[executor.scala 470:55]
  wire [7:0] _GEN_1539 = opcode_1 != 4'h0 ? _GEN_1031 : _GEN_771; // @[executor.scala 470:55]
  wire [7:0] _GEN_1540 = opcode_1 != 4'h0 ? _GEN_1032 : _GEN_772; // @[executor.scala 470:55]
  wire [7:0] _GEN_1541 = opcode_1 != 4'h0 ? _GEN_1033 : _GEN_773; // @[executor.scala 470:55]
  wire [7:0] _GEN_1542 = opcode_1 != 4'h0 ? _GEN_1038 : _GEN_774; // @[executor.scala 470:55]
  wire [7:0] _GEN_1543 = opcode_1 != 4'h0 ? _GEN_1039 : _GEN_775; // @[executor.scala 470:55]
  wire [7:0] _GEN_1544 = opcode_1 != 4'h0 ? _GEN_1040 : _GEN_776; // @[executor.scala 470:55]
  wire [7:0] _GEN_1545 = opcode_1 != 4'h0 ? _GEN_1041 : _GEN_777; // @[executor.scala 470:55]
  wire [7:0] _GEN_1546 = opcode_1 != 4'h0 ? _GEN_1046 : _GEN_778; // @[executor.scala 470:55]
  wire [7:0] _GEN_1547 = opcode_1 != 4'h0 ? _GEN_1047 : _GEN_779; // @[executor.scala 470:55]
  wire [7:0] _GEN_1548 = opcode_1 != 4'h0 ? _GEN_1048 : _GEN_780; // @[executor.scala 470:55]
  wire [7:0] _GEN_1549 = opcode_1 != 4'h0 ? _GEN_1049 : _GEN_781; // @[executor.scala 470:55]
  wire [7:0] _GEN_1550 = opcode_1 != 4'h0 ? _GEN_1054 : _GEN_782; // @[executor.scala 470:55]
  wire [7:0] _GEN_1551 = opcode_1 != 4'h0 ? _GEN_1055 : _GEN_783; // @[executor.scala 470:55]
  wire [7:0] _GEN_1552 = opcode_1 != 4'h0 ? _GEN_1056 : _GEN_784; // @[executor.scala 470:55]
  wire [7:0] _GEN_1553 = opcode_1 != 4'h0 ? _GEN_1057 : _GEN_785; // @[executor.scala 470:55]
  wire [7:0] _GEN_1554 = opcode_1 != 4'h0 ? _GEN_1062 : _GEN_786; // @[executor.scala 470:55]
  wire [7:0] _GEN_1555 = opcode_1 != 4'h0 ? _GEN_1063 : _GEN_787; // @[executor.scala 470:55]
  wire [7:0] _GEN_1556 = opcode_1 != 4'h0 ? _GEN_1064 : _GEN_788; // @[executor.scala 470:55]
  wire [7:0] _GEN_1557 = opcode_1 != 4'h0 ? _GEN_1065 : _GEN_789; // @[executor.scala 470:55]
  wire [7:0] _GEN_1558 = opcode_1 != 4'h0 ? _GEN_1070 : _GEN_790; // @[executor.scala 470:55]
  wire [7:0] _GEN_1559 = opcode_1 != 4'h0 ? _GEN_1071 : _GEN_791; // @[executor.scala 470:55]
  wire [7:0] _GEN_1560 = opcode_1 != 4'h0 ? _GEN_1072 : _GEN_792; // @[executor.scala 470:55]
  wire [7:0] _GEN_1561 = opcode_1 != 4'h0 ? _GEN_1073 : _GEN_793; // @[executor.scala 470:55]
  wire [7:0] _GEN_1562 = opcode_1 != 4'h0 ? _GEN_1078 : _GEN_794; // @[executor.scala 470:55]
  wire [7:0] _GEN_1563 = opcode_1 != 4'h0 ? _GEN_1079 : _GEN_795; // @[executor.scala 470:55]
  wire [7:0] _GEN_1564 = opcode_1 != 4'h0 ? _GEN_1080 : _GEN_796; // @[executor.scala 470:55]
  wire [7:0] _GEN_1565 = opcode_1 != 4'h0 ? _GEN_1081 : _GEN_797; // @[executor.scala 470:55]
  wire [7:0] _GEN_1566 = opcode_1 != 4'h0 ? _GEN_1086 : _GEN_798; // @[executor.scala 470:55]
  wire [7:0] _GEN_1567 = opcode_1 != 4'h0 ? _GEN_1087 : _GEN_799; // @[executor.scala 470:55]
  wire [7:0] _GEN_1568 = opcode_1 != 4'h0 ? _GEN_1088 : _GEN_800; // @[executor.scala 470:55]
  wire [7:0] _GEN_1569 = opcode_1 != 4'h0 ? _GEN_1089 : _GEN_801; // @[executor.scala 470:55]
  wire [7:0] _GEN_1570 = opcode_1 != 4'h0 ? _GEN_1094 : _GEN_802; // @[executor.scala 470:55]
  wire [7:0] _GEN_1571 = opcode_1 != 4'h0 ? _GEN_1095 : _GEN_803; // @[executor.scala 470:55]
  wire [7:0] _GEN_1572 = opcode_1 != 4'h0 ? _GEN_1096 : _GEN_804; // @[executor.scala 470:55]
  wire [7:0] _GEN_1573 = opcode_1 != 4'h0 ? _GEN_1097 : _GEN_805; // @[executor.scala 470:55]
  wire [7:0] _GEN_1574 = opcode_1 != 4'h0 ? _GEN_1102 : _GEN_806; // @[executor.scala 470:55]
  wire [7:0] _GEN_1575 = opcode_1 != 4'h0 ? _GEN_1103 : _GEN_807; // @[executor.scala 470:55]
  wire [7:0] _GEN_1576 = opcode_1 != 4'h0 ? _GEN_1104 : _GEN_808; // @[executor.scala 470:55]
  wire [7:0] _GEN_1577 = opcode_1 != 4'h0 ? _GEN_1105 : _GEN_809; // @[executor.scala 470:55]
  wire [7:0] _GEN_1578 = opcode_1 != 4'h0 ? _GEN_1110 : _GEN_810; // @[executor.scala 470:55]
  wire [7:0] _GEN_1579 = opcode_1 != 4'h0 ? _GEN_1111 : _GEN_811; // @[executor.scala 470:55]
  wire [7:0] _GEN_1580 = opcode_1 != 4'h0 ? _GEN_1112 : _GEN_812; // @[executor.scala 470:55]
  wire [7:0] _GEN_1581 = opcode_1 != 4'h0 ? _GEN_1113 : _GEN_813; // @[executor.scala 470:55]
  wire [7:0] _GEN_1582 = opcode_1 != 4'h0 ? _GEN_1118 : _GEN_814; // @[executor.scala 470:55]
  wire [7:0] _GEN_1583 = opcode_1 != 4'h0 ? _GEN_1119 : _GEN_815; // @[executor.scala 470:55]
  wire [7:0] _GEN_1584 = opcode_1 != 4'h0 ? _GEN_1120 : _GEN_816; // @[executor.scala 470:55]
  wire [7:0] _GEN_1585 = opcode_1 != 4'h0 ? _GEN_1121 : _GEN_817; // @[executor.scala 470:55]
  wire [7:0] _GEN_1586 = opcode_1 != 4'h0 ? _GEN_1126 : _GEN_818; // @[executor.scala 470:55]
  wire [7:0] _GEN_1587 = opcode_1 != 4'h0 ? _GEN_1127 : _GEN_819; // @[executor.scala 470:55]
  wire [7:0] _GEN_1588 = opcode_1 != 4'h0 ? _GEN_1128 : _GEN_820; // @[executor.scala 470:55]
  wire [7:0] _GEN_1589 = opcode_1 != 4'h0 ? _GEN_1129 : _GEN_821; // @[executor.scala 470:55]
  wire [7:0] _GEN_1590 = opcode_1 != 4'h0 ? _GEN_1134 : _GEN_822; // @[executor.scala 470:55]
  wire [7:0] _GEN_1591 = opcode_1 != 4'h0 ? _GEN_1135 : _GEN_823; // @[executor.scala 470:55]
  wire [7:0] _GEN_1592 = opcode_1 != 4'h0 ? _GEN_1136 : _GEN_824; // @[executor.scala 470:55]
  wire [7:0] _GEN_1593 = opcode_1 != 4'h0 ? _GEN_1137 : _GEN_825; // @[executor.scala 470:55]
  wire [7:0] _GEN_1594 = opcode_1 != 4'h0 ? _GEN_1142 : _GEN_826; // @[executor.scala 470:55]
  wire [7:0] _GEN_1595 = opcode_1 != 4'h0 ? _GEN_1143 : _GEN_827; // @[executor.scala 470:55]
  wire [7:0] _GEN_1596 = opcode_1 != 4'h0 ? _GEN_1144 : _GEN_828; // @[executor.scala 470:55]
  wire [7:0] _GEN_1597 = opcode_1 != 4'h0 ? _GEN_1145 : _GEN_829; // @[executor.scala 470:55]
  wire [7:0] _GEN_1598 = opcode_1 != 4'h0 ? _GEN_1150 : _GEN_830; // @[executor.scala 470:55]
  wire [7:0] _GEN_1599 = opcode_1 != 4'h0 ? _GEN_1151 : _GEN_831; // @[executor.scala 470:55]
  wire [7:0] _GEN_1600 = opcode_1 != 4'h0 ? _GEN_1152 : _GEN_832; // @[executor.scala 470:55]
  wire [7:0] _GEN_1601 = opcode_1 != 4'h0 ? _GEN_1153 : _GEN_833; // @[executor.scala 470:55]
  wire [7:0] _GEN_1602 = opcode_1 != 4'h0 ? _GEN_1158 : _GEN_834; // @[executor.scala 470:55]
  wire [7:0] _GEN_1603 = opcode_1 != 4'h0 ? _GEN_1159 : _GEN_835; // @[executor.scala 470:55]
  wire [7:0] _GEN_1604 = opcode_1 != 4'h0 ? _GEN_1160 : _GEN_836; // @[executor.scala 470:55]
  wire [7:0] _GEN_1605 = opcode_1 != 4'h0 ? _GEN_1161 : _GEN_837; // @[executor.scala 470:55]
  wire [7:0] _GEN_1606 = opcode_1 != 4'h0 ? _GEN_1166 : _GEN_838; // @[executor.scala 470:55]
  wire [7:0] _GEN_1607 = opcode_1 != 4'h0 ? _GEN_1167 : _GEN_839; // @[executor.scala 470:55]
  wire [7:0] _GEN_1608 = opcode_1 != 4'h0 ? _GEN_1168 : _GEN_840; // @[executor.scala 470:55]
  wire [7:0] _GEN_1609 = opcode_1 != 4'h0 ? _GEN_1169 : _GEN_841; // @[executor.scala 470:55]
  wire [7:0] _GEN_1610 = opcode_1 != 4'h0 ? _GEN_1174 : _GEN_842; // @[executor.scala 470:55]
  wire [7:0] _GEN_1611 = opcode_1 != 4'h0 ? _GEN_1175 : _GEN_843; // @[executor.scala 470:55]
  wire [7:0] _GEN_1612 = opcode_1 != 4'h0 ? _GEN_1176 : _GEN_844; // @[executor.scala 470:55]
  wire [7:0] _GEN_1613 = opcode_1 != 4'h0 ? _GEN_1177 : _GEN_845; // @[executor.scala 470:55]
  wire [7:0] _GEN_1614 = opcode_1 != 4'h0 ? _GEN_1182 : _GEN_846; // @[executor.scala 470:55]
  wire [7:0] _GEN_1615 = opcode_1 != 4'h0 ? _GEN_1183 : _GEN_847; // @[executor.scala 470:55]
  wire [7:0] _GEN_1616 = opcode_1 != 4'h0 ? _GEN_1184 : _GEN_848; // @[executor.scala 470:55]
  wire [7:0] _GEN_1617 = opcode_1 != 4'h0 ? _GEN_1185 : _GEN_849; // @[executor.scala 470:55]
  wire [7:0] _GEN_1618 = opcode_1 != 4'h0 ? _GEN_1190 : _GEN_850; // @[executor.scala 470:55]
  wire [7:0] _GEN_1619 = opcode_1 != 4'h0 ? _GEN_1191 : _GEN_851; // @[executor.scala 470:55]
  wire [7:0] _GEN_1620 = opcode_1 != 4'h0 ? _GEN_1192 : _GEN_852; // @[executor.scala 470:55]
  wire [7:0] _GEN_1621 = opcode_1 != 4'h0 ? _GEN_1193 : _GEN_853; // @[executor.scala 470:55]
  wire [7:0] _GEN_1622 = opcode_1 != 4'h0 ? _GEN_1198 : _GEN_854; // @[executor.scala 470:55]
  wire [7:0] _GEN_1623 = opcode_1 != 4'h0 ? _GEN_1199 : _GEN_855; // @[executor.scala 470:55]
  wire [7:0] _GEN_1624 = opcode_1 != 4'h0 ? _GEN_1200 : _GEN_856; // @[executor.scala 470:55]
  wire [7:0] _GEN_1625 = opcode_1 != 4'h0 ? _GEN_1201 : _GEN_857; // @[executor.scala 470:55]
  wire [7:0] _GEN_1626 = opcode_1 != 4'h0 ? _GEN_1206 : _GEN_858; // @[executor.scala 470:55]
  wire [7:0] _GEN_1627 = opcode_1 != 4'h0 ? _GEN_1207 : _GEN_859; // @[executor.scala 470:55]
  wire [7:0] _GEN_1628 = opcode_1 != 4'h0 ? _GEN_1208 : _GEN_860; // @[executor.scala 470:55]
  wire [7:0] _GEN_1629 = opcode_1 != 4'h0 ? _GEN_1209 : _GEN_861; // @[executor.scala 470:55]
  wire [7:0] _GEN_1630 = opcode_1 != 4'h0 ? _GEN_1214 : _GEN_862; // @[executor.scala 470:55]
  wire [7:0] _GEN_1631 = opcode_1 != 4'h0 ? _GEN_1215 : _GEN_863; // @[executor.scala 470:55]
  wire [7:0] _GEN_1632 = opcode_1 != 4'h0 ? _GEN_1216 : _GEN_864; // @[executor.scala 470:55]
  wire [7:0] _GEN_1633 = opcode_1 != 4'h0 ? _GEN_1217 : _GEN_865; // @[executor.scala 470:55]
  wire [7:0] _GEN_1634 = opcode_1 != 4'h0 ? _GEN_1222 : _GEN_866; // @[executor.scala 470:55]
  wire [7:0] _GEN_1635 = opcode_1 != 4'h0 ? _GEN_1223 : _GEN_867; // @[executor.scala 470:55]
  wire [7:0] _GEN_1636 = opcode_1 != 4'h0 ? _GEN_1224 : _GEN_868; // @[executor.scala 470:55]
  wire [7:0] _GEN_1637 = opcode_1 != 4'h0 ? _GEN_1225 : _GEN_869; // @[executor.scala 470:55]
  wire [7:0] _GEN_1638 = opcode_1 != 4'h0 ? _GEN_1230 : _GEN_870; // @[executor.scala 470:55]
  wire [7:0] _GEN_1639 = opcode_1 != 4'h0 ? _GEN_1231 : _GEN_871; // @[executor.scala 470:55]
  wire [7:0] _GEN_1640 = opcode_1 != 4'h0 ? _GEN_1232 : _GEN_872; // @[executor.scala 470:55]
  wire [7:0] _GEN_1641 = opcode_1 != 4'h0 ? _GEN_1233 : _GEN_873; // @[executor.scala 470:55]
  wire [7:0] _GEN_1642 = opcode_1 != 4'h0 ? _GEN_1238 : _GEN_874; // @[executor.scala 470:55]
  wire [7:0] _GEN_1643 = opcode_1 != 4'h0 ? _GEN_1239 : _GEN_875; // @[executor.scala 470:55]
  wire [7:0] _GEN_1644 = opcode_1 != 4'h0 ? _GEN_1240 : _GEN_876; // @[executor.scala 470:55]
  wire [7:0] _GEN_1645 = opcode_1 != 4'h0 ? _GEN_1241 : _GEN_877; // @[executor.scala 470:55]
  wire [7:0] _GEN_1646 = opcode_1 != 4'h0 ? _GEN_1246 : _GEN_878; // @[executor.scala 470:55]
  wire [7:0] _GEN_1647 = opcode_1 != 4'h0 ? _GEN_1247 : _GEN_879; // @[executor.scala 470:55]
  wire [7:0] _GEN_1648 = opcode_1 != 4'h0 ? _GEN_1248 : _GEN_880; // @[executor.scala 470:55]
  wire [7:0] _GEN_1649 = opcode_1 != 4'h0 ? _GEN_1249 : _GEN_881; // @[executor.scala 470:55]
  wire [7:0] _GEN_1650 = opcode_1 != 4'h0 ? _GEN_1254 : _GEN_882; // @[executor.scala 470:55]
  wire [7:0] _GEN_1651 = opcode_1 != 4'h0 ? _GEN_1255 : _GEN_883; // @[executor.scala 470:55]
  wire [7:0] _GEN_1652 = opcode_1 != 4'h0 ? _GEN_1256 : _GEN_884; // @[executor.scala 470:55]
  wire [7:0] _GEN_1653 = opcode_1 != 4'h0 ? _GEN_1257 : _GEN_885; // @[executor.scala 470:55]
  wire [7:0] _GEN_1654 = opcode_1 != 4'h0 ? _GEN_1262 : _GEN_886; // @[executor.scala 470:55]
  wire [7:0] _GEN_1655 = opcode_1 != 4'h0 ? _GEN_1263 : _GEN_887; // @[executor.scala 470:55]
  wire [7:0] _GEN_1656 = opcode_1 != 4'h0 ? _GEN_1264 : _GEN_888; // @[executor.scala 470:55]
  wire [7:0] _GEN_1657 = opcode_1 != 4'h0 ? _GEN_1265 : _GEN_889; // @[executor.scala 470:55]
  wire [7:0] _GEN_1658 = opcode_1 != 4'h0 ? _GEN_1270 : _GEN_890; // @[executor.scala 470:55]
  wire [7:0] _GEN_1659 = opcode_1 != 4'h0 ? _GEN_1271 : _GEN_891; // @[executor.scala 470:55]
  wire [7:0] _GEN_1660 = opcode_1 != 4'h0 ? _GEN_1272 : _GEN_892; // @[executor.scala 470:55]
  wire [7:0] _GEN_1661 = opcode_1 != 4'h0 ? _GEN_1273 : _GEN_893; // @[executor.scala 470:55]
  wire [7:0] _GEN_1662 = opcode_1 != 4'h0 ? _GEN_1278 : _GEN_894; // @[executor.scala 470:55]
  wire [7:0] _GEN_1663 = opcode_1 != 4'h0 ? _GEN_1279 : _GEN_895; // @[executor.scala 470:55]
  wire [7:0] _GEN_1664 = opcode_1 != 4'h0 ? _GEN_1280 : _GEN_896; // @[executor.scala 470:55]
  wire [7:0] _GEN_1665 = opcode_1 != 4'h0 ? _GEN_1281 : _GEN_897; // @[executor.scala 470:55]
  wire [7:0] _GEN_1666 = opcode_1 != 4'h0 ? _GEN_1286 : _GEN_898; // @[executor.scala 470:55]
  wire [7:0] _GEN_1667 = opcode_1 != 4'h0 ? _GEN_1287 : _GEN_899; // @[executor.scala 470:55]
  wire [7:0] _GEN_1668 = opcode_1 != 4'h0 ? _GEN_1288 : _GEN_900; // @[executor.scala 470:55]
  wire [7:0] _GEN_1669 = opcode_1 != 4'h0 ? _GEN_1289 : _GEN_901; // @[executor.scala 470:55]
  wire [7:0] _GEN_1670 = opcode_1 != 4'h0 ? _GEN_1294 : _GEN_902; // @[executor.scala 470:55]
  wire [7:0] _GEN_1671 = opcode_1 != 4'h0 ? _GEN_1295 : _GEN_903; // @[executor.scala 470:55]
  wire [7:0] _GEN_1672 = opcode_1 != 4'h0 ? _GEN_1296 : _GEN_904; // @[executor.scala 470:55]
  wire [7:0] _GEN_1673 = opcode_1 != 4'h0 ? _GEN_1297 : _GEN_905; // @[executor.scala 470:55]
  wire [7:0] _GEN_1674 = opcode_1 != 4'h0 ? _GEN_1302 : _GEN_906; // @[executor.scala 470:55]
  wire [7:0] _GEN_1675 = opcode_1 != 4'h0 ? _GEN_1303 : _GEN_907; // @[executor.scala 470:55]
  wire [7:0] _GEN_1676 = opcode_1 != 4'h0 ? _GEN_1304 : _GEN_908; // @[executor.scala 470:55]
  wire [7:0] _GEN_1677 = opcode_1 != 4'h0 ? _GEN_1305 : _GEN_909; // @[executor.scala 470:55]
  wire [7:0] _GEN_1678 = opcode_1 != 4'h0 ? _GEN_1310 : _GEN_910; // @[executor.scala 470:55]
  wire [7:0] _GEN_1679 = opcode_1 != 4'h0 ? _GEN_1311 : _GEN_911; // @[executor.scala 470:55]
  wire [7:0] _GEN_1680 = opcode_1 != 4'h0 ? _GEN_1312 : _GEN_912; // @[executor.scala 470:55]
  wire [7:0] _GEN_1681 = opcode_1 != 4'h0 ? _GEN_1313 : _GEN_913; // @[executor.scala 470:55]
  wire [7:0] _GEN_1682 = opcode_1 != 4'h0 ? _GEN_1318 : _GEN_914; // @[executor.scala 470:55]
  wire [7:0] _GEN_1683 = opcode_1 != 4'h0 ? _GEN_1319 : _GEN_915; // @[executor.scala 470:55]
  wire [7:0] _GEN_1684 = opcode_1 != 4'h0 ? _GEN_1320 : _GEN_916; // @[executor.scala 470:55]
  wire [7:0] _GEN_1685 = opcode_1 != 4'h0 ? _GEN_1321 : _GEN_917; // @[executor.scala 470:55]
  wire [7:0] _GEN_1686 = opcode_1 != 4'h0 ? _GEN_1326 : _GEN_918; // @[executor.scala 470:55]
  wire [7:0] _GEN_1687 = opcode_1 != 4'h0 ? _GEN_1327 : _GEN_919; // @[executor.scala 470:55]
  wire [7:0] _GEN_1688 = opcode_1 != 4'h0 ? _GEN_1328 : _GEN_920; // @[executor.scala 470:55]
  wire [7:0] _GEN_1689 = opcode_1 != 4'h0 ? _GEN_1329 : _GEN_921; // @[executor.scala 470:55]
  wire [7:0] _GEN_1690 = opcode_1 != 4'h0 ? _GEN_1334 : _GEN_922; // @[executor.scala 470:55]
  wire [7:0] _GEN_1691 = opcode_1 != 4'h0 ? _GEN_1335 : _GEN_923; // @[executor.scala 470:55]
  wire [7:0] _GEN_1692 = opcode_1 != 4'h0 ? _GEN_1336 : _GEN_924; // @[executor.scala 470:55]
  wire [7:0] _GEN_1693 = opcode_1 != 4'h0 ? _GEN_1337 : _GEN_925; // @[executor.scala 470:55]
  wire [7:0] _GEN_1694 = opcode_1 != 4'h0 ? _GEN_1342 : _GEN_926; // @[executor.scala 470:55]
  wire [7:0] _GEN_1695 = opcode_1 != 4'h0 ? _GEN_1343 : _GEN_927; // @[executor.scala 470:55]
  wire [7:0] _GEN_1696 = opcode_1 != 4'h0 ? _GEN_1344 : _GEN_928; // @[executor.scala 470:55]
  wire [7:0] _GEN_1697 = opcode_1 != 4'h0 ? _GEN_1345 : _GEN_929; // @[executor.scala 470:55]
  wire [7:0] _GEN_1698 = opcode_1 != 4'h0 ? _GEN_1350 : _GEN_930; // @[executor.scala 470:55]
  wire [7:0] _GEN_1699 = opcode_1 != 4'h0 ? _GEN_1351 : _GEN_931; // @[executor.scala 470:55]
  wire [7:0] _GEN_1700 = opcode_1 != 4'h0 ? _GEN_1352 : _GEN_932; // @[executor.scala 470:55]
  wire [7:0] _GEN_1701 = opcode_1 != 4'h0 ? _GEN_1353 : _GEN_933; // @[executor.scala 470:55]
  wire [7:0] _GEN_1702 = opcode_1 != 4'h0 ? _GEN_1358 : _GEN_934; // @[executor.scala 470:55]
  wire [7:0] _GEN_1703 = opcode_1 != 4'h0 ? _GEN_1359 : _GEN_935; // @[executor.scala 470:55]
  wire [7:0] _GEN_1704 = opcode_1 != 4'h0 ? _GEN_1360 : _GEN_936; // @[executor.scala 470:55]
  wire [7:0] _GEN_1705 = opcode_1 != 4'h0 ? _GEN_1361 : _GEN_937; // @[executor.scala 470:55]
  wire [7:0] _GEN_1706 = opcode_1 != 4'h0 ? _GEN_1366 : _GEN_938; // @[executor.scala 470:55]
  wire [7:0] _GEN_1707 = opcode_1 != 4'h0 ? _GEN_1367 : _GEN_939; // @[executor.scala 470:55]
  wire [7:0] _GEN_1708 = opcode_1 != 4'h0 ? _GEN_1368 : _GEN_940; // @[executor.scala 470:55]
  wire [7:0] _GEN_1709 = opcode_1 != 4'h0 ? _GEN_1369 : _GEN_941; // @[executor.scala 470:55]
  wire [7:0] _GEN_1710 = opcode_1 != 4'h0 ? _GEN_1374 : _GEN_942; // @[executor.scala 470:55]
  wire [7:0] _GEN_1711 = opcode_1 != 4'h0 ? _GEN_1375 : _GEN_943; // @[executor.scala 470:55]
  wire [7:0] _GEN_1712 = opcode_1 != 4'h0 ? _GEN_1376 : _GEN_944; // @[executor.scala 470:55]
  wire [7:0] _GEN_1713 = opcode_1 != 4'h0 ? _GEN_1377 : _GEN_945; // @[executor.scala 470:55]
  wire [7:0] _GEN_1714 = opcode_1 != 4'h0 ? _GEN_1382 : _GEN_946; // @[executor.scala 470:55]
  wire [7:0] _GEN_1715 = opcode_1 != 4'h0 ? _GEN_1383 : _GEN_947; // @[executor.scala 470:55]
  wire [7:0] _GEN_1716 = opcode_1 != 4'h0 ? _GEN_1384 : _GEN_948; // @[executor.scala 470:55]
  wire [7:0] _GEN_1717 = opcode_1 != 4'h0 ? _GEN_1385 : _GEN_949; // @[executor.scala 470:55]
  wire [7:0] _GEN_1718 = opcode_1 != 4'h0 ? _GEN_1390 : _GEN_950; // @[executor.scala 470:55]
  wire [7:0] _GEN_1719 = opcode_1 != 4'h0 ? _GEN_1391 : _GEN_951; // @[executor.scala 470:55]
  wire [7:0] _GEN_1720 = opcode_1 != 4'h0 ? _GEN_1392 : _GEN_952; // @[executor.scala 470:55]
  wire [7:0] _GEN_1721 = opcode_1 != 4'h0 ? _GEN_1393 : _GEN_953; // @[executor.scala 470:55]
  wire [7:0] _GEN_1722 = opcode_1 != 4'h0 ? _GEN_1398 : _GEN_954; // @[executor.scala 470:55]
  wire [7:0] _GEN_1723 = opcode_1 != 4'h0 ? _GEN_1399 : _GEN_955; // @[executor.scala 470:55]
  wire [7:0] _GEN_1724 = opcode_1 != 4'h0 ? _GEN_1400 : _GEN_956; // @[executor.scala 470:55]
  wire [7:0] _GEN_1725 = opcode_1 != 4'h0 ? _GEN_1401 : _GEN_957; // @[executor.scala 470:55]
  wire [7:0] _GEN_1726 = opcode_1 != 4'h0 ? _GEN_1406 : _GEN_958; // @[executor.scala 470:55]
  wire [7:0] _GEN_1727 = opcode_1 != 4'h0 ? _GEN_1407 : _GEN_959; // @[executor.scala 470:55]
  wire [7:0] _GEN_1728 = opcode_1 != 4'h0 ? _GEN_1408 : _GEN_960; // @[executor.scala 470:55]
  wire [7:0] _GEN_1729 = opcode_1 != 4'h0 ? _GEN_1409 : _GEN_961; // @[executor.scala 470:55]
  wire [7:0] _GEN_1730 = opcode_1 != 4'h0 ? _GEN_1414 : _GEN_962; // @[executor.scala 470:55]
  wire [7:0] _GEN_1731 = opcode_1 != 4'h0 ? _GEN_1415 : _GEN_963; // @[executor.scala 470:55]
  wire [7:0] _GEN_1732 = opcode_1 != 4'h0 ? _GEN_1416 : _GEN_964; // @[executor.scala 470:55]
  wire [7:0] _GEN_1733 = opcode_1 != 4'h0 ? _GEN_1417 : _GEN_965; // @[executor.scala 470:55]
  wire [7:0] _GEN_1734 = opcode_1 != 4'h0 ? _GEN_1422 : _GEN_966; // @[executor.scala 470:55]
  wire [7:0] _GEN_1735 = opcode_1 != 4'h0 ? _GEN_1423 : _GEN_967; // @[executor.scala 470:55]
  wire [7:0] _GEN_1736 = opcode_1 != 4'h0 ? _GEN_1424 : _GEN_968; // @[executor.scala 470:55]
  wire [7:0] _GEN_1737 = opcode_1 != 4'h0 ? _GEN_1425 : _GEN_969; // @[executor.scala 470:55]
  wire [7:0] _GEN_1738 = opcode_1 != 4'h0 ? _GEN_1430 : _GEN_970; // @[executor.scala 470:55]
  wire [7:0] _GEN_1739 = opcode_1 != 4'h0 ? _GEN_1431 : _GEN_971; // @[executor.scala 470:55]
  wire [7:0] _GEN_1740 = opcode_1 != 4'h0 ? _GEN_1432 : _GEN_972; // @[executor.scala 470:55]
  wire [7:0] _GEN_1741 = opcode_1 != 4'h0 ? _GEN_1433 : _GEN_973; // @[executor.scala 470:55]
  wire [7:0] _GEN_1742 = opcode_1 != 4'h0 ? _GEN_1438 : _GEN_974; // @[executor.scala 470:55]
  wire [7:0] _GEN_1743 = opcode_1 != 4'h0 ? _GEN_1439 : _GEN_975; // @[executor.scala 470:55]
  wire [7:0] _GEN_1744 = opcode_1 != 4'h0 ? _GEN_1440 : _GEN_976; // @[executor.scala 470:55]
  wire [7:0] _GEN_1745 = opcode_1 != 4'h0 ? _GEN_1441 : _GEN_977; // @[executor.scala 470:55]
  wire [7:0] _GEN_1746 = opcode_1 != 4'h0 ? _GEN_1446 : _GEN_978; // @[executor.scala 470:55]
  wire [7:0] _GEN_1747 = opcode_1 != 4'h0 ? _GEN_1447 : _GEN_979; // @[executor.scala 470:55]
  wire [7:0] _GEN_1748 = opcode_1 != 4'h0 ? _GEN_1448 : _GEN_980; // @[executor.scala 470:55]
  wire [7:0] _GEN_1749 = opcode_1 != 4'h0 ? _GEN_1449 : _GEN_981; // @[executor.scala 470:55]
  wire [7:0] _GEN_1750 = opcode_1 != 4'h0 ? _GEN_1454 : _GEN_982; // @[executor.scala 470:55]
  wire [7:0] _GEN_1751 = opcode_1 != 4'h0 ? _GEN_1455 : _GEN_983; // @[executor.scala 470:55]
  wire [7:0] _GEN_1752 = opcode_1 != 4'h0 ? _GEN_1456 : _GEN_984; // @[executor.scala 470:55]
  wire [7:0] _GEN_1753 = opcode_1 != 4'h0 ? _GEN_1457 : _GEN_985; // @[executor.scala 470:55]
  wire [7:0] _GEN_1754 = opcode_1 != 4'h0 ? _GEN_1462 : _GEN_986; // @[executor.scala 470:55]
  wire [7:0] _GEN_1755 = opcode_1 != 4'h0 ? _GEN_1463 : _GEN_987; // @[executor.scala 470:55]
  wire [7:0] _GEN_1756 = opcode_1 != 4'h0 ? _GEN_1464 : _GEN_988; // @[executor.scala 470:55]
  wire [7:0] _GEN_1757 = opcode_1 != 4'h0 ? _GEN_1465 : _GEN_989; // @[executor.scala 470:55]
  wire [7:0] _GEN_1758 = opcode_1 != 4'h0 ? _GEN_1470 : _GEN_990; // @[executor.scala 470:55]
  wire [7:0] _GEN_1759 = opcode_1 != 4'h0 ? _GEN_1471 : _GEN_991; // @[executor.scala 470:55]
  wire [7:0] _GEN_1760 = opcode_1 != 4'h0 ? _GEN_1472 : _GEN_992; // @[executor.scala 470:55]
  wire [7:0] _GEN_1761 = opcode_1 != 4'h0 ? _GEN_1473 : _GEN_993; // @[executor.scala 470:55]
  wire [7:0] _GEN_1762 = opcode_1 != 4'h0 ? _GEN_1478 : _GEN_994; // @[executor.scala 470:55]
  wire [7:0] _GEN_1763 = opcode_1 != 4'h0 ? _GEN_1479 : _GEN_995; // @[executor.scala 470:55]
  wire [7:0] _GEN_1764 = opcode_1 != 4'h0 ? _GEN_1480 : _GEN_996; // @[executor.scala 470:55]
  wire [7:0] _GEN_1765 = opcode_1 != 4'h0 ? _GEN_1481 : _GEN_997; // @[executor.scala 470:55]
  wire [7:0] _GEN_1766 = opcode_1 != 4'h0 ? _GEN_1486 : _GEN_998; // @[executor.scala 470:55]
  wire [7:0] _GEN_1767 = opcode_1 != 4'h0 ? _GEN_1487 : _GEN_999; // @[executor.scala 470:55]
  wire [7:0] _GEN_1768 = opcode_1 != 4'h0 ? _GEN_1488 : _GEN_1000; // @[executor.scala 470:55]
  wire [7:0] _GEN_1769 = opcode_1 != 4'h0 ? _GEN_1489 : _GEN_1001; // @[executor.scala 470:55]
  wire [7:0] _GEN_1770 = opcode_1 != 4'h0 ? _GEN_1494 : _GEN_1002; // @[executor.scala 470:55]
  wire [7:0] _GEN_1771 = opcode_1 != 4'h0 ? _GEN_1495 : _GEN_1003; // @[executor.scala 470:55]
  wire [7:0] _GEN_1772 = opcode_1 != 4'h0 ? _GEN_1496 : _GEN_1004; // @[executor.scala 470:55]
  wire [7:0] _GEN_1773 = opcode_1 != 4'h0 ? _GEN_1497 : _GEN_1005; // @[executor.scala 470:55]
  wire [7:0] _GEN_1774 = opcode_1 != 4'h0 ? _GEN_1502 : _GEN_1006; // @[executor.scala 470:55]
  wire [7:0] _GEN_1775 = opcode_1 != 4'h0 ? _GEN_1503 : _GEN_1007; // @[executor.scala 470:55]
  wire [7:0] _GEN_1776 = opcode_1 != 4'h0 ? _GEN_1504 : _GEN_1008; // @[executor.scala 470:55]
  wire [7:0] _GEN_1777 = opcode_1 != 4'h0 ? _GEN_1505 : _GEN_1009; // @[executor.scala 470:55]
  wire [7:0] _GEN_1778 = opcode_1 != 4'h0 ? _GEN_1510 : _GEN_1010; // @[executor.scala 470:55]
  wire [7:0] _GEN_1779 = opcode_1 != 4'h0 ? _GEN_1511 : _GEN_1011; // @[executor.scala 470:55]
  wire [7:0] _GEN_1780 = opcode_1 != 4'h0 ? _GEN_1512 : _GEN_1012; // @[executor.scala 470:55]
  wire [7:0] _GEN_1781 = opcode_1 != 4'h0 ? _GEN_1513 : _GEN_1013; // @[executor.scala 470:55]
  wire [7:0] _GEN_1782 = opcode_1 != 4'h0 ? _GEN_1518 : _GEN_1014; // @[executor.scala 470:55]
  wire [7:0] _GEN_1783 = opcode_1 != 4'h0 ? _GEN_1519 : _GEN_1015; // @[executor.scala 470:55]
  wire [7:0] _GEN_1784 = opcode_1 != 4'h0 ? _GEN_1520 : _GEN_1016; // @[executor.scala 470:55]
  wire [7:0] _GEN_1785 = opcode_1 != 4'h0 ? _GEN_1521 : _GEN_1017; // @[executor.scala 470:55]
  wire [7:0] _GEN_1786 = opcode_1 != 4'h0 ? _GEN_1526 : _GEN_1018; // @[executor.scala 470:55]
  wire [7:0] _GEN_1787 = opcode_1 != 4'h0 ? _GEN_1527 : _GEN_1019; // @[executor.scala 470:55]
  wire [7:0] _GEN_1788 = opcode_1 != 4'h0 ? _GEN_1528 : _GEN_1020; // @[executor.scala 470:55]
  wire [7:0] _GEN_1789 = opcode_1 != 4'h0 ? _GEN_1529 : _GEN_1021; // @[executor.scala 470:55]
  wire [7:0] _GEN_1790 = opcode_1 != 4'h0 ? _GEN_1534 : _GEN_1022; // @[executor.scala 470:55]
  wire [7:0] _GEN_1791 = opcode_1 != 4'h0 ? _GEN_1535 : _GEN_1023; // @[executor.scala 470:55]
  wire [7:0] _GEN_1792 = opcode_1 != 4'h0 ? _GEN_1536 : _GEN_1024; // @[executor.scala 470:55]
  wire [7:0] _GEN_1793 = opcode_1 != 4'h0 ? _GEN_1537 : _GEN_1025; // @[executor.scala 470:55]
  wire [7:0] _GEN_1796 = opcode_1 == 4'hf ? _GEN_770 : _GEN_1538; // @[executor.scala 466:52]
  wire [7:0] _GEN_1797 = opcode_1 == 4'hf ? _GEN_771 : _GEN_1539; // @[executor.scala 466:52]
  wire [7:0] _GEN_1798 = opcode_1 == 4'hf ? _GEN_772 : _GEN_1540; // @[executor.scala 466:52]
  wire [7:0] _GEN_1799 = opcode_1 == 4'hf ? _GEN_773 : _GEN_1541; // @[executor.scala 466:52]
  wire [7:0] _GEN_1800 = opcode_1 == 4'hf ? _GEN_774 : _GEN_1542; // @[executor.scala 466:52]
  wire [7:0] _GEN_1801 = opcode_1 == 4'hf ? _GEN_775 : _GEN_1543; // @[executor.scala 466:52]
  wire [7:0] _GEN_1802 = opcode_1 == 4'hf ? _GEN_776 : _GEN_1544; // @[executor.scala 466:52]
  wire [7:0] _GEN_1803 = opcode_1 == 4'hf ? _GEN_777 : _GEN_1545; // @[executor.scala 466:52]
  wire [7:0] _GEN_1804 = opcode_1 == 4'hf ? _GEN_778 : _GEN_1546; // @[executor.scala 466:52]
  wire [7:0] _GEN_1805 = opcode_1 == 4'hf ? _GEN_779 : _GEN_1547; // @[executor.scala 466:52]
  wire [7:0] _GEN_1806 = opcode_1 == 4'hf ? _GEN_780 : _GEN_1548; // @[executor.scala 466:52]
  wire [7:0] _GEN_1807 = opcode_1 == 4'hf ? _GEN_781 : _GEN_1549; // @[executor.scala 466:52]
  wire [7:0] _GEN_1808 = opcode_1 == 4'hf ? _GEN_782 : _GEN_1550; // @[executor.scala 466:52]
  wire [7:0] _GEN_1809 = opcode_1 == 4'hf ? _GEN_783 : _GEN_1551; // @[executor.scala 466:52]
  wire [7:0] _GEN_1810 = opcode_1 == 4'hf ? _GEN_784 : _GEN_1552; // @[executor.scala 466:52]
  wire [7:0] _GEN_1811 = opcode_1 == 4'hf ? _GEN_785 : _GEN_1553; // @[executor.scala 466:52]
  wire [7:0] _GEN_1812 = opcode_1 == 4'hf ? _GEN_786 : _GEN_1554; // @[executor.scala 466:52]
  wire [7:0] _GEN_1813 = opcode_1 == 4'hf ? _GEN_787 : _GEN_1555; // @[executor.scala 466:52]
  wire [7:0] _GEN_1814 = opcode_1 == 4'hf ? _GEN_788 : _GEN_1556; // @[executor.scala 466:52]
  wire [7:0] _GEN_1815 = opcode_1 == 4'hf ? _GEN_789 : _GEN_1557; // @[executor.scala 466:52]
  wire [7:0] _GEN_1816 = opcode_1 == 4'hf ? _GEN_790 : _GEN_1558; // @[executor.scala 466:52]
  wire [7:0] _GEN_1817 = opcode_1 == 4'hf ? _GEN_791 : _GEN_1559; // @[executor.scala 466:52]
  wire [7:0] _GEN_1818 = opcode_1 == 4'hf ? _GEN_792 : _GEN_1560; // @[executor.scala 466:52]
  wire [7:0] _GEN_1819 = opcode_1 == 4'hf ? _GEN_793 : _GEN_1561; // @[executor.scala 466:52]
  wire [7:0] _GEN_1820 = opcode_1 == 4'hf ? _GEN_794 : _GEN_1562; // @[executor.scala 466:52]
  wire [7:0] _GEN_1821 = opcode_1 == 4'hf ? _GEN_795 : _GEN_1563; // @[executor.scala 466:52]
  wire [7:0] _GEN_1822 = opcode_1 == 4'hf ? _GEN_796 : _GEN_1564; // @[executor.scala 466:52]
  wire [7:0] _GEN_1823 = opcode_1 == 4'hf ? _GEN_797 : _GEN_1565; // @[executor.scala 466:52]
  wire [7:0] _GEN_1824 = opcode_1 == 4'hf ? _GEN_798 : _GEN_1566; // @[executor.scala 466:52]
  wire [7:0] _GEN_1825 = opcode_1 == 4'hf ? _GEN_799 : _GEN_1567; // @[executor.scala 466:52]
  wire [7:0] _GEN_1826 = opcode_1 == 4'hf ? _GEN_800 : _GEN_1568; // @[executor.scala 466:52]
  wire [7:0] _GEN_1827 = opcode_1 == 4'hf ? _GEN_801 : _GEN_1569; // @[executor.scala 466:52]
  wire [7:0] _GEN_1828 = opcode_1 == 4'hf ? _GEN_802 : _GEN_1570; // @[executor.scala 466:52]
  wire [7:0] _GEN_1829 = opcode_1 == 4'hf ? _GEN_803 : _GEN_1571; // @[executor.scala 466:52]
  wire [7:0] _GEN_1830 = opcode_1 == 4'hf ? _GEN_804 : _GEN_1572; // @[executor.scala 466:52]
  wire [7:0] _GEN_1831 = opcode_1 == 4'hf ? _GEN_805 : _GEN_1573; // @[executor.scala 466:52]
  wire [7:0] _GEN_1832 = opcode_1 == 4'hf ? _GEN_806 : _GEN_1574; // @[executor.scala 466:52]
  wire [7:0] _GEN_1833 = opcode_1 == 4'hf ? _GEN_807 : _GEN_1575; // @[executor.scala 466:52]
  wire [7:0] _GEN_1834 = opcode_1 == 4'hf ? _GEN_808 : _GEN_1576; // @[executor.scala 466:52]
  wire [7:0] _GEN_1835 = opcode_1 == 4'hf ? _GEN_809 : _GEN_1577; // @[executor.scala 466:52]
  wire [7:0] _GEN_1836 = opcode_1 == 4'hf ? _GEN_810 : _GEN_1578; // @[executor.scala 466:52]
  wire [7:0] _GEN_1837 = opcode_1 == 4'hf ? _GEN_811 : _GEN_1579; // @[executor.scala 466:52]
  wire [7:0] _GEN_1838 = opcode_1 == 4'hf ? _GEN_812 : _GEN_1580; // @[executor.scala 466:52]
  wire [7:0] _GEN_1839 = opcode_1 == 4'hf ? _GEN_813 : _GEN_1581; // @[executor.scala 466:52]
  wire [7:0] _GEN_1840 = opcode_1 == 4'hf ? _GEN_814 : _GEN_1582; // @[executor.scala 466:52]
  wire [7:0] _GEN_1841 = opcode_1 == 4'hf ? _GEN_815 : _GEN_1583; // @[executor.scala 466:52]
  wire [7:0] _GEN_1842 = opcode_1 == 4'hf ? _GEN_816 : _GEN_1584; // @[executor.scala 466:52]
  wire [7:0] _GEN_1843 = opcode_1 == 4'hf ? _GEN_817 : _GEN_1585; // @[executor.scala 466:52]
  wire [7:0] _GEN_1844 = opcode_1 == 4'hf ? _GEN_818 : _GEN_1586; // @[executor.scala 466:52]
  wire [7:0] _GEN_1845 = opcode_1 == 4'hf ? _GEN_819 : _GEN_1587; // @[executor.scala 466:52]
  wire [7:0] _GEN_1846 = opcode_1 == 4'hf ? _GEN_820 : _GEN_1588; // @[executor.scala 466:52]
  wire [7:0] _GEN_1847 = opcode_1 == 4'hf ? _GEN_821 : _GEN_1589; // @[executor.scala 466:52]
  wire [7:0] _GEN_1848 = opcode_1 == 4'hf ? _GEN_822 : _GEN_1590; // @[executor.scala 466:52]
  wire [7:0] _GEN_1849 = opcode_1 == 4'hf ? _GEN_823 : _GEN_1591; // @[executor.scala 466:52]
  wire [7:0] _GEN_1850 = opcode_1 == 4'hf ? _GEN_824 : _GEN_1592; // @[executor.scala 466:52]
  wire [7:0] _GEN_1851 = opcode_1 == 4'hf ? _GEN_825 : _GEN_1593; // @[executor.scala 466:52]
  wire [7:0] _GEN_1852 = opcode_1 == 4'hf ? _GEN_826 : _GEN_1594; // @[executor.scala 466:52]
  wire [7:0] _GEN_1853 = opcode_1 == 4'hf ? _GEN_827 : _GEN_1595; // @[executor.scala 466:52]
  wire [7:0] _GEN_1854 = opcode_1 == 4'hf ? _GEN_828 : _GEN_1596; // @[executor.scala 466:52]
  wire [7:0] _GEN_1855 = opcode_1 == 4'hf ? _GEN_829 : _GEN_1597; // @[executor.scala 466:52]
  wire [7:0] _GEN_1856 = opcode_1 == 4'hf ? _GEN_830 : _GEN_1598; // @[executor.scala 466:52]
  wire [7:0] _GEN_1857 = opcode_1 == 4'hf ? _GEN_831 : _GEN_1599; // @[executor.scala 466:52]
  wire [7:0] _GEN_1858 = opcode_1 == 4'hf ? _GEN_832 : _GEN_1600; // @[executor.scala 466:52]
  wire [7:0] _GEN_1859 = opcode_1 == 4'hf ? _GEN_833 : _GEN_1601; // @[executor.scala 466:52]
  wire [7:0] _GEN_1860 = opcode_1 == 4'hf ? _GEN_834 : _GEN_1602; // @[executor.scala 466:52]
  wire [7:0] _GEN_1861 = opcode_1 == 4'hf ? _GEN_835 : _GEN_1603; // @[executor.scala 466:52]
  wire [7:0] _GEN_1862 = opcode_1 == 4'hf ? _GEN_836 : _GEN_1604; // @[executor.scala 466:52]
  wire [7:0] _GEN_1863 = opcode_1 == 4'hf ? _GEN_837 : _GEN_1605; // @[executor.scala 466:52]
  wire [7:0] _GEN_1864 = opcode_1 == 4'hf ? _GEN_838 : _GEN_1606; // @[executor.scala 466:52]
  wire [7:0] _GEN_1865 = opcode_1 == 4'hf ? _GEN_839 : _GEN_1607; // @[executor.scala 466:52]
  wire [7:0] _GEN_1866 = opcode_1 == 4'hf ? _GEN_840 : _GEN_1608; // @[executor.scala 466:52]
  wire [7:0] _GEN_1867 = opcode_1 == 4'hf ? _GEN_841 : _GEN_1609; // @[executor.scala 466:52]
  wire [7:0] _GEN_1868 = opcode_1 == 4'hf ? _GEN_842 : _GEN_1610; // @[executor.scala 466:52]
  wire [7:0] _GEN_1869 = opcode_1 == 4'hf ? _GEN_843 : _GEN_1611; // @[executor.scala 466:52]
  wire [7:0] _GEN_1870 = opcode_1 == 4'hf ? _GEN_844 : _GEN_1612; // @[executor.scala 466:52]
  wire [7:0] _GEN_1871 = opcode_1 == 4'hf ? _GEN_845 : _GEN_1613; // @[executor.scala 466:52]
  wire [7:0] _GEN_1872 = opcode_1 == 4'hf ? _GEN_846 : _GEN_1614; // @[executor.scala 466:52]
  wire [7:0] _GEN_1873 = opcode_1 == 4'hf ? _GEN_847 : _GEN_1615; // @[executor.scala 466:52]
  wire [7:0] _GEN_1874 = opcode_1 == 4'hf ? _GEN_848 : _GEN_1616; // @[executor.scala 466:52]
  wire [7:0] _GEN_1875 = opcode_1 == 4'hf ? _GEN_849 : _GEN_1617; // @[executor.scala 466:52]
  wire [7:0] _GEN_1876 = opcode_1 == 4'hf ? _GEN_850 : _GEN_1618; // @[executor.scala 466:52]
  wire [7:0] _GEN_1877 = opcode_1 == 4'hf ? _GEN_851 : _GEN_1619; // @[executor.scala 466:52]
  wire [7:0] _GEN_1878 = opcode_1 == 4'hf ? _GEN_852 : _GEN_1620; // @[executor.scala 466:52]
  wire [7:0] _GEN_1879 = opcode_1 == 4'hf ? _GEN_853 : _GEN_1621; // @[executor.scala 466:52]
  wire [7:0] _GEN_1880 = opcode_1 == 4'hf ? _GEN_854 : _GEN_1622; // @[executor.scala 466:52]
  wire [7:0] _GEN_1881 = opcode_1 == 4'hf ? _GEN_855 : _GEN_1623; // @[executor.scala 466:52]
  wire [7:0] _GEN_1882 = opcode_1 == 4'hf ? _GEN_856 : _GEN_1624; // @[executor.scala 466:52]
  wire [7:0] _GEN_1883 = opcode_1 == 4'hf ? _GEN_857 : _GEN_1625; // @[executor.scala 466:52]
  wire [7:0] _GEN_1884 = opcode_1 == 4'hf ? _GEN_858 : _GEN_1626; // @[executor.scala 466:52]
  wire [7:0] _GEN_1885 = opcode_1 == 4'hf ? _GEN_859 : _GEN_1627; // @[executor.scala 466:52]
  wire [7:0] _GEN_1886 = opcode_1 == 4'hf ? _GEN_860 : _GEN_1628; // @[executor.scala 466:52]
  wire [7:0] _GEN_1887 = opcode_1 == 4'hf ? _GEN_861 : _GEN_1629; // @[executor.scala 466:52]
  wire [7:0] _GEN_1888 = opcode_1 == 4'hf ? _GEN_862 : _GEN_1630; // @[executor.scala 466:52]
  wire [7:0] _GEN_1889 = opcode_1 == 4'hf ? _GEN_863 : _GEN_1631; // @[executor.scala 466:52]
  wire [7:0] _GEN_1890 = opcode_1 == 4'hf ? _GEN_864 : _GEN_1632; // @[executor.scala 466:52]
  wire [7:0] _GEN_1891 = opcode_1 == 4'hf ? _GEN_865 : _GEN_1633; // @[executor.scala 466:52]
  wire [7:0] _GEN_1892 = opcode_1 == 4'hf ? _GEN_866 : _GEN_1634; // @[executor.scala 466:52]
  wire [7:0] _GEN_1893 = opcode_1 == 4'hf ? _GEN_867 : _GEN_1635; // @[executor.scala 466:52]
  wire [7:0] _GEN_1894 = opcode_1 == 4'hf ? _GEN_868 : _GEN_1636; // @[executor.scala 466:52]
  wire [7:0] _GEN_1895 = opcode_1 == 4'hf ? _GEN_869 : _GEN_1637; // @[executor.scala 466:52]
  wire [7:0] _GEN_1896 = opcode_1 == 4'hf ? _GEN_870 : _GEN_1638; // @[executor.scala 466:52]
  wire [7:0] _GEN_1897 = opcode_1 == 4'hf ? _GEN_871 : _GEN_1639; // @[executor.scala 466:52]
  wire [7:0] _GEN_1898 = opcode_1 == 4'hf ? _GEN_872 : _GEN_1640; // @[executor.scala 466:52]
  wire [7:0] _GEN_1899 = opcode_1 == 4'hf ? _GEN_873 : _GEN_1641; // @[executor.scala 466:52]
  wire [7:0] _GEN_1900 = opcode_1 == 4'hf ? _GEN_874 : _GEN_1642; // @[executor.scala 466:52]
  wire [7:0] _GEN_1901 = opcode_1 == 4'hf ? _GEN_875 : _GEN_1643; // @[executor.scala 466:52]
  wire [7:0] _GEN_1902 = opcode_1 == 4'hf ? _GEN_876 : _GEN_1644; // @[executor.scala 466:52]
  wire [7:0] _GEN_1903 = opcode_1 == 4'hf ? _GEN_877 : _GEN_1645; // @[executor.scala 466:52]
  wire [7:0] _GEN_1904 = opcode_1 == 4'hf ? _GEN_878 : _GEN_1646; // @[executor.scala 466:52]
  wire [7:0] _GEN_1905 = opcode_1 == 4'hf ? _GEN_879 : _GEN_1647; // @[executor.scala 466:52]
  wire [7:0] _GEN_1906 = opcode_1 == 4'hf ? _GEN_880 : _GEN_1648; // @[executor.scala 466:52]
  wire [7:0] _GEN_1907 = opcode_1 == 4'hf ? _GEN_881 : _GEN_1649; // @[executor.scala 466:52]
  wire [7:0] _GEN_1908 = opcode_1 == 4'hf ? _GEN_882 : _GEN_1650; // @[executor.scala 466:52]
  wire [7:0] _GEN_1909 = opcode_1 == 4'hf ? _GEN_883 : _GEN_1651; // @[executor.scala 466:52]
  wire [7:0] _GEN_1910 = opcode_1 == 4'hf ? _GEN_884 : _GEN_1652; // @[executor.scala 466:52]
  wire [7:0] _GEN_1911 = opcode_1 == 4'hf ? _GEN_885 : _GEN_1653; // @[executor.scala 466:52]
  wire [7:0] _GEN_1912 = opcode_1 == 4'hf ? _GEN_886 : _GEN_1654; // @[executor.scala 466:52]
  wire [7:0] _GEN_1913 = opcode_1 == 4'hf ? _GEN_887 : _GEN_1655; // @[executor.scala 466:52]
  wire [7:0] _GEN_1914 = opcode_1 == 4'hf ? _GEN_888 : _GEN_1656; // @[executor.scala 466:52]
  wire [7:0] _GEN_1915 = opcode_1 == 4'hf ? _GEN_889 : _GEN_1657; // @[executor.scala 466:52]
  wire [7:0] _GEN_1916 = opcode_1 == 4'hf ? _GEN_890 : _GEN_1658; // @[executor.scala 466:52]
  wire [7:0] _GEN_1917 = opcode_1 == 4'hf ? _GEN_891 : _GEN_1659; // @[executor.scala 466:52]
  wire [7:0] _GEN_1918 = opcode_1 == 4'hf ? _GEN_892 : _GEN_1660; // @[executor.scala 466:52]
  wire [7:0] _GEN_1919 = opcode_1 == 4'hf ? _GEN_893 : _GEN_1661; // @[executor.scala 466:52]
  wire [7:0] _GEN_1920 = opcode_1 == 4'hf ? _GEN_894 : _GEN_1662; // @[executor.scala 466:52]
  wire [7:0] _GEN_1921 = opcode_1 == 4'hf ? _GEN_895 : _GEN_1663; // @[executor.scala 466:52]
  wire [7:0] _GEN_1922 = opcode_1 == 4'hf ? _GEN_896 : _GEN_1664; // @[executor.scala 466:52]
  wire [7:0] _GEN_1923 = opcode_1 == 4'hf ? _GEN_897 : _GEN_1665; // @[executor.scala 466:52]
  wire [7:0] _GEN_1924 = opcode_1 == 4'hf ? _GEN_898 : _GEN_1666; // @[executor.scala 466:52]
  wire [7:0] _GEN_1925 = opcode_1 == 4'hf ? _GEN_899 : _GEN_1667; // @[executor.scala 466:52]
  wire [7:0] _GEN_1926 = opcode_1 == 4'hf ? _GEN_900 : _GEN_1668; // @[executor.scala 466:52]
  wire [7:0] _GEN_1927 = opcode_1 == 4'hf ? _GEN_901 : _GEN_1669; // @[executor.scala 466:52]
  wire [7:0] _GEN_1928 = opcode_1 == 4'hf ? _GEN_902 : _GEN_1670; // @[executor.scala 466:52]
  wire [7:0] _GEN_1929 = opcode_1 == 4'hf ? _GEN_903 : _GEN_1671; // @[executor.scala 466:52]
  wire [7:0] _GEN_1930 = opcode_1 == 4'hf ? _GEN_904 : _GEN_1672; // @[executor.scala 466:52]
  wire [7:0] _GEN_1931 = opcode_1 == 4'hf ? _GEN_905 : _GEN_1673; // @[executor.scala 466:52]
  wire [7:0] _GEN_1932 = opcode_1 == 4'hf ? _GEN_906 : _GEN_1674; // @[executor.scala 466:52]
  wire [7:0] _GEN_1933 = opcode_1 == 4'hf ? _GEN_907 : _GEN_1675; // @[executor.scala 466:52]
  wire [7:0] _GEN_1934 = opcode_1 == 4'hf ? _GEN_908 : _GEN_1676; // @[executor.scala 466:52]
  wire [7:0] _GEN_1935 = opcode_1 == 4'hf ? _GEN_909 : _GEN_1677; // @[executor.scala 466:52]
  wire [7:0] _GEN_1936 = opcode_1 == 4'hf ? _GEN_910 : _GEN_1678; // @[executor.scala 466:52]
  wire [7:0] _GEN_1937 = opcode_1 == 4'hf ? _GEN_911 : _GEN_1679; // @[executor.scala 466:52]
  wire [7:0] _GEN_1938 = opcode_1 == 4'hf ? _GEN_912 : _GEN_1680; // @[executor.scala 466:52]
  wire [7:0] _GEN_1939 = opcode_1 == 4'hf ? _GEN_913 : _GEN_1681; // @[executor.scala 466:52]
  wire [7:0] _GEN_1940 = opcode_1 == 4'hf ? _GEN_914 : _GEN_1682; // @[executor.scala 466:52]
  wire [7:0] _GEN_1941 = opcode_1 == 4'hf ? _GEN_915 : _GEN_1683; // @[executor.scala 466:52]
  wire [7:0] _GEN_1942 = opcode_1 == 4'hf ? _GEN_916 : _GEN_1684; // @[executor.scala 466:52]
  wire [7:0] _GEN_1943 = opcode_1 == 4'hf ? _GEN_917 : _GEN_1685; // @[executor.scala 466:52]
  wire [7:0] _GEN_1944 = opcode_1 == 4'hf ? _GEN_918 : _GEN_1686; // @[executor.scala 466:52]
  wire [7:0] _GEN_1945 = opcode_1 == 4'hf ? _GEN_919 : _GEN_1687; // @[executor.scala 466:52]
  wire [7:0] _GEN_1946 = opcode_1 == 4'hf ? _GEN_920 : _GEN_1688; // @[executor.scala 466:52]
  wire [7:0] _GEN_1947 = opcode_1 == 4'hf ? _GEN_921 : _GEN_1689; // @[executor.scala 466:52]
  wire [7:0] _GEN_1948 = opcode_1 == 4'hf ? _GEN_922 : _GEN_1690; // @[executor.scala 466:52]
  wire [7:0] _GEN_1949 = opcode_1 == 4'hf ? _GEN_923 : _GEN_1691; // @[executor.scala 466:52]
  wire [7:0] _GEN_1950 = opcode_1 == 4'hf ? _GEN_924 : _GEN_1692; // @[executor.scala 466:52]
  wire [7:0] _GEN_1951 = opcode_1 == 4'hf ? _GEN_925 : _GEN_1693; // @[executor.scala 466:52]
  wire [7:0] _GEN_1952 = opcode_1 == 4'hf ? _GEN_926 : _GEN_1694; // @[executor.scala 466:52]
  wire [7:0] _GEN_1953 = opcode_1 == 4'hf ? _GEN_927 : _GEN_1695; // @[executor.scala 466:52]
  wire [7:0] _GEN_1954 = opcode_1 == 4'hf ? _GEN_928 : _GEN_1696; // @[executor.scala 466:52]
  wire [7:0] _GEN_1955 = opcode_1 == 4'hf ? _GEN_929 : _GEN_1697; // @[executor.scala 466:52]
  wire [7:0] _GEN_1956 = opcode_1 == 4'hf ? _GEN_930 : _GEN_1698; // @[executor.scala 466:52]
  wire [7:0] _GEN_1957 = opcode_1 == 4'hf ? _GEN_931 : _GEN_1699; // @[executor.scala 466:52]
  wire [7:0] _GEN_1958 = opcode_1 == 4'hf ? _GEN_932 : _GEN_1700; // @[executor.scala 466:52]
  wire [7:0] _GEN_1959 = opcode_1 == 4'hf ? _GEN_933 : _GEN_1701; // @[executor.scala 466:52]
  wire [7:0] _GEN_1960 = opcode_1 == 4'hf ? _GEN_934 : _GEN_1702; // @[executor.scala 466:52]
  wire [7:0] _GEN_1961 = opcode_1 == 4'hf ? _GEN_935 : _GEN_1703; // @[executor.scala 466:52]
  wire [7:0] _GEN_1962 = opcode_1 == 4'hf ? _GEN_936 : _GEN_1704; // @[executor.scala 466:52]
  wire [7:0] _GEN_1963 = opcode_1 == 4'hf ? _GEN_937 : _GEN_1705; // @[executor.scala 466:52]
  wire [7:0] _GEN_1964 = opcode_1 == 4'hf ? _GEN_938 : _GEN_1706; // @[executor.scala 466:52]
  wire [7:0] _GEN_1965 = opcode_1 == 4'hf ? _GEN_939 : _GEN_1707; // @[executor.scala 466:52]
  wire [7:0] _GEN_1966 = opcode_1 == 4'hf ? _GEN_940 : _GEN_1708; // @[executor.scala 466:52]
  wire [7:0] _GEN_1967 = opcode_1 == 4'hf ? _GEN_941 : _GEN_1709; // @[executor.scala 466:52]
  wire [7:0] _GEN_1968 = opcode_1 == 4'hf ? _GEN_942 : _GEN_1710; // @[executor.scala 466:52]
  wire [7:0] _GEN_1969 = opcode_1 == 4'hf ? _GEN_943 : _GEN_1711; // @[executor.scala 466:52]
  wire [7:0] _GEN_1970 = opcode_1 == 4'hf ? _GEN_944 : _GEN_1712; // @[executor.scala 466:52]
  wire [7:0] _GEN_1971 = opcode_1 == 4'hf ? _GEN_945 : _GEN_1713; // @[executor.scala 466:52]
  wire [7:0] _GEN_1972 = opcode_1 == 4'hf ? _GEN_946 : _GEN_1714; // @[executor.scala 466:52]
  wire [7:0] _GEN_1973 = opcode_1 == 4'hf ? _GEN_947 : _GEN_1715; // @[executor.scala 466:52]
  wire [7:0] _GEN_1974 = opcode_1 == 4'hf ? _GEN_948 : _GEN_1716; // @[executor.scala 466:52]
  wire [7:0] _GEN_1975 = opcode_1 == 4'hf ? _GEN_949 : _GEN_1717; // @[executor.scala 466:52]
  wire [7:0] _GEN_1976 = opcode_1 == 4'hf ? _GEN_950 : _GEN_1718; // @[executor.scala 466:52]
  wire [7:0] _GEN_1977 = opcode_1 == 4'hf ? _GEN_951 : _GEN_1719; // @[executor.scala 466:52]
  wire [7:0] _GEN_1978 = opcode_1 == 4'hf ? _GEN_952 : _GEN_1720; // @[executor.scala 466:52]
  wire [7:0] _GEN_1979 = opcode_1 == 4'hf ? _GEN_953 : _GEN_1721; // @[executor.scala 466:52]
  wire [7:0] _GEN_1980 = opcode_1 == 4'hf ? _GEN_954 : _GEN_1722; // @[executor.scala 466:52]
  wire [7:0] _GEN_1981 = opcode_1 == 4'hf ? _GEN_955 : _GEN_1723; // @[executor.scala 466:52]
  wire [7:0] _GEN_1982 = opcode_1 == 4'hf ? _GEN_956 : _GEN_1724; // @[executor.scala 466:52]
  wire [7:0] _GEN_1983 = opcode_1 == 4'hf ? _GEN_957 : _GEN_1725; // @[executor.scala 466:52]
  wire [7:0] _GEN_1984 = opcode_1 == 4'hf ? _GEN_958 : _GEN_1726; // @[executor.scala 466:52]
  wire [7:0] _GEN_1985 = opcode_1 == 4'hf ? _GEN_959 : _GEN_1727; // @[executor.scala 466:52]
  wire [7:0] _GEN_1986 = opcode_1 == 4'hf ? _GEN_960 : _GEN_1728; // @[executor.scala 466:52]
  wire [7:0] _GEN_1987 = opcode_1 == 4'hf ? _GEN_961 : _GEN_1729; // @[executor.scala 466:52]
  wire [7:0] _GEN_1988 = opcode_1 == 4'hf ? _GEN_962 : _GEN_1730; // @[executor.scala 466:52]
  wire [7:0] _GEN_1989 = opcode_1 == 4'hf ? _GEN_963 : _GEN_1731; // @[executor.scala 466:52]
  wire [7:0] _GEN_1990 = opcode_1 == 4'hf ? _GEN_964 : _GEN_1732; // @[executor.scala 466:52]
  wire [7:0] _GEN_1991 = opcode_1 == 4'hf ? _GEN_965 : _GEN_1733; // @[executor.scala 466:52]
  wire [7:0] _GEN_1992 = opcode_1 == 4'hf ? _GEN_966 : _GEN_1734; // @[executor.scala 466:52]
  wire [7:0] _GEN_1993 = opcode_1 == 4'hf ? _GEN_967 : _GEN_1735; // @[executor.scala 466:52]
  wire [7:0] _GEN_1994 = opcode_1 == 4'hf ? _GEN_968 : _GEN_1736; // @[executor.scala 466:52]
  wire [7:0] _GEN_1995 = opcode_1 == 4'hf ? _GEN_969 : _GEN_1737; // @[executor.scala 466:52]
  wire [7:0] _GEN_1996 = opcode_1 == 4'hf ? _GEN_970 : _GEN_1738; // @[executor.scala 466:52]
  wire [7:0] _GEN_1997 = opcode_1 == 4'hf ? _GEN_971 : _GEN_1739; // @[executor.scala 466:52]
  wire [7:0] _GEN_1998 = opcode_1 == 4'hf ? _GEN_972 : _GEN_1740; // @[executor.scala 466:52]
  wire [7:0] _GEN_1999 = opcode_1 == 4'hf ? _GEN_973 : _GEN_1741; // @[executor.scala 466:52]
  wire [7:0] _GEN_2000 = opcode_1 == 4'hf ? _GEN_974 : _GEN_1742; // @[executor.scala 466:52]
  wire [7:0] _GEN_2001 = opcode_1 == 4'hf ? _GEN_975 : _GEN_1743; // @[executor.scala 466:52]
  wire [7:0] _GEN_2002 = opcode_1 == 4'hf ? _GEN_976 : _GEN_1744; // @[executor.scala 466:52]
  wire [7:0] _GEN_2003 = opcode_1 == 4'hf ? _GEN_977 : _GEN_1745; // @[executor.scala 466:52]
  wire [7:0] _GEN_2004 = opcode_1 == 4'hf ? _GEN_978 : _GEN_1746; // @[executor.scala 466:52]
  wire [7:0] _GEN_2005 = opcode_1 == 4'hf ? _GEN_979 : _GEN_1747; // @[executor.scala 466:52]
  wire [7:0] _GEN_2006 = opcode_1 == 4'hf ? _GEN_980 : _GEN_1748; // @[executor.scala 466:52]
  wire [7:0] _GEN_2007 = opcode_1 == 4'hf ? _GEN_981 : _GEN_1749; // @[executor.scala 466:52]
  wire [7:0] _GEN_2008 = opcode_1 == 4'hf ? _GEN_982 : _GEN_1750; // @[executor.scala 466:52]
  wire [7:0] _GEN_2009 = opcode_1 == 4'hf ? _GEN_983 : _GEN_1751; // @[executor.scala 466:52]
  wire [7:0] _GEN_2010 = opcode_1 == 4'hf ? _GEN_984 : _GEN_1752; // @[executor.scala 466:52]
  wire [7:0] _GEN_2011 = opcode_1 == 4'hf ? _GEN_985 : _GEN_1753; // @[executor.scala 466:52]
  wire [7:0] _GEN_2012 = opcode_1 == 4'hf ? _GEN_986 : _GEN_1754; // @[executor.scala 466:52]
  wire [7:0] _GEN_2013 = opcode_1 == 4'hf ? _GEN_987 : _GEN_1755; // @[executor.scala 466:52]
  wire [7:0] _GEN_2014 = opcode_1 == 4'hf ? _GEN_988 : _GEN_1756; // @[executor.scala 466:52]
  wire [7:0] _GEN_2015 = opcode_1 == 4'hf ? _GEN_989 : _GEN_1757; // @[executor.scala 466:52]
  wire [7:0] _GEN_2016 = opcode_1 == 4'hf ? _GEN_990 : _GEN_1758; // @[executor.scala 466:52]
  wire [7:0] _GEN_2017 = opcode_1 == 4'hf ? _GEN_991 : _GEN_1759; // @[executor.scala 466:52]
  wire [7:0] _GEN_2018 = opcode_1 == 4'hf ? _GEN_992 : _GEN_1760; // @[executor.scala 466:52]
  wire [7:0] _GEN_2019 = opcode_1 == 4'hf ? _GEN_993 : _GEN_1761; // @[executor.scala 466:52]
  wire [7:0] _GEN_2020 = opcode_1 == 4'hf ? _GEN_994 : _GEN_1762; // @[executor.scala 466:52]
  wire [7:0] _GEN_2021 = opcode_1 == 4'hf ? _GEN_995 : _GEN_1763; // @[executor.scala 466:52]
  wire [7:0] _GEN_2022 = opcode_1 == 4'hf ? _GEN_996 : _GEN_1764; // @[executor.scala 466:52]
  wire [7:0] _GEN_2023 = opcode_1 == 4'hf ? _GEN_997 : _GEN_1765; // @[executor.scala 466:52]
  wire [7:0] _GEN_2024 = opcode_1 == 4'hf ? _GEN_998 : _GEN_1766; // @[executor.scala 466:52]
  wire [7:0] _GEN_2025 = opcode_1 == 4'hf ? _GEN_999 : _GEN_1767; // @[executor.scala 466:52]
  wire [7:0] _GEN_2026 = opcode_1 == 4'hf ? _GEN_1000 : _GEN_1768; // @[executor.scala 466:52]
  wire [7:0] _GEN_2027 = opcode_1 == 4'hf ? _GEN_1001 : _GEN_1769; // @[executor.scala 466:52]
  wire [7:0] _GEN_2028 = opcode_1 == 4'hf ? _GEN_1002 : _GEN_1770; // @[executor.scala 466:52]
  wire [7:0] _GEN_2029 = opcode_1 == 4'hf ? _GEN_1003 : _GEN_1771; // @[executor.scala 466:52]
  wire [7:0] _GEN_2030 = opcode_1 == 4'hf ? _GEN_1004 : _GEN_1772; // @[executor.scala 466:52]
  wire [7:0] _GEN_2031 = opcode_1 == 4'hf ? _GEN_1005 : _GEN_1773; // @[executor.scala 466:52]
  wire [7:0] _GEN_2032 = opcode_1 == 4'hf ? _GEN_1006 : _GEN_1774; // @[executor.scala 466:52]
  wire [7:0] _GEN_2033 = opcode_1 == 4'hf ? _GEN_1007 : _GEN_1775; // @[executor.scala 466:52]
  wire [7:0] _GEN_2034 = opcode_1 == 4'hf ? _GEN_1008 : _GEN_1776; // @[executor.scala 466:52]
  wire [7:0] _GEN_2035 = opcode_1 == 4'hf ? _GEN_1009 : _GEN_1777; // @[executor.scala 466:52]
  wire [7:0] _GEN_2036 = opcode_1 == 4'hf ? _GEN_1010 : _GEN_1778; // @[executor.scala 466:52]
  wire [7:0] _GEN_2037 = opcode_1 == 4'hf ? _GEN_1011 : _GEN_1779; // @[executor.scala 466:52]
  wire [7:0] _GEN_2038 = opcode_1 == 4'hf ? _GEN_1012 : _GEN_1780; // @[executor.scala 466:52]
  wire [7:0] _GEN_2039 = opcode_1 == 4'hf ? _GEN_1013 : _GEN_1781; // @[executor.scala 466:52]
  wire [7:0] _GEN_2040 = opcode_1 == 4'hf ? _GEN_1014 : _GEN_1782; // @[executor.scala 466:52]
  wire [7:0] _GEN_2041 = opcode_1 == 4'hf ? _GEN_1015 : _GEN_1783; // @[executor.scala 466:52]
  wire [7:0] _GEN_2042 = opcode_1 == 4'hf ? _GEN_1016 : _GEN_1784; // @[executor.scala 466:52]
  wire [7:0] _GEN_2043 = opcode_1 == 4'hf ? _GEN_1017 : _GEN_1785; // @[executor.scala 466:52]
  wire [7:0] _GEN_2044 = opcode_1 == 4'hf ? _GEN_1018 : _GEN_1786; // @[executor.scala 466:52]
  wire [7:0] _GEN_2045 = opcode_1 == 4'hf ? _GEN_1019 : _GEN_1787; // @[executor.scala 466:52]
  wire [7:0] _GEN_2046 = opcode_1 == 4'hf ? _GEN_1020 : _GEN_1788; // @[executor.scala 466:52]
  wire [7:0] _GEN_2047 = opcode_1 == 4'hf ? _GEN_1021 : _GEN_1789; // @[executor.scala 466:52]
  wire [7:0] _GEN_2048 = opcode_1 == 4'hf ? _GEN_1022 : _GEN_1790; // @[executor.scala 466:52]
  wire [7:0] _GEN_2049 = opcode_1 == 4'hf ? _GEN_1023 : _GEN_1791; // @[executor.scala 466:52]
  wire [7:0] _GEN_2050 = opcode_1 == 4'hf ? _GEN_1024 : _GEN_1792; // @[executor.scala 466:52]
  wire [7:0] _GEN_2051 = opcode_1 == 4'hf ? _GEN_1025 : _GEN_1793; // @[executor.scala 466:52]
  wire [3:0] opcode_2 = vliw_2[31:28]; // @[primitive.scala 9:44]
  wire [7:0] _GEN_4490 = {{2'd0}, dst_offset_2}; // @[executor.scala 473:49]
  wire [7:0] byte_512 = field_2[7:0]; // @[executor.scala 475:56]
  wire [7:0] _GEN_2052 = mask_2[0] ? byte_512 : _GEN_1796; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] byte_513 = field_2[15:8]; // @[executor.scala 475:56]
  wire [7:0] _GEN_2053 = mask_2[1] ? byte_513 : _GEN_1797; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] byte_514 = field_2[23:16]; // @[executor.scala 475:56]
  wire [7:0] _GEN_2054 = mask_2[2] ? byte_514 : _GEN_1798; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] byte_515 = field_2[31:24]; // @[executor.scala 475:56]
  wire [7:0] _GEN_2055 = mask_2[3] ? byte_515 : _GEN_1799; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2056 = _GEN_4490 == 8'h0 ? _GEN_2052 : _GEN_1796; // @[executor.scala 473:84]
  wire [7:0] _GEN_2057 = _GEN_4490 == 8'h0 ? _GEN_2053 : _GEN_1797; // @[executor.scala 473:84]
  wire [7:0] _GEN_2058 = _GEN_4490 == 8'h0 ? _GEN_2054 : _GEN_1798; // @[executor.scala 473:84]
  wire [7:0] _GEN_2059 = _GEN_4490 == 8'h0 ? _GEN_2055 : _GEN_1799; // @[executor.scala 473:84]
  wire [7:0] _GEN_2060 = mask_2[0] ? byte_512 : _GEN_1800; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2061 = mask_2[1] ? byte_513 : _GEN_1801; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2062 = mask_2[2] ? byte_514 : _GEN_1802; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2063 = mask_2[3] ? byte_515 : _GEN_1803; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2064 = _GEN_4490 == 8'h1 ? _GEN_2060 : _GEN_1800; // @[executor.scala 473:84]
  wire [7:0] _GEN_2065 = _GEN_4490 == 8'h1 ? _GEN_2061 : _GEN_1801; // @[executor.scala 473:84]
  wire [7:0] _GEN_2066 = _GEN_4490 == 8'h1 ? _GEN_2062 : _GEN_1802; // @[executor.scala 473:84]
  wire [7:0] _GEN_2067 = _GEN_4490 == 8'h1 ? _GEN_2063 : _GEN_1803; // @[executor.scala 473:84]
  wire [7:0] _GEN_2068 = mask_2[0] ? byte_512 : _GEN_1804; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2069 = mask_2[1] ? byte_513 : _GEN_1805; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2070 = mask_2[2] ? byte_514 : _GEN_1806; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2071 = mask_2[3] ? byte_515 : _GEN_1807; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2072 = _GEN_4490 == 8'h2 ? _GEN_2068 : _GEN_1804; // @[executor.scala 473:84]
  wire [7:0] _GEN_2073 = _GEN_4490 == 8'h2 ? _GEN_2069 : _GEN_1805; // @[executor.scala 473:84]
  wire [7:0] _GEN_2074 = _GEN_4490 == 8'h2 ? _GEN_2070 : _GEN_1806; // @[executor.scala 473:84]
  wire [7:0] _GEN_2075 = _GEN_4490 == 8'h2 ? _GEN_2071 : _GEN_1807; // @[executor.scala 473:84]
  wire [7:0] _GEN_2076 = mask_2[0] ? byte_512 : _GEN_1808; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2077 = mask_2[1] ? byte_513 : _GEN_1809; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2078 = mask_2[2] ? byte_514 : _GEN_1810; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2079 = mask_2[3] ? byte_515 : _GEN_1811; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2080 = _GEN_4490 == 8'h3 ? _GEN_2076 : _GEN_1808; // @[executor.scala 473:84]
  wire [7:0] _GEN_2081 = _GEN_4490 == 8'h3 ? _GEN_2077 : _GEN_1809; // @[executor.scala 473:84]
  wire [7:0] _GEN_2082 = _GEN_4490 == 8'h3 ? _GEN_2078 : _GEN_1810; // @[executor.scala 473:84]
  wire [7:0] _GEN_2083 = _GEN_4490 == 8'h3 ? _GEN_2079 : _GEN_1811; // @[executor.scala 473:84]
  wire [7:0] _GEN_2084 = mask_2[0] ? byte_512 : _GEN_1812; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2085 = mask_2[1] ? byte_513 : _GEN_1813; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2086 = mask_2[2] ? byte_514 : _GEN_1814; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2087 = mask_2[3] ? byte_515 : _GEN_1815; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2088 = _GEN_4490 == 8'h4 ? _GEN_2084 : _GEN_1812; // @[executor.scala 473:84]
  wire [7:0] _GEN_2089 = _GEN_4490 == 8'h4 ? _GEN_2085 : _GEN_1813; // @[executor.scala 473:84]
  wire [7:0] _GEN_2090 = _GEN_4490 == 8'h4 ? _GEN_2086 : _GEN_1814; // @[executor.scala 473:84]
  wire [7:0] _GEN_2091 = _GEN_4490 == 8'h4 ? _GEN_2087 : _GEN_1815; // @[executor.scala 473:84]
  wire [7:0] _GEN_2092 = mask_2[0] ? byte_512 : _GEN_1816; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2093 = mask_2[1] ? byte_513 : _GEN_1817; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2094 = mask_2[2] ? byte_514 : _GEN_1818; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2095 = mask_2[3] ? byte_515 : _GEN_1819; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2096 = _GEN_4490 == 8'h5 ? _GEN_2092 : _GEN_1816; // @[executor.scala 473:84]
  wire [7:0] _GEN_2097 = _GEN_4490 == 8'h5 ? _GEN_2093 : _GEN_1817; // @[executor.scala 473:84]
  wire [7:0] _GEN_2098 = _GEN_4490 == 8'h5 ? _GEN_2094 : _GEN_1818; // @[executor.scala 473:84]
  wire [7:0] _GEN_2099 = _GEN_4490 == 8'h5 ? _GEN_2095 : _GEN_1819; // @[executor.scala 473:84]
  wire [7:0] _GEN_2100 = mask_2[0] ? byte_512 : _GEN_1820; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2101 = mask_2[1] ? byte_513 : _GEN_1821; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2102 = mask_2[2] ? byte_514 : _GEN_1822; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2103 = mask_2[3] ? byte_515 : _GEN_1823; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2104 = _GEN_4490 == 8'h6 ? _GEN_2100 : _GEN_1820; // @[executor.scala 473:84]
  wire [7:0] _GEN_2105 = _GEN_4490 == 8'h6 ? _GEN_2101 : _GEN_1821; // @[executor.scala 473:84]
  wire [7:0] _GEN_2106 = _GEN_4490 == 8'h6 ? _GEN_2102 : _GEN_1822; // @[executor.scala 473:84]
  wire [7:0] _GEN_2107 = _GEN_4490 == 8'h6 ? _GEN_2103 : _GEN_1823; // @[executor.scala 473:84]
  wire [7:0] _GEN_2108 = mask_2[0] ? byte_512 : _GEN_1824; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2109 = mask_2[1] ? byte_513 : _GEN_1825; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2110 = mask_2[2] ? byte_514 : _GEN_1826; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2111 = mask_2[3] ? byte_515 : _GEN_1827; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2112 = _GEN_4490 == 8'h7 ? _GEN_2108 : _GEN_1824; // @[executor.scala 473:84]
  wire [7:0] _GEN_2113 = _GEN_4490 == 8'h7 ? _GEN_2109 : _GEN_1825; // @[executor.scala 473:84]
  wire [7:0] _GEN_2114 = _GEN_4490 == 8'h7 ? _GEN_2110 : _GEN_1826; // @[executor.scala 473:84]
  wire [7:0] _GEN_2115 = _GEN_4490 == 8'h7 ? _GEN_2111 : _GEN_1827; // @[executor.scala 473:84]
  wire [7:0] _GEN_2116 = mask_2[0] ? byte_512 : _GEN_1828; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2117 = mask_2[1] ? byte_513 : _GEN_1829; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2118 = mask_2[2] ? byte_514 : _GEN_1830; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2119 = mask_2[3] ? byte_515 : _GEN_1831; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2120 = _GEN_4490 == 8'h8 ? _GEN_2116 : _GEN_1828; // @[executor.scala 473:84]
  wire [7:0] _GEN_2121 = _GEN_4490 == 8'h8 ? _GEN_2117 : _GEN_1829; // @[executor.scala 473:84]
  wire [7:0] _GEN_2122 = _GEN_4490 == 8'h8 ? _GEN_2118 : _GEN_1830; // @[executor.scala 473:84]
  wire [7:0] _GEN_2123 = _GEN_4490 == 8'h8 ? _GEN_2119 : _GEN_1831; // @[executor.scala 473:84]
  wire [7:0] _GEN_2124 = mask_2[0] ? byte_512 : _GEN_1832; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2125 = mask_2[1] ? byte_513 : _GEN_1833; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2126 = mask_2[2] ? byte_514 : _GEN_1834; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2127 = mask_2[3] ? byte_515 : _GEN_1835; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2128 = _GEN_4490 == 8'h9 ? _GEN_2124 : _GEN_1832; // @[executor.scala 473:84]
  wire [7:0] _GEN_2129 = _GEN_4490 == 8'h9 ? _GEN_2125 : _GEN_1833; // @[executor.scala 473:84]
  wire [7:0] _GEN_2130 = _GEN_4490 == 8'h9 ? _GEN_2126 : _GEN_1834; // @[executor.scala 473:84]
  wire [7:0] _GEN_2131 = _GEN_4490 == 8'h9 ? _GEN_2127 : _GEN_1835; // @[executor.scala 473:84]
  wire [7:0] _GEN_2132 = mask_2[0] ? byte_512 : _GEN_1836; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2133 = mask_2[1] ? byte_513 : _GEN_1837; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2134 = mask_2[2] ? byte_514 : _GEN_1838; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2135 = mask_2[3] ? byte_515 : _GEN_1839; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2136 = _GEN_4490 == 8'ha ? _GEN_2132 : _GEN_1836; // @[executor.scala 473:84]
  wire [7:0] _GEN_2137 = _GEN_4490 == 8'ha ? _GEN_2133 : _GEN_1837; // @[executor.scala 473:84]
  wire [7:0] _GEN_2138 = _GEN_4490 == 8'ha ? _GEN_2134 : _GEN_1838; // @[executor.scala 473:84]
  wire [7:0] _GEN_2139 = _GEN_4490 == 8'ha ? _GEN_2135 : _GEN_1839; // @[executor.scala 473:84]
  wire [7:0] _GEN_2140 = mask_2[0] ? byte_512 : _GEN_1840; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2141 = mask_2[1] ? byte_513 : _GEN_1841; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2142 = mask_2[2] ? byte_514 : _GEN_1842; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2143 = mask_2[3] ? byte_515 : _GEN_1843; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2144 = _GEN_4490 == 8'hb ? _GEN_2140 : _GEN_1840; // @[executor.scala 473:84]
  wire [7:0] _GEN_2145 = _GEN_4490 == 8'hb ? _GEN_2141 : _GEN_1841; // @[executor.scala 473:84]
  wire [7:0] _GEN_2146 = _GEN_4490 == 8'hb ? _GEN_2142 : _GEN_1842; // @[executor.scala 473:84]
  wire [7:0] _GEN_2147 = _GEN_4490 == 8'hb ? _GEN_2143 : _GEN_1843; // @[executor.scala 473:84]
  wire [7:0] _GEN_2148 = mask_2[0] ? byte_512 : _GEN_1844; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2149 = mask_2[1] ? byte_513 : _GEN_1845; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2150 = mask_2[2] ? byte_514 : _GEN_1846; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2151 = mask_2[3] ? byte_515 : _GEN_1847; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2152 = _GEN_4490 == 8'hc ? _GEN_2148 : _GEN_1844; // @[executor.scala 473:84]
  wire [7:0] _GEN_2153 = _GEN_4490 == 8'hc ? _GEN_2149 : _GEN_1845; // @[executor.scala 473:84]
  wire [7:0] _GEN_2154 = _GEN_4490 == 8'hc ? _GEN_2150 : _GEN_1846; // @[executor.scala 473:84]
  wire [7:0] _GEN_2155 = _GEN_4490 == 8'hc ? _GEN_2151 : _GEN_1847; // @[executor.scala 473:84]
  wire [7:0] _GEN_2156 = mask_2[0] ? byte_512 : _GEN_1848; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2157 = mask_2[1] ? byte_513 : _GEN_1849; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2158 = mask_2[2] ? byte_514 : _GEN_1850; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2159 = mask_2[3] ? byte_515 : _GEN_1851; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2160 = _GEN_4490 == 8'hd ? _GEN_2156 : _GEN_1848; // @[executor.scala 473:84]
  wire [7:0] _GEN_2161 = _GEN_4490 == 8'hd ? _GEN_2157 : _GEN_1849; // @[executor.scala 473:84]
  wire [7:0] _GEN_2162 = _GEN_4490 == 8'hd ? _GEN_2158 : _GEN_1850; // @[executor.scala 473:84]
  wire [7:0] _GEN_2163 = _GEN_4490 == 8'hd ? _GEN_2159 : _GEN_1851; // @[executor.scala 473:84]
  wire [7:0] _GEN_2164 = mask_2[0] ? byte_512 : _GEN_1852; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2165 = mask_2[1] ? byte_513 : _GEN_1853; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2166 = mask_2[2] ? byte_514 : _GEN_1854; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2167 = mask_2[3] ? byte_515 : _GEN_1855; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2168 = _GEN_4490 == 8'he ? _GEN_2164 : _GEN_1852; // @[executor.scala 473:84]
  wire [7:0] _GEN_2169 = _GEN_4490 == 8'he ? _GEN_2165 : _GEN_1853; // @[executor.scala 473:84]
  wire [7:0] _GEN_2170 = _GEN_4490 == 8'he ? _GEN_2166 : _GEN_1854; // @[executor.scala 473:84]
  wire [7:0] _GEN_2171 = _GEN_4490 == 8'he ? _GEN_2167 : _GEN_1855; // @[executor.scala 473:84]
  wire [7:0] _GEN_2172 = mask_2[0] ? byte_512 : _GEN_1856; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2173 = mask_2[1] ? byte_513 : _GEN_1857; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2174 = mask_2[2] ? byte_514 : _GEN_1858; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2175 = mask_2[3] ? byte_515 : _GEN_1859; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2176 = _GEN_4490 == 8'hf ? _GEN_2172 : _GEN_1856; // @[executor.scala 473:84]
  wire [7:0] _GEN_2177 = _GEN_4490 == 8'hf ? _GEN_2173 : _GEN_1857; // @[executor.scala 473:84]
  wire [7:0] _GEN_2178 = _GEN_4490 == 8'hf ? _GEN_2174 : _GEN_1858; // @[executor.scala 473:84]
  wire [7:0] _GEN_2179 = _GEN_4490 == 8'hf ? _GEN_2175 : _GEN_1859; // @[executor.scala 473:84]
  wire [7:0] _GEN_2180 = mask_2[0] ? byte_512 : _GEN_1860; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2181 = mask_2[1] ? byte_513 : _GEN_1861; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2182 = mask_2[2] ? byte_514 : _GEN_1862; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2183 = mask_2[3] ? byte_515 : _GEN_1863; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2184 = _GEN_4490 == 8'h10 ? _GEN_2180 : _GEN_1860; // @[executor.scala 473:84]
  wire [7:0] _GEN_2185 = _GEN_4490 == 8'h10 ? _GEN_2181 : _GEN_1861; // @[executor.scala 473:84]
  wire [7:0] _GEN_2186 = _GEN_4490 == 8'h10 ? _GEN_2182 : _GEN_1862; // @[executor.scala 473:84]
  wire [7:0] _GEN_2187 = _GEN_4490 == 8'h10 ? _GEN_2183 : _GEN_1863; // @[executor.scala 473:84]
  wire [7:0] _GEN_2188 = mask_2[0] ? byte_512 : _GEN_1864; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2189 = mask_2[1] ? byte_513 : _GEN_1865; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2190 = mask_2[2] ? byte_514 : _GEN_1866; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2191 = mask_2[3] ? byte_515 : _GEN_1867; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2192 = _GEN_4490 == 8'h11 ? _GEN_2188 : _GEN_1864; // @[executor.scala 473:84]
  wire [7:0] _GEN_2193 = _GEN_4490 == 8'h11 ? _GEN_2189 : _GEN_1865; // @[executor.scala 473:84]
  wire [7:0] _GEN_2194 = _GEN_4490 == 8'h11 ? _GEN_2190 : _GEN_1866; // @[executor.scala 473:84]
  wire [7:0] _GEN_2195 = _GEN_4490 == 8'h11 ? _GEN_2191 : _GEN_1867; // @[executor.scala 473:84]
  wire [7:0] _GEN_2196 = mask_2[0] ? byte_512 : _GEN_1868; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2197 = mask_2[1] ? byte_513 : _GEN_1869; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2198 = mask_2[2] ? byte_514 : _GEN_1870; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2199 = mask_2[3] ? byte_515 : _GEN_1871; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2200 = _GEN_4490 == 8'h12 ? _GEN_2196 : _GEN_1868; // @[executor.scala 473:84]
  wire [7:0] _GEN_2201 = _GEN_4490 == 8'h12 ? _GEN_2197 : _GEN_1869; // @[executor.scala 473:84]
  wire [7:0] _GEN_2202 = _GEN_4490 == 8'h12 ? _GEN_2198 : _GEN_1870; // @[executor.scala 473:84]
  wire [7:0] _GEN_2203 = _GEN_4490 == 8'h12 ? _GEN_2199 : _GEN_1871; // @[executor.scala 473:84]
  wire [7:0] _GEN_2204 = mask_2[0] ? byte_512 : _GEN_1872; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2205 = mask_2[1] ? byte_513 : _GEN_1873; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2206 = mask_2[2] ? byte_514 : _GEN_1874; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2207 = mask_2[3] ? byte_515 : _GEN_1875; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2208 = _GEN_4490 == 8'h13 ? _GEN_2204 : _GEN_1872; // @[executor.scala 473:84]
  wire [7:0] _GEN_2209 = _GEN_4490 == 8'h13 ? _GEN_2205 : _GEN_1873; // @[executor.scala 473:84]
  wire [7:0] _GEN_2210 = _GEN_4490 == 8'h13 ? _GEN_2206 : _GEN_1874; // @[executor.scala 473:84]
  wire [7:0] _GEN_2211 = _GEN_4490 == 8'h13 ? _GEN_2207 : _GEN_1875; // @[executor.scala 473:84]
  wire [7:0] _GEN_2212 = mask_2[0] ? byte_512 : _GEN_1876; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2213 = mask_2[1] ? byte_513 : _GEN_1877; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2214 = mask_2[2] ? byte_514 : _GEN_1878; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2215 = mask_2[3] ? byte_515 : _GEN_1879; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2216 = _GEN_4490 == 8'h14 ? _GEN_2212 : _GEN_1876; // @[executor.scala 473:84]
  wire [7:0] _GEN_2217 = _GEN_4490 == 8'h14 ? _GEN_2213 : _GEN_1877; // @[executor.scala 473:84]
  wire [7:0] _GEN_2218 = _GEN_4490 == 8'h14 ? _GEN_2214 : _GEN_1878; // @[executor.scala 473:84]
  wire [7:0] _GEN_2219 = _GEN_4490 == 8'h14 ? _GEN_2215 : _GEN_1879; // @[executor.scala 473:84]
  wire [7:0] _GEN_2220 = mask_2[0] ? byte_512 : _GEN_1880; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2221 = mask_2[1] ? byte_513 : _GEN_1881; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2222 = mask_2[2] ? byte_514 : _GEN_1882; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2223 = mask_2[3] ? byte_515 : _GEN_1883; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2224 = _GEN_4490 == 8'h15 ? _GEN_2220 : _GEN_1880; // @[executor.scala 473:84]
  wire [7:0] _GEN_2225 = _GEN_4490 == 8'h15 ? _GEN_2221 : _GEN_1881; // @[executor.scala 473:84]
  wire [7:0] _GEN_2226 = _GEN_4490 == 8'h15 ? _GEN_2222 : _GEN_1882; // @[executor.scala 473:84]
  wire [7:0] _GEN_2227 = _GEN_4490 == 8'h15 ? _GEN_2223 : _GEN_1883; // @[executor.scala 473:84]
  wire [7:0] _GEN_2228 = mask_2[0] ? byte_512 : _GEN_1884; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2229 = mask_2[1] ? byte_513 : _GEN_1885; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2230 = mask_2[2] ? byte_514 : _GEN_1886; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2231 = mask_2[3] ? byte_515 : _GEN_1887; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2232 = _GEN_4490 == 8'h16 ? _GEN_2228 : _GEN_1884; // @[executor.scala 473:84]
  wire [7:0] _GEN_2233 = _GEN_4490 == 8'h16 ? _GEN_2229 : _GEN_1885; // @[executor.scala 473:84]
  wire [7:0] _GEN_2234 = _GEN_4490 == 8'h16 ? _GEN_2230 : _GEN_1886; // @[executor.scala 473:84]
  wire [7:0] _GEN_2235 = _GEN_4490 == 8'h16 ? _GEN_2231 : _GEN_1887; // @[executor.scala 473:84]
  wire [7:0] _GEN_2236 = mask_2[0] ? byte_512 : _GEN_1888; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2237 = mask_2[1] ? byte_513 : _GEN_1889; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2238 = mask_2[2] ? byte_514 : _GEN_1890; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2239 = mask_2[3] ? byte_515 : _GEN_1891; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2240 = _GEN_4490 == 8'h17 ? _GEN_2236 : _GEN_1888; // @[executor.scala 473:84]
  wire [7:0] _GEN_2241 = _GEN_4490 == 8'h17 ? _GEN_2237 : _GEN_1889; // @[executor.scala 473:84]
  wire [7:0] _GEN_2242 = _GEN_4490 == 8'h17 ? _GEN_2238 : _GEN_1890; // @[executor.scala 473:84]
  wire [7:0] _GEN_2243 = _GEN_4490 == 8'h17 ? _GEN_2239 : _GEN_1891; // @[executor.scala 473:84]
  wire [7:0] _GEN_2244 = mask_2[0] ? byte_512 : _GEN_1892; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2245 = mask_2[1] ? byte_513 : _GEN_1893; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2246 = mask_2[2] ? byte_514 : _GEN_1894; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2247 = mask_2[3] ? byte_515 : _GEN_1895; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2248 = _GEN_4490 == 8'h18 ? _GEN_2244 : _GEN_1892; // @[executor.scala 473:84]
  wire [7:0] _GEN_2249 = _GEN_4490 == 8'h18 ? _GEN_2245 : _GEN_1893; // @[executor.scala 473:84]
  wire [7:0] _GEN_2250 = _GEN_4490 == 8'h18 ? _GEN_2246 : _GEN_1894; // @[executor.scala 473:84]
  wire [7:0] _GEN_2251 = _GEN_4490 == 8'h18 ? _GEN_2247 : _GEN_1895; // @[executor.scala 473:84]
  wire [7:0] _GEN_2252 = mask_2[0] ? byte_512 : _GEN_1896; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2253 = mask_2[1] ? byte_513 : _GEN_1897; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2254 = mask_2[2] ? byte_514 : _GEN_1898; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2255 = mask_2[3] ? byte_515 : _GEN_1899; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2256 = _GEN_4490 == 8'h19 ? _GEN_2252 : _GEN_1896; // @[executor.scala 473:84]
  wire [7:0] _GEN_2257 = _GEN_4490 == 8'h19 ? _GEN_2253 : _GEN_1897; // @[executor.scala 473:84]
  wire [7:0] _GEN_2258 = _GEN_4490 == 8'h19 ? _GEN_2254 : _GEN_1898; // @[executor.scala 473:84]
  wire [7:0] _GEN_2259 = _GEN_4490 == 8'h19 ? _GEN_2255 : _GEN_1899; // @[executor.scala 473:84]
  wire [7:0] _GEN_2260 = mask_2[0] ? byte_512 : _GEN_1900; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2261 = mask_2[1] ? byte_513 : _GEN_1901; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2262 = mask_2[2] ? byte_514 : _GEN_1902; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2263 = mask_2[3] ? byte_515 : _GEN_1903; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2264 = _GEN_4490 == 8'h1a ? _GEN_2260 : _GEN_1900; // @[executor.scala 473:84]
  wire [7:0] _GEN_2265 = _GEN_4490 == 8'h1a ? _GEN_2261 : _GEN_1901; // @[executor.scala 473:84]
  wire [7:0] _GEN_2266 = _GEN_4490 == 8'h1a ? _GEN_2262 : _GEN_1902; // @[executor.scala 473:84]
  wire [7:0] _GEN_2267 = _GEN_4490 == 8'h1a ? _GEN_2263 : _GEN_1903; // @[executor.scala 473:84]
  wire [7:0] _GEN_2268 = mask_2[0] ? byte_512 : _GEN_1904; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2269 = mask_2[1] ? byte_513 : _GEN_1905; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2270 = mask_2[2] ? byte_514 : _GEN_1906; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2271 = mask_2[3] ? byte_515 : _GEN_1907; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2272 = _GEN_4490 == 8'h1b ? _GEN_2268 : _GEN_1904; // @[executor.scala 473:84]
  wire [7:0] _GEN_2273 = _GEN_4490 == 8'h1b ? _GEN_2269 : _GEN_1905; // @[executor.scala 473:84]
  wire [7:0] _GEN_2274 = _GEN_4490 == 8'h1b ? _GEN_2270 : _GEN_1906; // @[executor.scala 473:84]
  wire [7:0] _GEN_2275 = _GEN_4490 == 8'h1b ? _GEN_2271 : _GEN_1907; // @[executor.scala 473:84]
  wire [7:0] _GEN_2276 = mask_2[0] ? byte_512 : _GEN_1908; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2277 = mask_2[1] ? byte_513 : _GEN_1909; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2278 = mask_2[2] ? byte_514 : _GEN_1910; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2279 = mask_2[3] ? byte_515 : _GEN_1911; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2280 = _GEN_4490 == 8'h1c ? _GEN_2276 : _GEN_1908; // @[executor.scala 473:84]
  wire [7:0] _GEN_2281 = _GEN_4490 == 8'h1c ? _GEN_2277 : _GEN_1909; // @[executor.scala 473:84]
  wire [7:0] _GEN_2282 = _GEN_4490 == 8'h1c ? _GEN_2278 : _GEN_1910; // @[executor.scala 473:84]
  wire [7:0] _GEN_2283 = _GEN_4490 == 8'h1c ? _GEN_2279 : _GEN_1911; // @[executor.scala 473:84]
  wire [7:0] _GEN_2284 = mask_2[0] ? byte_512 : _GEN_1912; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2285 = mask_2[1] ? byte_513 : _GEN_1913; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2286 = mask_2[2] ? byte_514 : _GEN_1914; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2287 = mask_2[3] ? byte_515 : _GEN_1915; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2288 = _GEN_4490 == 8'h1d ? _GEN_2284 : _GEN_1912; // @[executor.scala 473:84]
  wire [7:0] _GEN_2289 = _GEN_4490 == 8'h1d ? _GEN_2285 : _GEN_1913; // @[executor.scala 473:84]
  wire [7:0] _GEN_2290 = _GEN_4490 == 8'h1d ? _GEN_2286 : _GEN_1914; // @[executor.scala 473:84]
  wire [7:0] _GEN_2291 = _GEN_4490 == 8'h1d ? _GEN_2287 : _GEN_1915; // @[executor.scala 473:84]
  wire [7:0] _GEN_2292 = mask_2[0] ? byte_512 : _GEN_1916; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2293 = mask_2[1] ? byte_513 : _GEN_1917; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2294 = mask_2[2] ? byte_514 : _GEN_1918; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2295 = mask_2[3] ? byte_515 : _GEN_1919; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2296 = _GEN_4490 == 8'h1e ? _GEN_2292 : _GEN_1916; // @[executor.scala 473:84]
  wire [7:0] _GEN_2297 = _GEN_4490 == 8'h1e ? _GEN_2293 : _GEN_1917; // @[executor.scala 473:84]
  wire [7:0] _GEN_2298 = _GEN_4490 == 8'h1e ? _GEN_2294 : _GEN_1918; // @[executor.scala 473:84]
  wire [7:0] _GEN_2299 = _GEN_4490 == 8'h1e ? _GEN_2295 : _GEN_1919; // @[executor.scala 473:84]
  wire [7:0] _GEN_2300 = mask_2[0] ? byte_512 : _GEN_1920; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2301 = mask_2[1] ? byte_513 : _GEN_1921; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2302 = mask_2[2] ? byte_514 : _GEN_1922; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2303 = mask_2[3] ? byte_515 : _GEN_1923; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2304 = _GEN_4490 == 8'h1f ? _GEN_2300 : _GEN_1920; // @[executor.scala 473:84]
  wire [7:0] _GEN_2305 = _GEN_4490 == 8'h1f ? _GEN_2301 : _GEN_1921; // @[executor.scala 473:84]
  wire [7:0] _GEN_2306 = _GEN_4490 == 8'h1f ? _GEN_2302 : _GEN_1922; // @[executor.scala 473:84]
  wire [7:0] _GEN_2307 = _GEN_4490 == 8'h1f ? _GEN_2303 : _GEN_1923; // @[executor.scala 473:84]
  wire [7:0] _GEN_2308 = mask_2[0] ? byte_512 : _GEN_1924; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2309 = mask_2[1] ? byte_513 : _GEN_1925; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2310 = mask_2[2] ? byte_514 : _GEN_1926; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2311 = mask_2[3] ? byte_515 : _GEN_1927; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2312 = _GEN_4490 == 8'h20 ? _GEN_2308 : _GEN_1924; // @[executor.scala 473:84]
  wire [7:0] _GEN_2313 = _GEN_4490 == 8'h20 ? _GEN_2309 : _GEN_1925; // @[executor.scala 473:84]
  wire [7:0] _GEN_2314 = _GEN_4490 == 8'h20 ? _GEN_2310 : _GEN_1926; // @[executor.scala 473:84]
  wire [7:0] _GEN_2315 = _GEN_4490 == 8'h20 ? _GEN_2311 : _GEN_1927; // @[executor.scala 473:84]
  wire [7:0] _GEN_2316 = mask_2[0] ? byte_512 : _GEN_1928; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2317 = mask_2[1] ? byte_513 : _GEN_1929; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2318 = mask_2[2] ? byte_514 : _GEN_1930; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2319 = mask_2[3] ? byte_515 : _GEN_1931; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2320 = _GEN_4490 == 8'h21 ? _GEN_2316 : _GEN_1928; // @[executor.scala 473:84]
  wire [7:0] _GEN_2321 = _GEN_4490 == 8'h21 ? _GEN_2317 : _GEN_1929; // @[executor.scala 473:84]
  wire [7:0] _GEN_2322 = _GEN_4490 == 8'h21 ? _GEN_2318 : _GEN_1930; // @[executor.scala 473:84]
  wire [7:0] _GEN_2323 = _GEN_4490 == 8'h21 ? _GEN_2319 : _GEN_1931; // @[executor.scala 473:84]
  wire [7:0] _GEN_2324 = mask_2[0] ? byte_512 : _GEN_1932; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2325 = mask_2[1] ? byte_513 : _GEN_1933; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2326 = mask_2[2] ? byte_514 : _GEN_1934; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2327 = mask_2[3] ? byte_515 : _GEN_1935; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2328 = _GEN_4490 == 8'h22 ? _GEN_2324 : _GEN_1932; // @[executor.scala 473:84]
  wire [7:0] _GEN_2329 = _GEN_4490 == 8'h22 ? _GEN_2325 : _GEN_1933; // @[executor.scala 473:84]
  wire [7:0] _GEN_2330 = _GEN_4490 == 8'h22 ? _GEN_2326 : _GEN_1934; // @[executor.scala 473:84]
  wire [7:0] _GEN_2331 = _GEN_4490 == 8'h22 ? _GEN_2327 : _GEN_1935; // @[executor.scala 473:84]
  wire [7:0] _GEN_2332 = mask_2[0] ? byte_512 : _GEN_1936; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2333 = mask_2[1] ? byte_513 : _GEN_1937; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2334 = mask_2[2] ? byte_514 : _GEN_1938; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2335 = mask_2[3] ? byte_515 : _GEN_1939; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2336 = _GEN_4490 == 8'h23 ? _GEN_2332 : _GEN_1936; // @[executor.scala 473:84]
  wire [7:0] _GEN_2337 = _GEN_4490 == 8'h23 ? _GEN_2333 : _GEN_1937; // @[executor.scala 473:84]
  wire [7:0] _GEN_2338 = _GEN_4490 == 8'h23 ? _GEN_2334 : _GEN_1938; // @[executor.scala 473:84]
  wire [7:0] _GEN_2339 = _GEN_4490 == 8'h23 ? _GEN_2335 : _GEN_1939; // @[executor.scala 473:84]
  wire [7:0] _GEN_2340 = mask_2[0] ? byte_512 : _GEN_1940; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2341 = mask_2[1] ? byte_513 : _GEN_1941; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2342 = mask_2[2] ? byte_514 : _GEN_1942; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2343 = mask_2[3] ? byte_515 : _GEN_1943; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2344 = _GEN_4490 == 8'h24 ? _GEN_2340 : _GEN_1940; // @[executor.scala 473:84]
  wire [7:0] _GEN_2345 = _GEN_4490 == 8'h24 ? _GEN_2341 : _GEN_1941; // @[executor.scala 473:84]
  wire [7:0] _GEN_2346 = _GEN_4490 == 8'h24 ? _GEN_2342 : _GEN_1942; // @[executor.scala 473:84]
  wire [7:0] _GEN_2347 = _GEN_4490 == 8'h24 ? _GEN_2343 : _GEN_1943; // @[executor.scala 473:84]
  wire [7:0] _GEN_2348 = mask_2[0] ? byte_512 : _GEN_1944; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2349 = mask_2[1] ? byte_513 : _GEN_1945; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2350 = mask_2[2] ? byte_514 : _GEN_1946; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2351 = mask_2[3] ? byte_515 : _GEN_1947; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2352 = _GEN_4490 == 8'h25 ? _GEN_2348 : _GEN_1944; // @[executor.scala 473:84]
  wire [7:0] _GEN_2353 = _GEN_4490 == 8'h25 ? _GEN_2349 : _GEN_1945; // @[executor.scala 473:84]
  wire [7:0] _GEN_2354 = _GEN_4490 == 8'h25 ? _GEN_2350 : _GEN_1946; // @[executor.scala 473:84]
  wire [7:0] _GEN_2355 = _GEN_4490 == 8'h25 ? _GEN_2351 : _GEN_1947; // @[executor.scala 473:84]
  wire [7:0] _GEN_2356 = mask_2[0] ? byte_512 : _GEN_1948; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2357 = mask_2[1] ? byte_513 : _GEN_1949; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2358 = mask_2[2] ? byte_514 : _GEN_1950; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2359 = mask_2[3] ? byte_515 : _GEN_1951; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2360 = _GEN_4490 == 8'h26 ? _GEN_2356 : _GEN_1948; // @[executor.scala 473:84]
  wire [7:0] _GEN_2361 = _GEN_4490 == 8'h26 ? _GEN_2357 : _GEN_1949; // @[executor.scala 473:84]
  wire [7:0] _GEN_2362 = _GEN_4490 == 8'h26 ? _GEN_2358 : _GEN_1950; // @[executor.scala 473:84]
  wire [7:0] _GEN_2363 = _GEN_4490 == 8'h26 ? _GEN_2359 : _GEN_1951; // @[executor.scala 473:84]
  wire [7:0] _GEN_2364 = mask_2[0] ? byte_512 : _GEN_1952; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2365 = mask_2[1] ? byte_513 : _GEN_1953; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2366 = mask_2[2] ? byte_514 : _GEN_1954; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2367 = mask_2[3] ? byte_515 : _GEN_1955; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2368 = _GEN_4490 == 8'h27 ? _GEN_2364 : _GEN_1952; // @[executor.scala 473:84]
  wire [7:0] _GEN_2369 = _GEN_4490 == 8'h27 ? _GEN_2365 : _GEN_1953; // @[executor.scala 473:84]
  wire [7:0] _GEN_2370 = _GEN_4490 == 8'h27 ? _GEN_2366 : _GEN_1954; // @[executor.scala 473:84]
  wire [7:0] _GEN_2371 = _GEN_4490 == 8'h27 ? _GEN_2367 : _GEN_1955; // @[executor.scala 473:84]
  wire [7:0] _GEN_2372 = mask_2[0] ? byte_512 : _GEN_1956; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2373 = mask_2[1] ? byte_513 : _GEN_1957; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2374 = mask_2[2] ? byte_514 : _GEN_1958; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2375 = mask_2[3] ? byte_515 : _GEN_1959; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2376 = _GEN_4490 == 8'h28 ? _GEN_2372 : _GEN_1956; // @[executor.scala 473:84]
  wire [7:0] _GEN_2377 = _GEN_4490 == 8'h28 ? _GEN_2373 : _GEN_1957; // @[executor.scala 473:84]
  wire [7:0] _GEN_2378 = _GEN_4490 == 8'h28 ? _GEN_2374 : _GEN_1958; // @[executor.scala 473:84]
  wire [7:0] _GEN_2379 = _GEN_4490 == 8'h28 ? _GEN_2375 : _GEN_1959; // @[executor.scala 473:84]
  wire [7:0] _GEN_2380 = mask_2[0] ? byte_512 : _GEN_1960; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2381 = mask_2[1] ? byte_513 : _GEN_1961; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2382 = mask_2[2] ? byte_514 : _GEN_1962; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2383 = mask_2[3] ? byte_515 : _GEN_1963; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2384 = _GEN_4490 == 8'h29 ? _GEN_2380 : _GEN_1960; // @[executor.scala 473:84]
  wire [7:0] _GEN_2385 = _GEN_4490 == 8'h29 ? _GEN_2381 : _GEN_1961; // @[executor.scala 473:84]
  wire [7:0] _GEN_2386 = _GEN_4490 == 8'h29 ? _GEN_2382 : _GEN_1962; // @[executor.scala 473:84]
  wire [7:0] _GEN_2387 = _GEN_4490 == 8'h29 ? _GEN_2383 : _GEN_1963; // @[executor.scala 473:84]
  wire [7:0] _GEN_2388 = mask_2[0] ? byte_512 : _GEN_1964; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2389 = mask_2[1] ? byte_513 : _GEN_1965; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2390 = mask_2[2] ? byte_514 : _GEN_1966; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2391 = mask_2[3] ? byte_515 : _GEN_1967; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2392 = _GEN_4490 == 8'h2a ? _GEN_2388 : _GEN_1964; // @[executor.scala 473:84]
  wire [7:0] _GEN_2393 = _GEN_4490 == 8'h2a ? _GEN_2389 : _GEN_1965; // @[executor.scala 473:84]
  wire [7:0] _GEN_2394 = _GEN_4490 == 8'h2a ? _GEN_2390 : _GEN_1966; // @[executor.scala 473:84]
  wire [7:0] _GEN_2395 = _GEN_4490 == 8'h2a ? _GEN_2391 : _GEN_1967; // @[executor.scala 473:84]
  wire [7:0] _GEN_2396 = mask_2[0] ? byte_512 : _GEN_1968; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2397 = mask_2[1] ? byte_513 : _GEN_1969; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2398 = mask_2[2] ? byte_514 : _GEN_1970; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2399 = mask_2[3] ? byte_515 : _GEN_1971; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2400 = _GEN_4490 == 8'h2b ? _GEN_2396 : _GEN_1968; // @[executor.scala 473:84]
  wire [7:0] _GEN_2401 = _GEN_4490 == 8'h2b ? _GEN_2397 : _GEN_1969; // @[executor.scala 473:84]
  wire [7:0] _GEN_2402 = _GEN_4490 == 8'h2b ? _GEN_2398 : _GEN_1970; // @[executor.scala 473:84]
  wire [7:0] _GEN_2403 = _GEN_4490 == 8'h2b ? _GEN_2399 : _GEN_1971; // @[executor.scala 473:84]
  wire [7:0] _GEN_2404 = mask_2[0] ? byte_512 : _GEN_1972; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2405 = mask_2[1] ? byte_513 : _GEN_1973; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2406 = mask_2[2] ? byte_514 : _GEN_1974; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2407 = mask_2[3] ? byte_515 : _GEN_1975; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2408 = _GEN_4490 == 8'h2c ? _GEN_2404 : _GEN_1972; // @[executor.scala 473:84]
  wire [7:0] _GEN_2409 = _GEN_4490 == 8'h2c ? _GEN_2405 : _GEN_1973; // @[executor.scala 473:84]
  wire [7:0] _GEN_2410 = _GEN_4490 == 8'h2c ? _GEN_2406 : _GEN_1974; // @[executor.scala 473:84]
  wire [7:0] _GEN_2411 = _GEN_4490 == 8'h2c ? _GEN_2407 : _GEN_1975; // @[executor.scala 473:84]
  wire [7:0] _GEN_2412 = mask_2[0] ? byte_512 : _GEN_1976; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2413 = mask_2[1] ? byte_513 : _GEN_1977; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2414 = mask_2[2] ? byte_514 : _GEN_1978; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2415 = mask_2[3] ? byte_515 : _GEN_1979; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2416 = _GEN_4490 == 8'h2d ? _GEN_2412 : _GEN_1976; // @[executor.scala 473:84]
  wire [7:0] _GEN_2417 = _GEN_4490 == 8'h2d ? _GEN_2413 : _GEN_1977; // @[executor.scala 473:84]
  wire [7:0] _GEN_2418 = _GEN_4490 == 8'h2d ? _GEN_2414 : _GEN_1978; // @[executor.scala 473:84]
  wire [7:0] _GEN_2419 = _GEN_4490 == 8'h2d ? _GEN_2415 : _GEN_1979; // @[executor.scala 473:84]
  wire [7:0] _GEN_2420 = mask_2[0] ? byte_512 : _GEN_1980; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2421 = mask_2[1] ? byte_513 : _GEN_1981; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2422 = mask_2[2] ? byte_514 : _GEN_1982; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2423 = mask_2[3] ? byte_515 : _GEN_1983; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2424 = _GEN_4490 == 8'h2e ? _GEN_2420 : _GEN_1980; // @[executor.scala 473:84]
  wire [7:0] _GEN_2425 = _GEN_4490 == 8'h2e ? _GEN_2421 : _GEN_1981; // @[executor.scala 473:84]
  wire [7:0] _GEN_2426 = _GEN_4490 == 8'h2e ? _GEN_2422 : _GEN_1982; // @[executor.scala 473:84]
  wire [7:0] _GEN_2427 = _GEN_4490 == 8'h2e ? _GEN_2423 : _GEN_1983; // @[executor.scala 473:84]
  wire [7:0] _GEN_2428 = mask_2[0] ? byte_512 : _GEN_1984; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2429 = mask_2[1] ? byte_513 : _GEN_1985; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2430 = mask_2[2] ? byte_514 : _GEN_1986; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2431 = mask_2[3] ? byte_515 : _GEN_1987; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2432 = _GEN_4490 == 8'h2f ? _GEN_2428 : _GEN_1984; // @[executor.scala 473:84]
  wire [7:0] _GEN_2433 = _GEN_4490 == 8'h2f ? _GEN_2429 : _GEN_1985; // @[executor.scala 473:84]
  wire [7:0] _GEN_2434 = _GEN_4490 == 8'h2f ? _GEN_2430 : _GEN_1986; // @[executor.scala 473:84]
  wire [7:0] _GEN_2435 = _GEN_4490 == 8'h2f ? _GEN_2431 : _GEN_1987; // @[executor.scala 473:84]
  wire [7:0] _GEN_2436 = mask_2[0] ? byte_512 : _GEN_1988; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2437 = mask_2[1] ? byte_513 : _GEN_1989; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2438 = mask_2[2] ? byte_514 : _GEN_1990; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2439 = mask_2[3] ? byte_515 : _GEN_1991; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2440 = _GEN_4490 == 8'h30 ? _GEN_2436 : _GEN_1988; // @[executor.scala 473:84]
  wire [7:0] _GEN_2441 = _GEN_4490 == 8'h30 ? _GEN_2437 : _GEN_1989; // @[executor.scala 473:84]
  wire [7:0] _GEN_2442 = _GEN_4490 == 8'h30 ? _GEN_2438 : _GEN_1990; // @[executor.scala 473:84]
  wire [7:0] _GEN_2443 = _GEN_4490 == 8'h30 ? _GEN_2439 : _GEN_1991; // @[executor.scala 473:84]
  wire [7:0] _GEN_2444 = mask_2[0] ? byte_512 : _GEN_1992; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2445 = mask_2[1] ? byte_513 : _GEN_1993; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2446 = mask_2[2] ? byte_514 : _GEN_1994; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2447 = mask_2[3] ? byte_515 : _GEN_1995; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2448 = _GEN_4490 == 8'h31 ? _GEN_2444 : _GEN_1992; // @[executor.scala 473:84]
  wire [7:0] _GEN_2449 = _GEN_4490 == 8'h31 ? _GEN_2445 : _GEN_1993; // @[executor.scala 473:84]
  wire [7:0] _GEN_2450 = _GEN_4490 == 8'h31 ? _GEN_2446 : _GEN_1994; // @[executor.scala 473:84]
  wire [7:0] _GEN_2451 = _GEN_4490 == 8'h31 ? _GEN_2447 : _GEN_1995; // @[executor.scala 473:84]
  wire [7:0] _GEN_2452 = mask_2[0] ? byte_512 : _GEN_1996; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2453 = mask_2[1] ? byte_513 : _GEN_1997; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2454 = mask_2[2] ? byte_514 : _GEN_1998; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2455 = mask_2[3] ? byte_515 : _GEN_1999; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2456 = _GEN_4490 == 8'h32 ? _GEN_2452 : _GEN_1996; // @[executor.scala 473:84]
  wire [7:0] _GEN_2457 = _GEN_4490 == 8'h32 ? _GEN_2453 : _GEN_1997; // @[executor.scala 473:84]
  wire [7:0] _GEN_2458 = _GEN_4490 == 8'h32 ? _GEN_2454 : _GEN_1998; // @[executor.scala 473:84]
  wire [7:0] _GEN_2459 = _GEN_4490 == 8'h32 ? _GEN_2455 : _GEN_1999; // @[executor.scala 473:84]
  wire [7:0] _GEN_2460 = mask_2[0] ? byte_512 : _GEN_2000; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2461 = mask_2[1] ? byte_513 : _GEN_2001; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2462 = mask_2[2] ? byte_514 : _GEN_2002; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2463 = mask_2[3] ? byte_515 : _GEN_2003; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2464 = _GEN_4490 == 8'h33 ? _GEN_2460 : _GEN_2000; // @[executor.scala 473:84]
  wire [7:0] _GEN_2465 = _GEN_4490 == 8'h33 ? _GEN_2461 : _GEN_2001; // @[executor.scala 473:84]
  wire [7:0] _GEN_2466 = _GEN_4490 == 8'h33 ? _GEN_2462 : _GEN_2002; // @[executor.scala 473:84]
  wire [7:0] _GEN_2467 = _GEN_4490 == 8'h33 ? _GEN_2463 : _GEN_2003; // @[executor.scala 473:84]
  wire [7:0] _GEN_2468 = mask_2[0] ? byte_512 : _GEN_2004; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2469 = mask_2[1] ? byte_513 : _GEN_2005; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2470 = mask_2[2] ? byte_514 : _GEN_2006; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2471 = mask_2[3] ? byte_515 : _GEN_2007; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2472 = _GEN_4490 == 8'h34 ? _GEN_2468 : _GEN_2004; // @[executor.scala 473:84]
  wire [7:0] _GEN_2473 = _GEN_4490 == 8'h34 ? _GEN_2469 : _GEN_2005; // @[executor.scala 473:84]
  wire [7:0] _GEN_2474 = _GEN_4490 == 8'h34 ? _GEN_2470 : _GEN_2006; // @[executor.scala 473:84]
  wire [7:0] _GEN_2475 = _GEN_4490 == 8'h34 ? _GEN_2471 : _GEN_2007; // @[executor.scala 473:84]
  wire [7:0] _GEN_2476 = mask_2[0] ? byte_512 : _GEN_2008; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2477 = mask_2[1] ? byte_513 : _GEN_2009; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2478 = mask_2[2] ? byte_514 : _GEN_2010; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2479 = mask_2[3] ? byte_515 : _GEN_2011; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2480 = _GEN_4490 == 8'h35 ? _GEN_2476 : _GEN_2008; // @[executor.scala 473:84]
  wire [7:0] _GEN_2481 = _GEN_4490 == 8'h35 ? _GEN_2477 : _GEN_2009; // @[executor.scala 473:84]
  wire [7:0] _GEN_2482 = _GEN_4490 == 8'h35 ? _GEN_2478 : _GEN_2010; // @[executor.scala 473:84]
  wire [7:0] _GEN_2483 = _GEN_4490 == 8'h35 ? _GEN_2479 : _GEN_2011; // @[executor.scala 473:84]
  wire [7:0] _GEN_2484 = mask_2[0] ? byte_512 : _GEN_2012; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2485 = mask_2[1] ? byte_513 : _GEN_2013; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2486 = mask_2[2] ? byte_514 : _GEN_2014; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2487 = mask_2[3] ? byte_515 : _GEN_2015; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2488 = _GEN_4490 == 8'h36 ? _GEN_2484 : _GEN_2012; // @[executor.scala 473:84]
  wire [7:0] _GEN_2489 = _GEN_4490 == 8'h36 ? _GEN_2485 : _GEN_2013; // @[executor.scala 473:84]
  wire [7:0] _GEN_2490 = _GEN_4490 == 8'h36 ? _GEN_2486 : _GEN_2014; // @[executor.scala 473:84]
  wire [7:0] _GEN_2491 = _GEN_4490 == 8'h36 ? _GEN_2487 : _GEN_2015; // @[executor.scala 473:84]
  wire [7:0] _GEN_2492 = mask_2[0] ? byte_512 : _GEN_2016; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2493 = mask_2[1] ? byte_513 : _GEN_2017; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2494 = mask_2[2] ? byte_514 : _GEN_2018; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2495 = mask_2[3] ? byte_515 : _GEN_2019; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2496 = _GEN_4490 == 8'h37 ? _GEN_2492 : _GEN_2016; // @[executor.scala 473:84]
  wire [7:0] _GEN_2497 = _GEN_4490 == 8'h37 ? _GEN_2493 : _GEN_2017; // @[executor.scala 473:84]
  wire [7:0] _GEN_2498 = _GEN_4490 == 8'h37 ? _GEN_2494 : _GEN_2018; // @[executor.scala 473:84]
  wire [7:0] _GEN_2499 = _GEN_4490 == 8'h37 ? _GEN_2495 : _GEN_2019; // @[executor.scala 473:84]
  wire [7:0] _GEN_2500 = mask_2[0] ? byte_512 : _GEN_2020; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2501 = mask_2[1] ? byte_513 : _GEN_2021; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2502 = mask_2[2] ? byte_514 : _GEN_2022; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2503 = mask_2[3] ? byte_515 : _GEN_2023; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2504 = _GEN_4490 == 8'h38 ? _GEN_2500 : _GEN_2020; // @[executor.scala 473:84]
  wire [7:0] _GEN_2505 = _GEN_4490 == 8'h38 ? _GEN_2501 : _GEN_2021; // @[executor.scala 473:84]
  wire [7:0] _GEN_2506 = _GEN_4490 == 8'h38 ? _GEN_2502 : _GEN_2022; // @[executor.scala 473:84]
  wire [7:0] _GEN_2507 = _GEN_4490 == 8'h38 ? _GEN_2503 : _GEN_2023; // @[executor.scala 473:84]
  wire [7:0] _GEN_2508 = mask_2[0] ? byte_512 : _GEN_2024; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2509 = mask_2[1] ? byte_513 : _GEN_2025; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2510 = mask_2[2] ? byte_514 : _GEN_2026; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2511 = mask_2[3] ? byte_515 : _GEN_2027; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2512 = _GEN_4490 == 8'h39 ? _GEN_2508 : _GEN_2024; // @[executor.scala 473:84]
  wire [7:0] _GEN_2513 = _GEN_4490 == 8'h39 ? _GEN_2509 : _GEN_2025; // @[executor.scala 473:84]
  wire [7:0] _GEN_2514 = _GEN_4490 == 8'h39 ? _GEN_2510 : _GEN_2026; // @[executor.scala 473:84]
  wire [7:0] _GEN_2515 = _GEN_4490 == 8'h39 ? _GEN_2511 : _GEN_2027; // @[executor.scala 473:84]
  wire [7:0] _GEN_2516 = mask_2[0] ? byte_512 : _GEN_2028; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2517 = mask_2[1] ? byte_513 : _GEN_2029; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2518 = mask_2[2] ? byte_514 : _GEN_2030; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2519 = mask_2[3] ? byte_515 : _GEN_2031; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2520 = _GEN_4490 == 8'h3a ? _GEN_2516 : _GEN_2028; // @[executor.scala 473:84]
  wire [7:0] _GEN_2521 = _GEN_4490 == 8'h3a ? _GEN_2517 : _GEN_2029; // @[executor.scala 473:84]
  wire [7:0] _GEN_2522 = _GEN_4490 == 8'h3a ? _GEN_2518 : _GEN_2030; // @[executor.scala 473:84]
  wire [7:0] _GEN_2523 = _GEN_4490 == 8'h3a ? _GEN_2519 : _GEN_2031; // @[executor.scala 473:84]
  wire [7:0] _GEN_2524 = mask_2[0] ? byte_512 : _GEN_2032; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2525 = mask_2[1] ? byte_513 : _GEN_2033; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2526 = mask_2[2] ? byte_514 : _GEN_2034; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2527 = mask_2[3] ? byte_515 : _GEN_2035; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2528 = _GEN_4490 == 8'h3b ? _GEN_2524 : _GEN_2032; // @[executor.scala 473:84]
  wire [7:0] _GEN_2529 = _GEN_4490 == 8'h3b ? _GEN_2525 : _GEN_2033; // @[executor.scala 473:84]
  wire [7:0] _GEN_2530 = _GEN_4490 == 8'h3b ? _GEN_2526 : _GEN_2034; // @[executor.scala 473:84]
  wire [7:0] _GEN_2531 = _GEN_4490 == 8'h3b ? _GEN_2527 : _GEN_2035; // @[executor.scala 473:84]
  wire [7:0] _GEN_2532 = mask_2[0] ? byte_512 : _GEN_2036; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2533 = mask_2[1] ? byte_513 : _GEN_2037; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2534 = mask_2[2] ? byte_514 : _GEN_2038; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2535 = mask_2[3] ? byte_515 : _GEN_2039; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2536 = _GEN_4490 == 8'h3c ? _GEN_2532 : _GEN_2036; // @[executor.scala 473:84]
  wire [7:0] _GEN_2537 = _GEN_4490 == 8'h3c ? _GEN_2533 : _GEN_2037; // @[executor.scala 473:84]
  wire [7:0] _GEN_2538 = _GEN_4490 == 8'h3c ? _GEN_2534 : _GEN_2038; // @[executor.scala 473:84]
  wire [7:0] _GEN_2539 = _GEN_4490 == 8'h3c ? _GEN_2535 : _GEN_2039; // @[executor.scala 473:84]
  wire [7:0] _GEN_2540 = mask_2[0] ? byte_512 : _GEN_2040; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2541 = mask_2[1] ? byte_513 : _GEN_2041; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2542 = mask_2[2] ? byte_514 : _GEN_2042; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2543 = mask_2[3] ? byte_515 : _GEN_2043; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2544 = _GEN_4490 == 8'h3d ? _GEN_2540 : _GEN_2040; // @[executor.scala 473:84]
  wire [7:0] _GEN_2545 = _GEN_4490 == 8'h3d ? _GEN_2541 : _GEN_2041; // @[executor.scala 473:84]
  wire [7:0] _GEN_2546 = _GEN_4490 == 8'h3d ? _GEN_2542 : _GEN_2042; // @[executor.scala 473:84]
  wire [7:0] _GEN_2547 = _GEN_4490 == 8'h3d ? _GEN_2543 : _GEN_2043; // @[executor.scala 473:84]
  wire [7:0] _GEN_2548 = mask_2[0] ? byte_512 : _GEN_2044; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2549 = mask_2[1] ? byte_513 : _GEN_2045; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2550 = mask_2[2] ? byte_514 : _GEN_2046; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2551 = mask_2[3] ? byte_515 : _GEN_2047; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2552 = _GEN_4490 == 8'h3e ? _GEN_2548 : _GEN_2044; // @[executor.scala 473:84]
  wire [7:0] _GEN_2553 = _GEN_4490 == 8'h3e ? _GEN_2549 : _GEN_2045; // @[executor.scala 473:84]
  wire [7:0] _GEN_2554 = _GEN_4490 == 8'h3e ? _GEN_2550 : _GEN_2046; // @[executor.scala 473:84]
  wire [7:0] _GEN_2555 = _GEN_4490 == 8'h3e ? _GEN_2551 : _GEN_2047; // @[executor.scala 473:84]
  wire [7:0] _GEN_2556 = mask_2[0] ? byte_512 : _GEN_2048; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2557 = mask_2[1] ? byte_513 : _GEN_2049; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2558 = mask_2[2] ? byte_514 : _GEN_2050; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2559 = mask_2[3] ? byte_515 : _GEN_2051; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2560 = _GEN_4490 == 8'h3f ? _GEN_2556 : _GEN_2048; // @[executor.scala 473:84]
  wire [7:0] _GEN_2561 = _GEN_4490 == 8'h3f ? _GEN_2557 : _GEN_2049; // @[executor.scala 473:84]
  wire [7:0] _GEN_2562 = _GEN_4490 == 8'h3f ? _GEN_2558 : _GEN_2050; // @[executor.scala 473:84]
  wire [7:0] _GEN_2563 = _GEN_4490 == 8'h3f ? _GEN_2559 : _GEN_2051; // @[executor.scala 473:84]
  wire [7:0] _GEN_2564 = opcode_2 != 4'h0 ? _GEN_2056 : _GEN_1796; // @[executor.scala 470:55]
  wire [7:0] _GEN_2565 = opcode_2 != 4'h0 ? _GEN_2057 : _GEN_1797; // @[executor.scala 470:55]
  wire [7:0] _GEN_2566 = opcode_2 != 4'h0 ? _GEN_2058 : _GEN_1798; // @[executor.scala 470:55]
  wire [7:0] _GEN_2567 = opcode_2 != 4'h0 ? _GEN_2059 : _GEN_1799; // @[executor.scala 470:55]
  wire [7:0] _GEN_2568 = opcode_2 != 4'h0 ? _GEN_2064 : _GEN_1800; // @[executor.scala 470:55]
  wire [7:0] _GEN_2569 = opcode_2 != 4'h0 ? _GEN_2065 : _GEN_1801; // @[executor.scala 470:55]
  wire [7:0] _GEN_2570 = opcode_2 != 4'h0 ? _GEN_2066 : _GEN_1802; // @[executor.scala 470:55]
  wire [7:0] _GEN_2571 = opcode_2 != 4'h0 ? _GEN_2067 : _GEN_1803; // @[executor.scala 470:55]
  wire [7:0] _GEN_2572 = opcode_2 != 4'h0 ? _GEN_2072 : _GEN_1804; // @[executor.scala 470:55]
  wire [7:0] _GEN_2573 = opcode_2 != 4'h0 ? _GEN_2073 : _GEN_1805; // @[executor.scala 470:55]
  wire [7:0] _GEN_2574 = opcode_2 != 4'h0 ? _GEN_2074 : _GEN_1806; // @[executor.scala 470:55]
  wire [7:0] _GEN_2575 = opcode_2 != 4'h0 ? _GEN_2075 : _GEN_1807; // @[executor.scala 470:55]
  wire [7:0] _GEN_2576 = opcode_2 != 4'h0 ? _GEN_2080 : _GEN_1808; // @[executor.scala 470:55]
  wire [7:0] _GEN_2577 = opcode_2 != 4'h0 ? _GEN_2081 : _GEN_1809; // @[executor.scala 470:55]
  wire [7:0] _GEN_2578 = opcode_2 != 4'h0 ? _GEN_2082 : _GEN_1810; // @[executor.scala 470:55]
  wire [7:0] _GEN_2579 = opcode_2 != 4'h0 ? _GEN_2083 : _GEN_1811; // @[executor.scala 470:55]
  wire [7:0] _GEN_2580 = opcode_2 != 4'h0 ? _GEN_2088 : _GEN_1812; // @[executor.scala 470:55]
  wire [7:0] _GEN_2581 = opcode_2 != 4'h0 ? _GEN_2089 : _GEN_1813; // @[executor.scala 470:55]
  wire [7:0] _GEN_2582 = opcode_2 != 4'h0 ? _GEN_2090 : _GEN_1814; // @[executor.scala 470:55]
  wire [7:0] _GEN_2583 = opcode_2 != 4'h0 ? _GEN_2091 : _GEN_1815; // @[executor.scala 470:55]
  wire [7:0] _GEN_2584 = opcode_2 != 4'h0 ? _GEN_2096 : _GEN_1816; // @[executor.scala 470:55]
  wire [7:0] _GEN_2585 = opcode_2 != 4'h0 ? _GEN_2097 : _GEN_1817; // @[executor.scala 470:55]
  wire [7:0] _GEN_2586 = opcode_2 != 4'h0 ? _GEN_2098 : _GEN_1818; // @[executor.scala 470:55]
  wire [7:0] _GEN_2587 = opcode_2 != 4'h0 ? _GEN_2099 : _GEN_1819; // @[executor.scala 470:55]
  wire [7:0] _GEN_2588 = opcode_2 != 4'h0 ? _GEN_2104 : _GEN_1820; // @[executor.scala 470:55]
  wire [7:0] _GEN_2589 = opcode_2 != 4'h0 ? _GEN_2105 : _GEN_1821; // @[executor.scala 470:55]
  wire [7:0] _GEN_2590 = opcode_2 != 4'h0 ? _GEN_2106 : _GEN_1822; // @[executor.scala 470:55]
  wire [7:0] _GEN_2591 = opcode_2 != 4'h0 ? _GEN_2107 : _GEN_1823; // @[executor.scala 470:55]
  wire [7:0] _GEN_2592 = opcode_2 != 4'h0 ? _GEN_2112 : _GEN_1824; // @[executor.scala 470:55]
  wire [7:0] _GEN_2593 = opcode_2 != 4'h0 ? _GEN_2113 : _GEN_1825; // @[executor.scala 470:55]
  wire [7:0] _GEN_2594 = opcode_2 != 4'h0 ? _GEN_2114 : _GEN_1826; // @[executor.scala 470:55]
  wire [7:0] _GEN_2595 = opcode_2 != 4'h0 ? _GEN_2115 : _GEN_1827; // @[executor.scala 470:55]
  wire [7:0] _GEN_2596 = opcode_2 != 4'h0 ? _GEN_2120 : _GEN_1828; // @[executor.scala 470:55]
  wire [7:0] _GEN_2597 = opcode_2 != 4'h0 ? _GEN_2121 : _GEN_1829; // @[executor.scala 470:55]
  wire [7:0] _GEN_2598 = opcode_2 != 4'h0 ? _GEN_2122 : _GEN_1830; // @[executor.scala 470:55]
  wire [7:0] _GEN_2599 = opcode_2 != 4'h0 ? _GEN_2123 : _GEN_1831; // @[executor.scala 470:55]
  wire [7:0] _GEN_2600 = opcode_2 != 4'h0 ? _GEN_2128 : _GEN_1832; // @[executor.scala 470:55]
  wire [7:0] _GEN_2601 = opcode_2 != 4'h0 ? _GEN_2129 : _GEN_1833; // @[executor.scala 470:55]
  wire [7:0] _GEN_2602 = opcode_2 != 4'h0 ? _GEN_2130 : _GEN_1834; // @[executor.scala 470:55]
  wire [7:0] _GEN_2603 = opcode_2 != 4'h0 ? _GEN_2131 : _GEN_1835; // @[executor.scala 470:55]
  wire [7:0] _GEN_2604 = opcode_2 != 4'h0 ? _GEN_2136 : _GEN_1836; // @[executor.scala 470:55]
  wire [7:0] _GEN_2605 = opcode_2 != 4'h0 ? _GEN_2137 : _GEN_1837; // @[executor.scala 470:55]
  wire [7:0] _GEN_2606 = opcode_2 != 4'h0 ? _GEN_2138 : _GEN_1838; // @[executor.scala 470:55]
  wire [7:0] _GEN_2607 = opcode_2 != 4'h0 ? _GEN_2139 : _GEN_1839; // @[executor.scala 470:55]
  wire [7:0] _GEN_2608 = opcode_2 != 4'h0 ? _GEN_2144 : _GEN_1840; // @[executor.scala 470:55]
  wire [7:0] _GEN_2609 = opcode_2 != 4'h0 ? _GEN_2145 : _GEN_1841; // @[executor.scala 470:55]
  wire [7:0] _GEN_2610 = opcode_2 != 4'h0 ? _GEN_2146 : _GEN_1842; // @[executor.scala 470:55]
  wire [7:0] _GEN_2611 = opcode_2 != 4'h0 ? _GEN_2147 : _GEN_1843; // @[executor.scala 470:55]
  wire [7:0] _GEN_2612 = opcode_2 != 4'h0 ? _GEN_2152 : _GEN_1844; // @[executor.scala 470:55]
  wire [7:0] _GEN_2613 = opcode_2 != 4'h0 ? _GEN_2153 : _GEN_1845; // @[executor.scala 470:55]
  wire [7:0] _GEN_2614 = opcode_2 != 4'h0 ? _GEN_2154 : _GEN_1846; // @[executor.scala 470:55]
  wire [7:0] _GEN_2615 = opcode_2 != 4'h0 ? _GEN_2155 : _GEN_1847; // @[executor.scala 470:55]
  wire [7:0] _GEN_2616 = opcode_2 != 4'h0 ? _GEN_2160 : _GEN_1848; // @[executor.scala 470:55]
  wire [7:0] _GEN_2617 = opcode_2 != 4'h0 ? _GEN_2161 : _GEN_1849; // @[executor.scala 470:55]
  wire [7:0] _GEN_2618 = opcode_2 != 4'h0 ? _GEN_2162 : _GEN_1850; // @[executor.scala 470:55]
  wire [7:0] _GEN_2619 = opcode_2 != 4'h0 ? _GEN_2163 : _GEN_1851; // @[executor.scala 470:55]
  wire [7:0] _GEN_2620 = opcode_2 != 4'h0 ? _GEN_2168 : _GEN_1852; // @[executor.scala 470:55]
  wire [7:0] _GEN_2621 = opcode_2 != 4'h0 ? _GEN_2169 : _GEN_1853; // @[executor.scala 470:55]
  wire [7:0] _GEN_2622 = opcode_2 != 4'h0 ? _GEN_2170 : _GEN_1854; // @[executor.scala 470:55]
  wire [7:0] _GEN_2623 = opcode_2 != 4'h0 ? _GEN_2171 : _GEN_1855; // @[executor.scala 470:55]
  wire [7:0] _GEN_2624 = opcode_2 != 4'h0 ? _GEN_2176 : _GEN_1856; // @[executor.scala 470:55]
  wire [7:0] _GEN_2625 = opcode_2 != 4'h0 ? _GEN_2177 : _GEN_1857; // @[executor.scala 470:55]
  wire [7:0] _GEN_2626 = opcode_2 != 4'h0 ? _GEN_2178 : _GEN_1858; // @[executor.scala 470:55]
  wire [7:0] _GEN_2627 = opcode_2 != 4'h0 ? _GEN_2179 : _GEN_1859; // @[executor.scala 470:55]
  wire [7:0] _GEN_2628 = opcode_2 != 4'h0 ? _GEN_2184 : _GEN_1860; // @[executor.scala 470:55]
  wire [7:0] _GEN_2629 = opcode_2 != 4'h0 ? _GEN_2185 : _GEN_1861; // @[executor.scala 470:55]
  wire [7:0] _GEN_2630 = opcode_2 != 4'h0 ? _GEN_2186 : _GEN_1862; // @[executor.scala 470:55]
  wire [7:0] _GEN_2631 = opcode_2 != 4'h0 ? _GEN_2187 : _GEN_1863; // @[executor.scala 470:55]
  wire [7:0] _GEN_2632 = opcode_2 != 4'h0 ? _GEN_2192 : _GEN_1864; // @[executor.scala 470:55]
  wire [7:0] _GEN_2633 = opcode_2 != 4'h0 ? _GEN_2193 : _GEN_1865; // @[executor.scala 470:55]
  wire [7:0] _GEN_2634 = opcode_2 != 4'h0 ? _GEN_2194 : _GEN_1866; // @[executor.scala 470:55]
  wire [7:0] _GEN_2635 = opcode_2 != 4'h0 ? _GEN_2195 : _GEN_1867; // @[executor.scala 470:55]
  wire [7:0] _GEN_2636 = opcode_2 != 4'h0 ? _GEN_2200 : _GEN_1868; // @[executor.scala 470:55]
  wire [7:0] _GEN_2637 = opcode_2 != 4'h0 ? _GEN_2201 : _GEN_1869; // @[executor.scala 470:55]
  wire [7:0] _GEN_2638 = opcode_2 != 4'h0 ? _GEN_2202 : _GEN_1870; // @[executor.scala 470:55]
  wire [7:0] _GEN_2639 = opcode_2 != 4'h0 ? _GEN_2203 : _GEN_1871; // @[executor.scala 470:55]
  wire [7:0] _GEN_2640 = opcode_2 != 4'h0 ? _GEN_2208 : _GEN_1872; // @[executor.scala 470:55]
  wire [7:0] _GEN_2641 = opcode_2 != 4'h0 ? _GEN_2209 : _GEN_1873; // @[executor.scala 470:55]
  wire [7:0] _GEN_2642 = opcode_2 != 4'h0 ? _GEN_2210 : _GEN_1874; // @[executor.scala 470:55]
  wire [7:0] _GEN_2643 = opcode_2 != 4'h0 ? _GEN_2211 : _GEN_1875; // @[executor.scala 470:55]
  wire [7:0] _GEN_2644 = opcode_2 != 4'h0 ? _GEN_2216 : _GEN_1876; // @[executor.scala 470:55]
  wire [7:0] _GEN_2645 = opcode_2 != 4'h0 ? _GEN_2217 : _GEN_1877; // @[executor.scala 470:55]
  wire [7:0] _GEN_2646 = opcode_2 != 4'h0 ? _GEN_2218 : _GEN_1878; // @[executor.scala 470:55]
  wire [7:0] _GEN_2647 = opcode_2 != 4'h0 ? _GEN_2219 : _GEN_1879; // @[executor.scala 470:55]
  wire [7:0] _GEN_2648 = opcode_2 != 4'h0 ? _GEN_2224 : _GEN_1880; // @[executor.scala 470:55]
  wire [7:0] _GEN_2649 = opcode_2 != 4'h0 ? _GEN_2225 : _GEN_1881; // @[executor.scala 470:55]
  wire [7:0] _GEN_2650 = opcode_2 != 4'h0 ? _GEN_2226 : _GEN_1882; // @[executor.scala 470:55]
  wire [7:0] _GEN_2651 = opcode_2 != 4'h0 ? _GEN_2227 : _GEN_1883; // @[executor.scala 470:55]
  wire [7:0] _GEN_2652 = opcode_2 != 4'h0 ? _GEN_2232 : _GEN_1884; // @[executor.scala 470:55]
  wire [7:0] _GEN_2653 = opcode_2 != 4'h0 ? _GEN_2233 : _GEN_1885; // @[executor.scala 470:55]
  wire [7:0] _GEN_2654 = opcode_2 != 4'h0 ? _GEN_2234 : _GEN_1886; // @[executor.scala 470:55]
  wire [7:0] _GEN_2655 = opcode_2 != 4'h0 ? _GEN_2235 : _GEN_1887; // @[executor.scala 470:55]
  wire [7:0] _GEN_2656 = opcode_2 != 4'h0 ? _GEN_2240 : _GEN_1888; // @[executor.scala 470:55]
  wire [7:0] _GEN_2657 = opcode_2 != 4'h0 ? _GEN_2241 : _GEN_1889; // @[executor.scala 470:55]
  wire [7:0] _GEN_2658 = opcode_2 != 4'h0 ? _GEN_2242 : _GEN_1890; // @[executor.scala 470:55]
  wire [7:0] _GEN_2659 = opcode_2 != 4'h0 ? _GEN_2243 : _GEN_1891; // @[executor.scala 470:55]
  wire [7:0] _GEN_2660 = opcode_2 != 4'h0 ? _GEN_2248 : _GEN_1892; // @[executor.scala 470:55]
  wire [7:0] _GEN_2661 = opcode_2 != 4'h0 ? _GEN_2249 : _GEN_1893; // @[executor.scala 470:55]
  wire [7:0] _GEN_2662 = opcode_2 != 4'h0 ? _GEN_2250 : _GEN_1894; // @[executor.scala 470:55]
  wire [7:0] _GEN_2663 = opcode_2 != 4'h0 ? _GEN_2251 : _GEN_1895; // @[executor.scala 470:55]
  wire [7:0] _GEN_2664 = opcode_2 != 4'h0 ? _GEN_2256 : _GEN_1896; // @[executor.scala 470:55]
  wire [7:0] _GEN_2665 = opcode_2 != 4'h0 ? _GEN_2257 : _GEN_1897; // @[executor.scala 470:55]
  wire [7:0] _GEN_2666 = opcode_2 != 4'h0 ? _GEN_2258 : _GEN_1898; // @[executor.scala 470:55]
  wire [7:0] _GEN_2667 = opcode_2 != 4'h0 ? _GEN_2259 : _GEN_1899; // @[executor.scala 470:55]
  wire [7:0] _GEN_2668 = opcode_2 != 4'h0 ? _GEN_2264 : _GEN_1900; // @[executor.scala 470:55]
  wire [7:0] _GEN_2669 = opcode_2 != 4'h0 ? _GEN_2265 : _GEN_1901; // @[executor.scala 470:55]
  wire [7:0] _GEN_2670 = opcode_2 != 4'h0 ? _GEN_2266 : _GEN_1902; // @[executor.scala 470:55]
  wire [7:0] _GEN_2671 = opcode_2 != 4'h0 ? _GEN_2267 : _GEN_1903; // @[executor.scala 470:55]
  wire [7:0] _GEN_2672 = opcode_2 != 4'h0 ? _GEN_2272 : _GEN_1904; // @[executor.scala 470:55]
  wire [7:0] _GEN_2673 = opcode_2 != 4'h0 ? _GEN_2273 : _GEN_1905; // @[executor.scala 470:55]
  wire [7:0] _GEN_2674 = opcode_2 != 4'h0 ? _GEN_2274 : _GEN_1906; // @[executor.scala 470:55]
  wire [7:0] _GEN_2675 = opcode_2 != 4'h0 ? _GEN_2275 : _GEN_1907; // @[executor.scala 470:55]
  wire [7:0] _GEN_2676 = opcode_2 != 4'h0 ? _GEN_2280 : _GEN_1908; // @[executor.scala 470:55]
  wire [7:0] _GEN_2677 = opcode_2 != 4'h0 ? _GEN_2281 : _GEN_1909; // @[executor.scala 470:55]
  wire [7:0] _GEN_2678 = opcode_2 != 4'h0 ? _GEN_2282 : _GEN_1910; // @[executor.scala 470:55]
  wire [7:0] _GEN_2679 = opcode_2 != 4'h0 ? _GEN_2283 : _GEN_1911; // @[executor.scala 470:55]
  wire [7:0] _GEN_2680 = opcode_2 != 4'h0 ? _GEN_2288 : _GEN_1912; // @[executor.scala 470:55]
  wire [7:0] _GEN_2681 = opcode_2 != 4'h0 ? _GEN_2289 : _GEN_1913; // @[executor.scala 470:55]
  wire [7:0] _GEN_2682 = opcode_2 != 4'h0 ? _GEN_2290 : _GEN_1914; // @[executor.scala 470:55]
  wire [7:0] _GEN_2683 = opcode_2 != 4'h0 ? _GEN_2291 : _GEN_1915; // @[executor.scala 470:55]
  wire [7:0] _GEN_2684 = opcode_2 != 4'h0 ? _GEN_2296 : _GEN_1916; // @[executor.scala 470:55]
  wire [7:0] _GEN_2685 = opcode_2 != 4'h0 ? _GEN_2297 : _GEN_1917; // @[executor.scala 470:55]
  wire [7:0] _GEN_2686 = opcode_2 != 4'h0 ? _GEN_2298 : _GEN_1918; // @[executor.scala 470:55]
  wire [7:0] _GEN_2687 = opcode_2 != 4'h0 ? _GEN_2299 : _GEN_1919; // @[executor.scala 470:55]
  wire [7:0] _GEN_2688 = opcode_2 != 4'h0 ? _GEN_2304 : _GEN_1920; // @[executor.scala 470:55]
  wire [7:0] _GEN_2689 = opcode_2 != 4'h0 ? _GEN_2305 : _GEN_1921; // @[executor.scala 470:55]
  wire [7:0] _GEN_2690 = opcode_2 != 4'h0 ? _GEN_2306 : _GEN_1922; // @[executor.scala 470:55]
  wire [7:0] _GEN_2691 = opcode_2 != 4'h0 ? _GEN_2307 : _GEN_1923; // @[executor.scala 470:55]
  wire [7:0] _GEN_2692 = opcode_2 != 4'h0 ? _GEN_2312 : _GEN_1924; // @[executor.scala 470:55]
  wire [7:0] _GEN_2693 = opcode_2 != 4'h0 ? _GEN_2313 : _GEN_1925; // @[executor.scala 470:55]
  wire [7:0] _GEN_2694 = opcode_2 != 4'h0 ? _GEN_2314 : _GEN_1926; // @[executor.scala 470:55]
  wire [7:0] _GEN_2695 = opcode_2 != 4'h0 ? _GEN_2315 : _GEN_1927; // @[executor.scala 470:55]
  wire [7:0] _GEN_2696 = opcode_2 != 4'h0 ? _GEN_2320 : _GEN_1928; // @[executor.scala 470:55]
  wire [7:0] _GEN_2697 = opcode_2 != 4'h0 ? _GEN_2321 : _GEN_1929; // @[executor.scala 470:55]
  wire [7:0] _GEN_2698 = opcode_2 != 4'h0 ? _GEN_2322 : _GEN_1930; // @[executor.scala 470:55]
  wire [7:0] _GEN_2699 = opcode_2 != 4'h0 ? _GEN_2323 : _GEN_1931; // @[executor.scala 470:55]
  wire [7:0] _GEN_2700 = opcode_2 != 4'h0 ? _GEN_2328 : _GEN_1932; // @[executor.scala 470:55]
  wire [7:0] _GEN_2701 = opcode_2 != 4'h0 ? _GEN_2329 : _GEN_1933; // @[executor.scala 470:55]
  wire [7:0] _GEN_2702 = opcode_2 != 4'h0 ? _GEN_2330 : _GEN_1934; // @[executor.scala 470:55]
  wire [7:0] _GEN_2703 = opcode_2 != 4'h0 ? _GEN_2331 : _GEN_1935; // @[executor.scala 470:55]
  wire [7:0] _GEN_2704 = opcode_2 != 4'h0 ? _GEN_2336 : _GEN_1936; // @[executor.scala 470:55]
  wire [7:0] _GEN_2705 = opcode_2 != 4'h0 ? _GEN_2337 : _GEN_1937; // @[executor.scala 470:55]
  wire [7:0] _GEN_2706 = opcode_2 != 4'h0 ? _GEN_2338 : _GEN_1938; // @[executor.scala 470:55]
  wire [7:0] _GEN_2707 = opcode_2 != 4'h0 ? _GEN_2339 : _GEN_1939; // @[executor.scala 470:55]
  wire [7:0] _GEN_2708 = opcode_2 != 4'h0 ? _GEN_2344 : _GEN_1940; // @[executor.scala 470:55]
  wire [7:0] _GEN_2709 = opcode_2 != 4'h0 ? _GEN_2345 : _GEN_1941; // @[executor.scala 470:55]
  wire [7:0] _GEN_2710 = opcode_2 != 4'h0 ? _GEN_2346 : _GEN_1942; // @[executor.scala 470:55]
  wire [7:0] _GEN_2711 = opcode_2 != 4'h0 ? _GEN_2347 : _GEN_1943; // @[executor.scala 470:55]
  wire [7:0] _GEN_2712 = opcode_2 != 4'h0 ? _GEN_2352 : _GEN_1944; // @[executor.scala 470:55]
  wire [7:0] _GEN_2713 = opcode_2 != 4'h0 ? _GEN_2353 : _GEN_1945; // @[executor.scala 470:55]
  wire [7:0] _GEN_2714 = opcode_2 != 4'h0 ? _GEN_2354 : _GEN_1946; // @[executor.scala 470:55]
  wire [7:0] _GEN_2715 = opcode_2 != 4'h0 ? _GEN_2355 : _GEN_1947; // @[executor.scala 470:55]
  wire [7:0] _GEN_2716 = opcode_2 != 4'h0 ? _GEN_2360 : _GEN_1948; // @[executor.scala 470:55]
  wire [7:0] _GEN_2717 = opcode_2 != 4'h0 ? _GEN_2361 : _GEN_1949; // @[executor.scala 470:55]
  wire [7:0] _GEN_2718 = opcode_2 != 4'h0 ? _GEN_2362 : _GEN_1950; // @[executor.scala 470:55]
  wire [7:0] _GEN_2719 = opcode_2 != 4'h0 ? _GEN_2363 : _GEN_1951; // @[executor.scala 470:55]
  wire [7:0] _GEN_2720 = opcode_2 != 4'h0 ? _GEN_2368 : _GEN_1952; // @[executor.scala 470:55]
  wire [7:0] _GEN_2721 = opcode_2 != 4'h0 ? _GEN_2369 : _GEN_1953; // @[executor.scala 470:55]
  wire [7:0] _GEN_2722 = opcode_2 != 4'h0 ? _GEN_2370 : _GEN_1954; // @[executor.scala 470:55]
  wire [7:0] _GEN_2723 = opcode_2 != 4'h0 ? _GEN_2371 : _GEN_1955; // @[executor.scala 470:55]
  wire [7:0] _GEN_2724 = opcode_2 != 4'h0 ? _GEN_2376 : _GEN_1956; // @[executor.scala 470:55]
  wire [7:0] _GEN_2725 = opcode_2 != 4'h0 ? _GEN_2377 : _GEN_1957; // @[executor.scala 470:55]
  wire [7:0] _GEN_2726 = opcode_2 != 4'h0 ? _GEN_2378 : _GEN_1958; // @[executor.scala 470:55]
  wire [7:0] _GEN_2727 = opcode_2 != 4'h0 ? _GEN_2379 : _GEN_1959; // @[executor.scala 470:55]
  wire [7:0] _GEN_2728 = opcode_2 != 4'h0 ? _GEN_2384 : _GEN_1960; // @[executor.scala 470:55]
  wire [7:0] _GEN_2729 = opcode_2 != 4'h0 ? _GEN_2385 : _GEN_1961; // @[executor.scala 470:55]
  wire [7:0] _GEN_2730 = opcode_2 != 4'h0 ? _GEN_2386 : _GEN_1962; // @[executor.scala 470:55]
  wire [7:0] _GEN_2731 = opcode_2 != 4'h0 ? _GEN_2387 : _GEN_1963; // @[executor.scala 470:55]
  wire [7:0] _GEN_2732 = opcode_2 != 4'h0 ? _GEN_2392 : _GEN_1964; // @[executor.scala 470:55]
  wire [7:0] _GEN_2733 = opcode_2 != 4'h0 ? _GEN_2393 : _GEN_1965; // @[executor.scala 470:55]
  wire [7:0] _GEN_2734 = opcode_2 != 4'h0 ? _GEN_2394 : _GEN_1966; // @[executor.scala 470:55]
  wire [7:0] _GEN_2735 = opcode_2 != 4'h0 ? _GEN_2395 : _GEN_1967; // @[executor.scala 470:55]
  wire [7:0] _GEN_2736 = opcode_2 != 4'h0 ? _GEN_2400 : _GEN_1968; // @[executor.scala 470:55]
  wire [7:0] _GEN_2737 = opcode_2 != 4'h0 ? _GEN_2401 : _GEN_1969; // @[executor.scala 470:55]
  wire [7:0] _GEN_2738 = opcode_2 != 4'h0 ? _GEN_2402 : _GEN_1970; // @[executor.scala 470:55]
  wire [7:0] _GEN_2739 = opcode_2 != 4'h0 ? _GEN_2403 : _GEN_1971; // @[executor.scala 470:55]
  wire [7:0] _GEN_2740 = opcode_2 != 4'h0 ? _GEN_2408 : _GEN_1972; // @[executor.scala 470:55]
  wire [7:0] _GEN_2741 = opcode_2 != 4'h0 ? _GEN_2409 : _GEN_1973; // @[executor.scala 470:55]
  wire [7:0] _GEN_2742 = opcode_2 != 4'h0 ? _GEN_2410 : _GEN_1974; // @[executor.scala 470:55]
  wire [7:0] _GEN_2743 = opcode_2 != 4'h0 ? _GEN_2411 : _GEN_1975; // @[executor.scala 470:55]
  wire [7:0] _GEN_2744 = opcode_2 != 4'h0 ? _GEN_2416 : _GEN_1976; // @[executor.scala 470:55]
  wire [7:0] _GEN_2745 = opcode_2 != 4'h0 ? _GEN_2417 : _GEN_1977; // @[executor.scala 470:55]
  wire [7:0] _GEN_2746 = opcode_2 != 4'h0 ? _GEN_2418 : _GEN_1978; // @[executor.scala 470:55]
  wire [7:0] _GEN_2747 = opcode_2 != 4'h0 ? _GEN_2419 : _GEN_1979; // @[executor.scala 470:55]
  wire [7:0] _GEN_2748 = opcode_2 != 4'h0 ? _GEN_2424 : _GEN_1980; // @[executor.scala 470:55]
  wire [7:0] _GEN_2749 = opcode_2 != 4'h0 ? _GEN_2425 : _GEN_1981; // @[executor.scala 470:55]
  wire [7:0] _GEN_2750 = opcode_2 != 4'h0 ? _GEN_2426 : _GEN_1982; // @[executor.scala 470:55]
  wire [7:0] _GEN_2751 = opcode_2 != 4'h0 ? _GEN_2427 : _GEN_1983; // @[executor.scala 470:55]
  wire [7:0] _GEN_2752 = opcode_2 != 4'h0 ? _GEN_2432 : _GEN_1984; // @[executor.scala 470:55]
  wire [7:0] _GEN_2753 = opcode_2 != 4'h0 ? _GEN_2433 : _GEN_1985; // @[executor.scala 470:55]
  wire [7:0] _GEN_2754 = opcode_2 != 4'h0 ? _GEN_2434 : _GEN_1986; // @[executor.scala 470:55]
  wire [7:0] _GEN_2755 = opcode_2 != 4'h0 ? _GEN_2435 : _GEN_1987; // @[executor.scala 470:55]
  wire [7:0] _GEN_2756 = opcode_2 != 4'h0 ? _GEN_2440 : _GEN_1988; // @[executor.scala 470:55]
  wire [7:0] _GEN_2757 = opcode_2 != 4'h0 ? _GEN_2441 : _GEN_1989; // @[executor.scala 470:55]
  wire [7:0] _GEN_2758 = opcode_2 != 4'h0 ? _GEN_2442 : _GEN_1990; // @[executor.scala 470:55]
  wire [7:0] _GEN_2759 = opcode_2 != 4'h0 ? _GEN_2443 : _GEN_1991; // @[executor.scala 470:55]
  wire [7:0] _GEN_2760 = opcode_2 != 4'h0 ? _GEN_2448 : _GEN_1992; // @[executor.scala 470:55]
  wire [7:0] _GEN_2761 = opcode_2 != 4'h0 ? _GEN_2449 : _GEN_1993; // @[executor.scala 470:55]
  wire [7:0] _GEN_2762 = opcode_2 != 4'h0 ? _GEN_2450 : _GEN_1994; // @[executor.scala 470:55]
  wire [7:0] _GEN_2763 = opcode_2 != 4'h0 ? _GEN_2451 : _GEN_1995; // @[executor.scala 470:55]
  wire [7:0] _GEN_2764 = opcode_2 != 4'h0 ? _GEN_2456 : _GEN_1996; // @[executor.scala 470:55]
  wire [7:0] _GEN_2765 = opcode_2 != 4'h0 ? _GEN_2457 : _GEN_1997; // @[executor.scala 470:55]
  wire [7:0] _GEN_2766 = opcode_2 != 4'h0 ? _GEN_2458 : _GEN_1998; // @[executor.scala 470:55]
  wire [7:0] _GEN_2767 = opcode_2 != 4'h0 ? _GEN_2459 : _GEN_1999; // @[executor.scala 470:55]
  wire [7:0] _GEN_2768 = opcode_2 != 4'h0 ? _GEN_2464 : _GEN_2000; // @[executor.scala 470:55]
  wire [7:0] _GEN_2769 = opcode_2 != 4'h0 ? _GEN_2465 : _GEN_2001; // @[executor.scala 470:55]
  wire [7:0] _GEN_2770 = opcode_2 != 4'h0 ? _GEN_2466 : _GEN_2002; // @[executor.scala 470:55]
  wire [7:0] _GEN_2771 = opcode_2 != 4'h0 ? _GEN_2467 : _GEN_2003; // @[executor.scala 470:55]
  wire [7:0] _GEN_2772 = opcode_2 != 4'h0 ? _GEN_2472 : _GEN_2004; // @[executor.scala 470:55]
  wire [7:0] _GEN_2773 = opcode_2 != 4'h0 ? _GEN_2473 : _GEN_2005; // @[executor.scala 470:55]
  wire [7:0] _GEN_2774 = opcode_2 != 4'h0 ? _GEN_2474 : _GEN_2006; // @[executor.scala 470:55]
  wire [7:0] _GEN_2775 = opcode_2 != 4'h0 ? _GEN_2475 : _GEN_2007; // @[executor.scala 470:55]
  wire [7:0] _GEN_2776 = opcode_2 != 4'h0 ? _GEN_2480 : _GEN_2008; // @[executor.scala 470:55]
  wire [7:0] _GEN_2777 = opcode_2 != 4'h0 ? _GEN_2481 : _GEN_2009; // @[executor.scala 470:55]
  wire [7:0] _GEN_2778 = opcode_2 != 4'h0 ? _GEN_2482 : _GEN_2010; // @[executor.scala 470:55]
  wire [7:0] _GEN_2779 = opcode_2 != 4'h0 ? _GEN_2483 : _GEN_2011; // @[executor.scala 470:55]
  wire [7:0] _GEN_2780 = opcode_2 != 4'h0 ? _GEN_2488 : _GEN_2012; // @[executor.scala 470:55]
  wire [7:0] _GEN_2781 = opcode_2 != 4'h0 ? _GEN_2489 : _GEN_2013; // @[executor.scala 470:55]
  wire [7:0] _GEN_2782 = opcode_2 != 4'h0 ? _GEN_2490 : _GEN_2014; // @[executor.scala 470:55]
  wire [7:0] _GEN_2783 = opcode_2 != 4'h0 ? _GEN_2491 : _GEN_2015; // @[executor.scala 470:55]
  wire [7:0] _GEN_2784 = opcode_2 != 4'h0 ? _GEN_2496 : _GEN_2016; // @[executor.scala 470:55]
  wire [7:0] _GEN_2785 = opcode_2 != 4'h0 ? _GEN_2497 : _GEN_2017; // @[executor.scala 470:55]
  wire [7:0] _GEN_2786 = opcode_2 != 4'h0 ? _GEN_2498 : _GEN_2018; // @[executor.scala 470:55]
  wire [7:0] _GEN_2787 = opcode_2 != 4'h0 ? _GEN_2499 : _GEN_2019; // @[executor.scala 470:55]
  wire [7:0] _GEN_2788 = opcode_2 != 4'h0 ? _GEN_2504 : _GEN_2020; // @[executor.scala 470:55]
  wire [7:0] _GEN_2789 = opcode_2 != 4'h0 ? _GEN_2505 : _GEN_2021; // @[executor.scala 470:55]
  wire [7:0] _GEN_2790 = opcode_2 != 4'h0 ? _GEN_2506 : _GEN_2022; // @[executor.scala 470:55]
  wire [7:0] _GEN_2791 = opcode_2 != 4'h0 ? _GEN_2507 : _GEN_2023; // @[executor.scala 470:55]
  wire [7:0] _GEN_2792 = opcode_2 != 4'h0 ? _GEN_2512 : _GEN_2024; // @[executor.scala 470:55]
  wire [7:0] _GEN_2793 = opcode_2 != 4'h0 ? _GEN_2513 : _GEN_2025; // @[executor.scala 470:55]
  wire [7:0] _GEN_2794 = opcode_2 != 4'h0 ? _GEN_2514 : _GEN_2026; // @[executor.scala 470:55]
  wire [7:0] _GEN_2795 = opcode_2 != 4'h0 ? _GEN_2515 : _GEN_2027; // @[executor.scala 470:55]
  wire [7:0] _GEN_2796 = opcode_2 != 4'h0 ? _GEN_2520 : _GEN_2028; // @[executor.scala 470:55]
  wire [7:0] _GEN_2797 = opcode_2 != 4'h0 ? _GEN_2521 : _GEN_2029; // @[executor.scala 470:55]
  wire [7:0] _GEN_2798 = opcode_2 != 4'h0 ? _GEN_2522 : _GEN_2030; // @[executor.scala 470:55]
  wire [7:0] _GEN_2799 = opcode_2 != 4'h0 ? _GEN_2523 : _GEN_2031; // @[executor.scala 470:55]
  wire [7:0] _GEN_2800 = opcode_2 != 4'h0 ? _GEN_2528 : _GEN_2032; // @[executor.scala 470:55]
  wire [7:0] _GEN_2801 = opcode_2 != 4'h0 ? _GEN_2529 : _GEN_2033; // @[executor.scala 470:55]
  wire [7:0] _GEN_2802 = opcode_2 != 4'h0 ? _GEN_2530 : _GEN_2034; // @[executor.scala 470:55]
  wire [7:0] _GEN_2803 = opcode_2 != 4'h0 ? _GEN_2531 : _GEN_2035; // @[executor.scala 470:55]
  wire [7:0] _GEN_2804 = opcode_2 != 4'h0 ? _GEN_2536 : _GEN_2036; // @[executor.scala 470:55]
  wire [7:0] _GEN_2805 = opcode_2 != 4'h0 ? _GEN_2537 : _GEN_2037; // @[executor.scala 470:55]
  wire [7:0] _GEN_2806 = opcode_2 != 4'h0 ? _GEN_2538 : _GEN_2038; // @[executor.scala 470:55]
  wire [7:0] _GEN_2807 = opcode_2 != 4'h0 ? _GEN_2539 : _GEN_2039; // @[executor.scala 470:55]
  wire [7:0] _GEN_2808 = opcode_2 != 4'h0 ? _GEN_2544 : _GEN_2040; // @[executor.scala 470:55]
  wire [7:0] _GEN_2809 = opcode_2 != 4'h0 ? _GEN_2545 : _GEN_2041; // @[executor.scala 470:55]
  wire [7:0] _GEN_2810 = opcode_2 != 4'h0 ? _GEN_2546 : _GEN_2042; // @[executor.scala 470:55]
  wire [7:0] _GEN_2811 = opcode_2 != 4'h0 ? _GEN_2547 : _GEN_2043; // @[executor.scala 470:55]
  wire [7:0] _GEN_2812 = opcode_2 != 4'h0 ? _GEN_2552 : _GEN_2044; // @[executor.scala 470:55]
  wire [7:0] _GEN_2813 = opcode_2 != 4'h0 ? _GEN_2553 : _GEN_2045; // @[executor.scala 470:55]
  wire [7:0] _GEN_2814 = opcode_2 != 4'h0 ? _GEN_2554 : _GEN_2046; // @[executor.scala 470:55]
  wire [7:0] _GEN_2815 = opcode_2 != 4'h0 ? _GEN_2555 : _GEN_2047; // @[executor.scala 470:55]
  wire [7:0] _GEN_2816 = opcode_2 != 4'h0 ? _GEN_2560 : _GEN_2048; // @[executor.scala 470:55]
  wire [7:0] _GEN_2817 = opcode_2 != 4'h0 ? _GEN_2561 : _GEN_2049; // @[executor.scala 470:55]
  wire [7:0] _GEN_2818 = opcode_2 != 4'h0 ? _GEN_2562 : _GEN_2050; // @[executor.scala 470:55]
  wire [7:0] _GEN_2819 = opcode_2 != 4'h0 ? _GEN_2563 : _GEN_2051; // @[executor.scala 470:55]
  wire [7:0] _GEN_2822 = opcode_2 == 4'hf ? _GEN_1796 : _GEN_2564; // @[executor.scala 466:52]
  wire [7:0] _GEN_2823 = opcode_2 == 4'hf ? _GEN_1797 : _GEN_2565; // @[executor.scala 466:52]
  wire [7:0] _GEN_2824 = opcode_2 == 4'hf ? _GEN_1798 : _GEN_2566; // @[executor.scala 466:52]
  wire [7:0] _GEN_2825 = opcode_2 == 4'hf ? _GEN_1799 : _GEN_2567; // @[executor.scala 466:52]
  wire [7:0] _GEN_2826 = opcode_2 == 4'hf ? _GEN_1800 : _GEN_2568; // @[executor.scala 466:52]
  wire [7:0] _GEN_2827 = opcode_2 == 4'hf ? _GEN_1801 : _GEN_2569; // @[executor.scala 466:52]
  wire [7:0] _GEN_2828 = opcode_2 == 4'hf ? _GEN_1802 : _GEN_2570; // @[executor.scala 466:52]
  wire [7:0] _GEN_2829 = opcode_2 == 4'hf ? _GEN_1803 : _GEN_2571; // @[executor.scala 466:52]
  wire [7:0] _GEN_2830 = opcode_2 == 4'hf ? _GEN_1804 : _GEN_2572; // @[executor.scala 466:52]
  wire [7:0] _GEN_2831 = opcode_2 == 4'hf ? _GEN_1805 : _GEN_2573; // @[executor.scala 466:52]
  wire [7:0] _GEN_2832 = opcode_2 == 4'hf ? _GEN_1806 : _GEN_2574; // @[executor.scala 466:52]
  wire [7:0] _GEN_2833 = opcode_2 == 4'hf ? _GEN_1807 : _GEN_2575; // @[executor.scala 466:52]
  wire [7:0] _GEN_2834 = opcode_2 == 4'hf ? _GEN_1808 : _GEN_2576; // @[executor.scala 466:52]
  wire [7:0] _GEN_2835 = opcode_2 == 4'hf ? _GEN_1809 : _GEN_2577; // @[executor.scala 466:52]
  wire [7:0] _GEN_2836 = opcode_2 == 4'hf ? _GEN_1810 : _GEN_2578; // @[executor.scala 466:52]
  wire [7:0] _GEN_2837 = opcode_2 == 4'hf ? _GEN_1811 : _GEN_2579; // @[executor.scala 466:52]
  wire [7:0] _GEN_2838 = opcode_2 == 4'hf ? _GEN_1812 : _GEN_2580; // @[executor.scala 466:52]
  wire [7:0] _GEN_2839 = opcode_2 == 4'hf ? _GEN_1813 : _GEN_2581; // @[executor.scala 466:52]
  wire [7:0] _GEN_2840 = opcode_2 == 4'hf ? _GEN_1814 : _GEN_2582; // @[executor.scala 466:52]
  wire [7:0] _GEN_2841 = opcode_2 == 4'hf ? _GEN_1815 : _GEN_2583; // @[executor.scala 466:52]
  wire [7:0] _GEN_2842 = opcode_2 == 4'hf ? _GEN_1816 : _GEN_2584; // @[executor.scala 466:52]
  wire [7:0] _GEN_2843 = opcode_2 == 4'hf ? _GEN_1817 : _GEN_2585; // @[executor.scala 466:52]
  wire [7:0] _GEN_2844 = opcode_2 == 4'hf ? _GEN_1818 : _GEN_2586; // @[executor.scala 466:52]
  wire [7:0] _GEN_2845 = opcode_2 == 4'hf ? _GEN_1819 : _GEN_2587; // @[executor.scala 466:52]
  wire [7:0] _GEN_2846 = opcode_2 == 4'hf ? _GEN_1820 : _GEN_2588; // @[executor.scala 466:52]
  wire [7:0] _GEN_2847 = opcode_2 == 4'hf ? _GEN_1821 : _GEN_2589; // @[executor.scala 466:52]
  wire [7:0] _GEN_2848 = opcode_2 == 4'hf ? _GEN_1822 : _GEN_2590; // @[executor.scala 466:52]
  wire [7:0] _GEN_2849 = opcode_2 == 4'hf ? _GEN_1823 : _GEN_2591; // @[executor.scala 466:52]
  wire [7:0] _GEN_2850 = opcode_2 == 4'hf ? _GEN_1824 : _GEN_2592; // @[executor.scala 466:52]
  wire [7:0] _GEN_2851 = opcode_2 == 4'hf ? _GEN_1825 : _GEN_2593; // @[executor.scala 466:52]
  wire [7:0] _GEN_2852 = opcode_2 == 4'hf ? _GEN_1826 : _GEN_2594; // @[executor.scala 466:52]
  wire [7:0] _GEN_2853 = opcode_2 == 4'hf ? _GEN_1827 : _GEN_2595; // @[executor.scala 466:52]
  wire [7:0] _GEN_2854 = opcode_2 == 4'hf ? _GEN_1828 : _GEN_2596; // @[executor.scala 466:52]
  wire [7:0] _GEN_2855 = opcode_2 == 4'hf ? _GEN_1829 : _GEN_2597; // @[executor.scala 466:52]
  wire [7:0] _GEN_2856 = opcode_2 == 4'hf ? _GEN_1830 : _GEN_2598; // @[executor.scala 466:52]
  wire [7:0] _GEN_2857 = opcode_2 == 4'hf ? _GEN_1831 : _GEN_2599; // @[executor.scala 466:52]
  wire [7:0] _GEN_2858 = opcode_2 == 4'hf ? _GEN_1832 : _GEN_2600; // @[executor.scala 466:52]
  wire [7:0] _GEN_2859 = opcode_2 == 4'hf ? _GEN_1833 : _GEN_2601; // @[executor.scala 466:52]
  wire [7:0] _GEN_2860 = opcode_2 == 4'hf ? _GEN_1834 : _GEN_2602; // @[executor.scala 466:52]
  wire [7:0] _GEN_2861 = opcode_2 == 4'hf ? _GEN_1835 : _GEN_2603; // @[executor.scala 466:52]
  wire [7:0] _GEN_2862 = opcode_2 == 4'hf ? _GEN_1836 : _GEN_2604; // @[executor.scala 466:52]
  wire [7:0] _GEN_2863 = opcode_2 == 4'hf ? _GEN_1837 : _GEN_2605; // @[executor.scala 466:52]
  wire [7:0] _GEN_2864 = opcode_2 == 4'hf ? _GEN_1838 : _GEN_2606; // @[executor.scala 466:52]
  wire [7:0] _GEN_2865 = opcode_2 == 4'hf ? _GEN_1839 : _GEN_2607; // @[executor.scala 466:52]
  wire [7:0] _GEN_2866 = opcode_2 == 4'hf ? _GEN_1840 : _GEN_2608; // @[executor.scala 466:52]
  wire [7:0] _GEN_2867 = opcode_2 == 4'hf ? _GEN_1841 : _GEN_2609; // @[executor.scala 466:52]
  wire [7:0] _GEN_2868 = opcode_2 == 4'hf ? _GEN_1842 : _GEN_2610; // @[executor.scala 466:52]
  wire [7:0] _GEN_2869 = opcode_2 == 4'hf ? _GEN_1843 : _GEN_2611; // @[executor.scala 466:52]
  wire [7:0] _GEN_2870 = opcode_2 == 4'hf ? _GEN_1844 : _GEN_2612; // @[executor.scala 466:52]
  wire [7:0] _GEN_2871 = opcode_2 == 4'hf ? _GEN_1845 : _GEN_2613; // @[executor.scala 466:52]
  wire [7:0] _GEN_2872 = opcode_2 == 4'hf ? _GEN_1846 : _GEN_2614; // @[executor.scala 466:52]
  wire [7:0] _GEN_2873 = opcode_2 == 4'hf ? _GEN_1847 : _GEN_2615; // @[executor.scala 466:52]
  wire [7:0] _GEN_2874 = opcode_2 == 4'hf ? _GEN_1848 : _GEN_2616; // @[executor.scala 466:52]
  wire [7:0] _GEN_2875 = opcode_2 == 4'hf ? _GEN_1849 : _GEN_2617; // @[executor.scala 466:52]
  wire [7:0] _GEN_2876 = opcode_2 == 4'hf ? _GEN_1850 : _GEN_2618; // @[executor.scala 466:52]
  wire [7:0] _GEN_2877 = opcode_2 == 4'hf ? _GEN_1851 : _GEN_2619; // @[executor.scala 466:52]
  wire [7:0] _GEN_2878 = opcode_2 == 4'hf ? _GEN_1852 : _GEN_2620; // @[executor.scala 466:52]
  wire [7:0] _GEN_2879 = opcode_2 == 4'hf ? _GEN_1853 : _GEN_2621; // @[executor.scala 466:52]
  wire [7:0] _GEN_2880 = opcode_2 == 4'hf ? _GEN_1854 : _GEN_2622; // @[executor.scala 466:52]
  wire [7:0] _GEN_2881 = opcode_2 == 4'hf ? _GEN_1855 : _GEN_2623; // @[executor.scala 466:52]
  wire [7:0] _GEN_2882 = opcode_2 == 4'hf ? _GEN_1856 : _GEN_2624; // @[executor.scala 466:52]
  wire [7:0] _GEN_2883 = opcode_2 == 4'hf ? _GEN_1857 : _GEN_2625; // @[executor.scala 466:52]
  wire [7:0] _GEN_2884 = opcode_2 == 4'hf ? _GEN_1858 : _GEN_2626; // @[executor.scala 466:52]
  wire [7:0] _GEN_2885 = opcode_2 == 4'hf ? _GEN_1859 : _GEN_2627; // @[executor.scala 466:52]
  wire [7:0] _GEN_2886 = opcode_2 == 4'hf ? _GEN_1860 : _GEN_2628; // @[executor.scala 466:52]
  wire [7:0] _GEN_2887 = opcode_2 == 4'hf ? _GEN_1861 : _GEN_2629; // @[executor.scala 466:52]
  wire [7:0] _GEN_2888 = opcode_2 == 4'hf ? _GEN_1862 : _GEN_2630; // @[executor.scala 466:52]
  wire [7:0] _GEN_2889 = opcode_2 == 4'hf ? _GEN_1863 : _GEN_2631; // @[executor.scala 466:52]
  wire [7:0] _GEN_2890 = opcode_2 == 4'hf ? _GEN_1864 : _GEN_2632; // @[executor.scala 466:52]
  wire [7:0] _GEN_2891 = opcode_2 == 4'hf ? _GEN_1865 : _GEN_2633; // @[executor.scala 466:52]
  wire [7:0] _GEN_2892 = opcode_2 == 4'hf ? _GEN_1866 : _GEN_2634; // @[executor.scala 466:52]
  wire [7:0] _GEN_2893 = opcode_2 == 4'hf ? _GEN_1867 : _GEN_2635; // @[executor.scala 466:52]
  wire [7:0] _GEN_2894 = opcode_2 == 4'hf ? _GEN_1868 : _GEN_2636; // @[executor.scala 466:52]
  wire [7:0] _GEN_2895 = opcode_2 == 4'hf ? _GEN_1869 : _GEN_2637; // @[executor.scala 466:52]
  wire [7:0] _GEN_2896 = opcode_2 == 4'hf ? _GEN_1870 : _GEN_2638; // @[executor.scala 466:52]
  wire [7:0] _GEN_2897 = opcode_2 == 4'hf ? _GEN_1871 : _GEN_2639; // @[executor.scala 466:52]
  wire [7:0] _GEN_2898 = opcode_2 == 4'hf ? _GEN_1872 : _GEN_2640; // @[executor.scala 466:52]
  wire [7:0] _GEN_2899 = opcode_2 == 4'hf ? _GEN_1873 : _GEN_2641; // @[executor.scala 466:52]
  wire [7:0] _GEN_2900 = opcode_2 == 4'hf ? _GEN_1874 : _GEN_2642; // @[executor.scala 466:52]
  wire [7:0] _GEN_2901 = opcode_2 == 4'hf ? _GEN_1875 : _GEN_2643; // @[executor.scala 466:52]
  wire [7:0] _GEN_2902 = opcode_2 == 4'hf ? _GEN_1876 : _GEN_2644; // @[executor.scala 466:52]
  wire [7:0] _GEN_2903 = opcode_2 == 4'hf ? _GEN_1877 : _GEN_2645; // @[executor.scala 466:52]
  wire [7:0] _GEN_2904 = opcode_2 == 4'hf ? _GEN_1878 : _GEN_2646; // @[executor.scala 466:52]
  wire [7:0] _GEN_2905 = opcode_2 == 4'hf ? _GEN_1879 : _GEN_2647; // @[executor.scala 466:52]
  wire [7:0] _GEN_2906 = opcode_2 == 4'hf ? _GEN_1880 : _GEN_2648; // @[executor.scala 466:52]
  wire [7:0] _GEN_2907 = opcode_2 == 4'hf ? _GEN_1881 : _GEN_2649; // @[executor.scala 466:52]
  wire [7:0] _GEN_2908 = opcode_2 == 4'hf ? _GEN_1882 : _GEN_2650; // @[executor.scala 466:52]
  wire [7:0] _GEN_2909 = opcode_2 == 4'hf ? _GEN_1883 : _GEN_2651; // @[executor.scala 466:52]
  wire [7:0] _GEN_2910 = opcode_2 == 4'hf ? _GEN_1884 : _GEN_2652; // @[executor.scala 466:52]
  wire [7:0] _GEN_2911 = opcode_2 == 4'hf ? _GEN_1885 : _GEN_2653; // @[executor.scala 466:52]
  wire [7:0] _GEN_2912 = opcode_2 == 4'hf ? _GEN_1886 : _GEN_2654; // @[executor.scala 466:52]
  wire [7:0] _GEN_2913 = opcode_2 == 4'hf ? _GEN_1887 : _GEN_2655; // @[executor.scala 466:52]
  wire [7:0] _GEN_2914 = opcode_2 == 4'hf ? _GEN_1888 : _GEN_2656; // @[executor.scala 466:52]
  wire [7:0] _GEN_2915 = opcode_2 == 4'hf ? _GEN_1889 : _GEN_2657; // @[executor.scala 466:52]
  wire [7:0] _GEN_2916 = opcode_2 == 4'hf ? _GEN_1890 : _GEN_2658; // @[executor.scala 466:52]
  wire [7:0] _GEN_2917 = opcode_2 == 4'hf ? _GEN_1891 : _GEN_2659; // @[executor.scala 466:52]
  wire [7:0] _GEN_2918 = opcode_2 == 4'hf ? _GEN_1892 : _GEN_2660; // @[executor.scala 466:52]
  wire [7:0] _GEN_2919 = opcode_2 == 4'hf ? _GEN_1893 : _GEN_2661; // @[executor.scala 466:52]
  wire [7:0] _GEN_2920 = opcode_2 == 4'hf ? _GEN_1894 : _GEN_2662; // @[executor.scala 466:52]
  wire [7:0] _GEN_2921 = opcode_2 == 4'hf ? _GEN_1895 : _GEN_2663; // @[executor.scala 466:52]
  wire [7:0] _GEN_2922 = opcode_2 == 4'hf ? _GEN_1896 : _GEN_2664; // @[executor.scala 466:52]
  wire [7:0] _GEN_2923 = opcode_2 == 4'hf ? _GEN_1897 : _GEN_2665; // @[executor.scala 466:52]
  wire [7:0] _GEN_2924 = opcode_2 == 4'hf ? _GEN_1898 : _GEN_2666; // @[executor.scala 466:52]
  wire [7:0] _GEN_2925 = opcode_2 == 4'hf ? _GEN_1899 : _GEN_2667; // @[executor.scala 466:52]
  wire [7:0] _GEN_2926 = opcode_2 == 4'hf ? _GEN_1900 : _GEN_2668; // @[executor.scala 466:52]
  wire [7:0] _GEN_2927 = opcode_2 == 4'hf ? _GEN_1901 : _GEN_2669; // @[executor.scala 466:52]
  wire [7:0] _GEN_2928 = opcode_2 == 4'hf ? _GEN_1902 : _GEN_2670; // @[executor.scala 466:52]
  wire [7:0] _GEN_2929 = opcode_2 == 4'hf ? _GEN_1903 : _GEN_2671; // @[executor.scala 466:52]
  wire [7:0] _GEN_2930 = opcode_2 == 4'hf ? _GEN_1904 : _GEN_2672; // @[executor.scala 466:52]
  wire [7:0] _GEN_2931 = opcode_2 == 4'hf ? _GEN_1905 : _GEN_2673; // @[executor.scala 466:52]
  wire [7:0] _GEN_2932 = opcode_2 == 4'hf ? _GEN_1906 : _GEN_2674; // @[executor.scala 466:52]
  wire [7:0] _GEN_2933 = opcode_2 == 4'hf ? _GEN_1907 : _GEN_2675; // @[executor.scala 466:52]
  wire [7:0] _GEN_2934 = opcode_2 == 4'hf ? _GEN_1908 : _GEN_2676; // @[executor.scala 466:52]
  wire [7:0] _GEN_2935 = opcode_2 == 4'hf ? _GEN_1909 : _GEN_2677; // @[executor.scala 466:52]
  wire [7:0] _GEN_2936 = opcode_2 == 4'hf ? _GEN_1910 : _GEN_2678; // @[executor.scala 466:52]
  wire [7:0] _GEN_2937 = opcode_2 == 4'hf ? _GEN_1911 : _GEN_2679; // @[executor.scala 466:52]
  wire [7:0] _GEN_2938 = opcode_2 == 4'hf ? _GEN_1912 : _GEN_2680; // @[executor.scala 466:52]
  wire [7:0] _GEN_2939 = opcode_2 == 4'hf ? _GEN_1913 : _GEN_2681; // @[executor.scala 466:52]
  wire [7:0] _GEN_2940 = opcode_2 == 4'hf ? _GEN_1914 : _GEN_2682; // @[executor.scala 466:52]
  wire [7:0] _GEN_2941 = opcode_2 == 4'hf ? _GEN_1915 : _GEN_2683; // @[executor.scala 466:52]
  wire [7:0] _GEN_2942 = opcode_2 == 4'hf ? _GEN_1916 : _GEN_2684; // @[executor.scala 466:52]
  wire [7:0] _GEN_2943 = opcode_2 == 4'hf ? _GEN_1917 : _GEN_2685; // @[executor.scala 466:52]
  wire [7:0] _GEN_2944 = opcode_2 == 4'hf ? _GEN_1918 : _GEN_2686; // @[executor.scala 466:52]
  wire [7:0] _GEN_2945 = opcode_2 == 4'hf ? _GEN_1919 : _GEN_2687; // @[executor.scala 466:52]
  wire [7:0] _GEN_2946 = opcode_2 == 4'hf ? _GEN_1920 : _GEN_2688; // @[executor.scala 466:52]
  wire [7:0] _GEN_2947 = opcode_2 == 4'hf ? _GEN_1921 : _GEN_2689; // @[executor.scala 466:52]
  wire [7:0] _GEN_2948 = opcode_2 == 4'hf ? _GEN_1922 : _GEN_2690; // @[executor.scala 466:52]
  wire [7:0] _GEN_2949 = opcode_2 == 4'hf ? _GEN_1923 : _GEN_2691; // @[executor.scala 466:52]
  wire [7:0] _GEN_2950 = opcode_2 == 4'hf ? _GEN_1924 : _GEN_2692; // @[executor.scala 466:52]
  wire [7:0] _GEN_2951 = opcode_2 == 4'hf ? _GEN_1925 : _GEN_2693; // @[executor.scala 466:52]
  wire [7:0] _GEN_2952 = opcode_2 == 4'hf ? _GEN_1926 : _GEN_2694; // @[executor.scala 466:52]
  wire [7:0] _GEN_2953 = opcode_2 == 4'hf ? _GEN_1927 : _GEN_2695; // @[executor.scala 466:52]
  wire [7:0] _GEN_2954 = opcode_2 == 4'hf ? _GEN_1928 : _GEN_2696; // @[executor.scala 466:52]
  wire [7:0] _GEN_2955 = opcode_2 == 4'hf ? _GEN_1929 : _GEN_2697; // @[executor.scala 466:52]
  wire [7:0] _GEN_2956 = opcode_2 == 4'hf ? _GEN_1930 : _GEN_2698; // @[executor.scala 466:52]
  wire [7:0] _GEN_2957 = opcode_2 == 4'hf ? _GEN_1931 : _GEN_2699; // @[executor.scala 466:52]
  wire [7:0] _GEN_2958 = opcode_2 == 4'hf ? _GEN_1932 : _GEN_2700; // @[executor.scala 466:52]
  wire [7:0] _GEN_2959 = opcode_2 == 4'hf ? _GEN_1933 : _GEN_2701; // @[executor.scala 466:52]
  wire [7:0] _GEN_2960 = opcode_2 == 4'hf ? _GEN_1934 : _GEN_2702; // @[executor.scala 466:52]
  wire [7:0] _GEN_2961 = opcode_2 == 4'hf ? _GEN_1935 : _GEN_2703; // @[executor.scala 466:52]
  wire [7:0] _GEN_2962 = opcode_2 == 4'hf ? _GEN_1936 : _GEN_2704; // @[executor.scala 466:52]
  wire [7:0] _GEN_2963 = opcode_2 == 4'hf ? _GEN_1937 : _GEN_2705; // @[executor.scala 466:52]
  wire [7:0] _GEN_2964 = opcode_2 == 4'hf ? _GEN_1938 : _GEN_2706; // @[executor.scala 466:52]
  wire [7:0] _GEN_2965 = opcode_2 == 4'hf ? _GEN_1939 : _GEN_2707; // @[executor.scala 466:52]
  wire [7:0] _GEN_2966 = opcode_2 == 4'hf ? _GEN_1940 : _GEN_2708; // @[executor.scala 466:52]
  wire [7:0] _GEN_2967 = opcode_2 == 4'hf ? _GEN_1941 : _GEN_2709; // @[executor.scala 466:52]
  wire [7:0] _GEN_2968 = opcode_2 == 4'hf ? _GEN_1942 : _GEN_2710; // @[executor.scala 466:52]
  wire [7:0] _GEN_2969 = opcode_2 == 4'hf ? _GEN_1943 : _GEN_2711; // @[executor.scala 466:52]
  wire [7:0] _GEN_2970 = opcode_2 == 4'hf ? _GEN_1944 : _GEN_2712; // @[executor.scala 466:52]
  wire [7:0] _GEN_2971 = opcode_2 == 4'hf ? _GEN_1945 : _GEN_2713; // @[executor.scala 466:52]
  wire [7:0] _GEN_2972 = opcode_2 == 4'hf ? _GEN_1946 : _GEN_2714; // @[executor.scala 466:52]
  wire [7:0] _GEN_2973 = opcode_2 == 4'hf ? _GEN_1947 : _GEN_2715; // @[executor.scala 466:52]
  wire [7:0] _GEN_2974 = opcode_2 == 4'hf ? _GEN_1948 : _GEN_2716; // @[executor.scala 466:52]
  wire [7:0] _GEN_2975 = opcode_2 == 4'hf ? _GEN_1949 : _GEN_2717; // @[executor.scala 466:52]
  wire [7:0] _GEN_2976 = opcode_2 == 4'hf ? _GEN_1950 : _GEN_2718; // @[executor.scala 466:52]
  wire [7:0] _GEN_2977 = opcode_2 == 4'hf ? _GEN_1951 : _GEN_2719; // @[executor.scala 466:52]
  wire [7:0] _GEN_2978 = opcode_2 == 4'hf ? _GEN_1952 : _GEN_2720; // @[executor.scala 466:52]
  wire [7:0] _GEN_2979 = opcode_2 == 4'hf ? _GEN_1953 : _GEN_2721; // @[executor.scala 466:52]
  wire [7:0] _GEN_2980 = opcode_2 == 4'hf ? _GEN_1954 : _GEN_2722; // @[executor.scala 466:52]
  wire [7:0] _GEN_2981 = opcode_2 == 4'hf ? _GEN_1955 : _GEN_2723; // @[executor.scala 466:52]
  wire [7:0] _GEN_2982 = opcode_2 == 4'hf ? _GEN_1956 : _GEN_2724; // @[executor.scala 466:52]
  wire [7:0] _GEN_2983 = opcode_2 == 4'hf ? _GEN_1957 : _GEN_2725; // @[executor.scala 466:52]
  wire [7:0] _GEN_2984 = opcode_2 == 4'hf ? _GEN_1958 : _GEN_2726; // @[executor.scala 466:52]
  wire [7:0] _GEN_2985 = opcode_2 == 4'hf ? _GEN_1959 : _GEN_2727; // @[executor.scala 466:52]
  wire [7:0] _GEN_2986 = opcode_2 == 4'hf ? _GEN_1960 : _GEN_2728; // @[executor.scala 466:52]
  wire [7:0] _GEN_2987 = opcode_2 == 4'hf ? _GEN_1961 : _GEN_2729; // @[executor.scala 466:52]
  wire [7:0] _GEN_2988 = opcode_2 == 4'hf ? _GEN_1962 : _GEN_2730; // @[executor.scala 466:52]
  wire [7:0] _GEN_2989 = opcode_2 == 4'hf ? _GEN_1963 : _GEN_2731; // @[executor.scala 466:52]
  wire [7:0] _GEN_2990 = opcode_2 == 4'hf ? _GEN_1964 : _GEN_2732; // @[executor.scala 466:52]
  wire [7:0] _GEN_2991 = opcode_2 == 4'hf ? _GEN_1965 : _GEN_2733; // @[executor.scala 466:52]
  wire [7:0] _GEN_2992 = opcode_2 == 4'hf ? _GEN_1966 : _GEN_2734; // @[executor.scala 466:52]
  wire [7:0] _GEN_2993 = opcode_2 == 4'hf ? _GEN_1967 : _GEN_2735; // @[executor.scala 466:52]
  wire [7:0] _GEN_2994 = opcode_2 == 4'hf ? _GEN_1968 : _GEN_2736; // @[executor.scala 466:52]
  wire [7:0] _GEN_2995 = opcode_2 == 4'hf ? _GEN_1969 : _GEN_2737; // @[executor.scala 466:52]
  wire [7:0] _GEN_2996 = opcode_2 == 4'hf ? _GEN_1970 : _GEN_2738; // @[executor.scala 466:52]
  wire [7:0] _GEN_2997 = opcode_2 == 4'hf ? _GEN_1971 : _GEN_2739; // @[executor.scala 466:52]
  wire [7:0] _GEN_2998 = opcode_2 == 4'hf ? _GEN_1972 : _GEN_2740; // @[executor.scala 466:52]
  wire [7:0] _GEN_2999 = opcode_2 == 4'hf ? _GEN_1973 : _GEN_2741; // @[executor.scala 466:52]
  wire [7:0] _GEN_3000 = opcode_2 == 4'hf ? _GEN_1974 : _GEN_2742; // @[executor.scala 466:52]
  wire [7:0] _GEN_3001 = opcode_2 == 4'hf ? _GEN_1975 : _GEN_2743; // @[executor.scala 466:52]
  wire [7:0] _GEN_3002 = opcode_2 == 4'hf ? _GEN_1976 : _GEN_2744; // @[executor.scala 466:52]
  wire [7:0] _GEN_3003 = opcode_2 == 4'hf ? _GEN_1977 : _GEN_2745; // @[executor.scala 466:52]
  wire [7:0] _GEN_3004 = opcode_2 == 4'hf ? _GEN_1978 : _GEN_2746; // @[executor.scala 466:52]
  wire [7:0] _GEN_3005 = opcode_2 == 4'hf ? _GEN_1979 : _GEN_2747; // @[executor.scala 466:52]
  wire [7:0] _GEN_3006 = opcode_2 == 4'hf ? _GEN_1980 : _GEN_2748; // @[executor.scala 466:52]
  wire [7:0] _GEN_3007 = opcode_2 == 4'hf ? _GEN_1981 : _GEN_2749; // @[executor.scala 466:52]
  wire [7:0] _GEN_3008 = opcode_2 == 4'hf ? _GEN_1982 : _GEN_2750; // @[executor.scala 466:52]
  wire [7:0] _GEN_3009 = opcode_2 == 4'hf ? _GEN_1983 : _GEN_2751; // @[executor.scala 466:52]
  wire [7:0] _GEN_3010 = opcode_2 == 4'hf ? _GEN_1984 : _GEN_2752; // @[executor.scala 466:52]
  wire [7:0] _GEN_3011 = opcode_2 == 4'hf ? _GEN_1985 : _GEN_2753; // @[executor.scala 466:52]
  wire [7:0] _GEN_3012 = opcode_2 == 4'hf ? _GEN_1986 : _GEN_2754; // @[executor.scala 466:52]
  wire [7:0] _GEN_3013 = opcode_2 == 4'hf ? _GEN_1987 : _GEN_2755; // @[executor.scala 466:52]
  wire [7:0] _GEN_3014 = opcode_2 == 4'hf ? _GEN_1988 : _GEN_2756; // @[executor.scala 466:52]
  wire [7:0] _GEN_3015 = opcode_2 == 4'hf ? _GEN_1989 : _GEN_2757; // @[executor.scala 466:52]
  wire [7:0] _GEN_3016 = opcode_2 == 4'hf ? _GEN_1990 : _GEN_2758; // @[executor.scala 466:52]
  wire [7:0] _GEN_3017 = opcode_2 == 4'hf ? _GEN_1991 : _GEN_2759; // @[executor.scala 466:52]
  wire [7:0] _GEN_3018 = opcode_2 == 4'hf ? _GEN_1992 : _GEN_2760; // @[executor.scala 466:52]
  wire [7:0] _GEN_3019 = opcode_2 == 4'hf ? _GEN_1993 : _GEN_2761; // @[executor.scala 466:52]
  wire [7:0] _GEN_3020 = opcode_2 == 4'hf ? _GEN_1994 : _GEN_2762; // @[executor.scala 466:52]
  wire [7:0] _GEN_3021 = opcode_2 == 4'hf ? _GEN_1995 : _GEN_2763; // @[executor.scala 466:52]
  wire [7:0] _GEN_3022 = opcode_2 == 4'hf ? _GEN_1996 : _GEN_2764; // @[executor.scala 466:52]
  wire [7:0] _GEN_3023 = opcode_2 == 4'hf ? _GEN_1997 : _GEN_2765; // @[executor.scala 466:52]
  wire [7:0] _GEN_3024 = opcode_2 == 4'hf ? _GEN_1998 : _GEN_2766; // @[executor.scala 466:52]
  wire [7:0] _GEN_3025 = opcode_2 == 4'hf ? _GEN_1999 : _GEN_2767; // @[executor.scala 466:52]
  wire [7:0] _GEN_3026 = opcode_2 == 4'hf ? _GEN_2000 : _GEN_2768; // @[executor.scala 466:52]
  wire [7:0] _GEN_3027 = opcode_2 == 4'hf ? _GEN_2001 : _GEN_2769; // @[executor.scala 466:52]
  wire [7:0] _GEN_3028 = opcode_2 == 4'hf ? _GEN_2002 : _GEN_2770; // @[executor.scala 466:52]
  wire [7:0] _GEN_3029 = opcode_2 == 4'hf ? _GEN_2003 : _GEN_2771; // @[executor.scala 466:52]
  wire [7:0] _GEN_3030 = opcode_2 == 4'hf ? _GEN_2004 : _GEN_2772; // @[executor.scala 466:52]
  wire [7:0] _GEN_3031 = opcode_2 == 4'hf ? _GEN_2005 : _GEN_2773; // @[executor.scala 466:52]
  wire [7:0] _GEN_3032 = opcode_2 == 4'hf ? _GEN_2006 : _GEN_2774; // @[executor.scala 466:52]
  wire [7:0] _GEN_3033 = opcode_2 == 4'hf ? _GEN_2007 : _GEN_2775; // @[executor.scala 466:52]
  wire [7:0] _GEN_3034 = opcode_2 == 4'hf ? _GEN_2008 : _GEN_2776; // @[executor.scala 466:52]
  wire [7:0] _GEN_3035 = opcode_2 == 4'hf ? _GEN_2009 : _GEN_2777; // @[executor.scala 466:52]
  wire [7:0] _GEN_3036 = opcode_2 == 4'hf ? _GEN_2010 : _GEN_2778; // @[executor.scala 466:52]
  wire [7:0] _GEN_3037 = opcode_2 == 4'hf ? _GEN_2011 : _GEN_2779; // @[executor.scala 466:52]
  wire [7:0] _GEN_3038 = opcode_2 == 4'hf ? _GEN_2012 : _GEN_2780; // @[executor.scala 466:52]
  wire [7:0] _GEN_3039 = opcode_2 == 4'hf ? _GEN_2013 : _GEN_2781; // @[executor.scala 466:52]
  wire [7:0] _GEN_3040 = opcode_2 == 4'hf ? _GEN_2014 : _GEN_2782; // @[executor.scala 466:52]
  wire [7:0] _GEN_3041 = opcode_2 == 4'hf ? _GEN_2015 : _GEN_2783; // @[executor.scala 466:52]
  wire [7:0] _GEN_3042 = opcode_2 == 4'hf ? _GEN_2016 : _GEN_2784; // @[executor.scala 466:52]
  wire [7:0] _GEN_3043 = opcode_2 == 4'hf ? _GEN_2017 : _GEN_2785; // @[executor.scala 466:52]
  wire [7:0] _GEN_3044 = opcode_2 == 4'hf ? _GEN_2018 : _GEN_2786; // @[executor.scala 466:52]
  wire [7:0] _GEN_3045 = opcode_2 == 4'hf ? _GEN_2019 : _GEN_2787; // @[executor.scala 466:52]
  wire [7:0] _GEN_3046 = opcode_2 == 4'hf ? _GEN_2020 : _GEN_2788; // @[executor.scala 466:52]
  wire [7:0] _GEN_3047 = opcode_2 == 4'hf ? _GEN_2021 : _GEN_2789; // @[executor.scala 466:52]
  wire [7:0] _GEN_3048 = opcode_2 == 4'hf ? _GEN_2022 : _GEN_2790; // @[executor.scala 466:52]
  wire [7:0] _GEN_3049 = opcode_2 == 4'hf ? _GEN_2023 : _GEN_2791; // @[executor.scala 466:52]
  wire [7:0] _GEN_3050 = opcode_2 == 4'hf ? _GEN_2024 : _GEN_2792; // @[executor.scala 466:52]
  wire [7:0] _GEN_3051 = opcode_2 == 4'hf ? _GEN_2025 : _GEN_2793; // @[executor.scala 466:52]
  wire [7:0] _GEN_3052 = opcode_2 == 4'hf ? _GEN_2026 : _GEN_2794; // @[executor.scala 466:52]
  wire [7:0] _GEN_3053 = opcode_2 == 4'hf ? _GEN_2027 : _GEN_2795; // @[executor.scala 466:52]
  wire [7:0] _GEN_3054 = opcode_2 == 4'hf ? _GEN_2028 : _GEN_2796; // @[executor.scala 466:52]
  wire [7:0] _GEN_3055 = opcode_2 == 4'hf ? _GEN_2029 : _GEN_2797; // @[executor.scala 466:52]
  wire [7:0] _GEN_3056 = opcode_2 == 4'hf ? _GEN_2030 : _GEN_2798; // @[executor.scala 466:52]
  wire [7:0] _GEN_3057 = opcode_2 == 4'hf ? _GEN_2031 : _GEN_2799; // @[executor.scala 466:52]
  wire [7:0] _GEN_3058 = opcode_2 == 4'hf ? _GEN_2032 : _GEN_2800; // @[executor.scala 466:52]
  wire [7:0] _GEN_3059 = opcode_2 == 4'hf ? _GEN_2033 : _GEN_2801; // @[executor.scala 466:52]
  wire [7:0] _GEN_3060 = opcode_2 == 4'hf ? _GEN_2034 : _GEN_2802; // @[executor.scala 466:52]
  wire [7:0] _GEN_3061 = opcode_2 == 4'hf ? _GEN_2035 : _GEN_2803; // @[executor.scala 466:52]
  wire [7:0] _GEN_3062 = opcode_2 == 4'hf ? _GEN_2036 : _GEN_2804; // @[executor.scala 466:52]
  wire [7:0] _GEN_3063 = opcode_2 == 4'hf ? _GEN_2037 : _GEN_2805; // @[executor.scala 466:52]
  wire [7:0] _GEN_3064 = opcode_2 == 4'hf ? _GEN_2038 : _GEN_2806; // @[executor.scala 466:52]
  wire [7:0] _GEN_3065 = opcode_2 == 4'hf ? _GEN_2039 : _GEN_2807; // @[executor.scala 466:52]
  wire [7:0] _GEN_3066 = opcode_2 == 4'hf ? _GEN_2040 : _GEN_2808; // @[executor.scala 466:52]
  wire [7:0] _GEN_3067 = opcode_2 == 4'hf ? _GEN_2041 : _GEN_2809; // @[executor.scala 466:52]
  wire [7:0] _GEN_3068 = opcode_2 == 4'hf ? _GEN_2042 : _GEN_2810; // @[executor.scala 466:52]
  wire [7:0] _GEN_3069 = opcode_2 == 4'hf ? _GEN_2043 : _GEN_2811; // @[executor.scala 466:52]
  wire [7:0] _GEN_3070 = opcode_2 == 4'hf ? _GEN_2044 : _GEN_2812; // @[executor.scala 466:52]
  wire [7:0] _GEN_3071 = opcode_2 == 4'hf ? _GEN_2045 : _GEN_2813; // @[executor.scala 466:52]
  wire [7:0] _GEN_3072 = opcode_2 == 4'hf ? _GEN_2046 : _GEN_2814; // @[executor.scala 466:52]
  wire [7:0] _GEN_3073 = opcode_2 == 4'hf ? _GEN_2047 : _GEN_2815; // @[executor.scala 466:52]
  wire [7:0] _GEN_3074 = opcode_2 == 4'hf ? _GEN_2048 : _GEN_2816; // @[executor.scala 466:52]
  wire [7:0] _GEN_3075 = opcode_2 == 4'hf ? _GEN_2049 : _GEN_2817; // @[executor.scala 466:52]
  wire [7:0] _GEN_3076 = opcode_2 == 4'hf ? _GEN_2050 : _GEN_2818; // @[executor.scala 466:52]
  wire [7:0] _GEN_3077 = opcode_2 == 4'hf ? _GEN_2051 : _GEN_2819; // @[executor.scala 466:52]
  wire [3:0] opcode_3 = vliw_3[31:28]; // @[primitive.scala 9:44]
  wire [7:0] _GEN_4554 = {{2'd0}, dst_offset_3}; // @[executor.scala 473:49]
  wire [7:0] byte_768 = field_3[7:0]; // @[executor.scala 475:56]
  wire [7:0] _GEN_3078 = mask_3[0] ? byte_768 : _GEN_2822; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] byte_769 = field_3[15:8]; // @[executor.scala 475:56]
  wire [7:0] _GEN_3079 = mask_3[1] ? byte_769 : _GEN_2823; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] byte_770 = field_3[23:16]; // @[executor.scala 475:56]
  wire [7:0] _GEN_3080 = mask_3[2] ? byte_770 : _GEN_2824; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] byte_771 = field_3[31:24]; // @[executor.scala 475:56]
  wire [7:0] _GEN_3081 = mask_3[3] ? byte_771 : _GEN_2825; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3082 = _GEN_4554 == 8'h0 ? _GEN_3078 : _GEN_2822; // @[executor.scala 473:84]
  wire [7:0] _GEN_3083 = _GEN_4554 == 8'h0 ? _GEN_3079 : _GEN_2823; // @[executor.scala 473:84]
  wire [7:0] _GEN_3084 = _GEN_4554 == 8'h0 ? _GEN_3080 : _GEN_2824; // @[executor.scala 473:84]
  wire [7:0] _GEN_3085 = _GEN_4554 == 8'h0 ? _GEN_3081 : _GEN_2825; // @[executor.scala 473:84]
  wire [7:0] _GEN_3086 = mask_3[0] ? byte_768 : _GEN_2826; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3087 = mask_3[1] ? byte_769 : _GEN_2827; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3088 = mask_3[2] ? byte_770 : _GEN_2828; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3089 = mask_3[3] ? byte_771 : _GEN_2829; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3090 = _GEN_4554 == 8'h1 ? _GEN_3086 : _GEN_2826; // @[executor.scala 473:84]
  wire [7:0] _GEN_3091 = _GEN_4554 == 8'h1 ? _GEN_3087 : _GEN_2827; // @[executor.scala 473:84]
  wire [7:0] _GEN_3092 = _GEN_4554 == 8'h1 ? _GEN_3088 : _GEN_2828; // @[executor.scala 473:84]
  wire [7:0] _GEN_3093 = _GEN_4554 == 8'h1 ? _GEN_3089 : _GEN_2829; // @[executor.scala 473:84]
  wire [7:0] _GEN_3094 = mask_3[0] ? byte_768 : _GEN_2830; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3095 = mask_3[1] ? byte_769 : _GEN_2831; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3096 = mask_3[2] ? byte_770 : _GEN_2832; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3097 = mask_3[3] ? byte_771 : _GEN_2833; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3098 = _GEN_4554 == 8'h2 ? _GEN_3094 : _GEN_2830; // @[executor.scala 473:84]
  wire [7:0] _GEN_3099 = _GEN_4554 == 8'h2 ? _GEN_3095 : _GEN_2831; // @[executor.scala 473:84]
  wire [7:0] _GEN_3100 = _GEN_4554 == 8'h2 ? _GEN_3096 : _GEN_2832; // @[executor.scala 473:84]
  wire [7:0] _GEN_3101 = _GEN_4554 == 8'h2 ? _GEN_3097 : _GEN_2833; // @[executor.scala 473:84]
  wire [7:0] _GEN_3102 = mask_3[0] ? byte_768 : _GEN_2834; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3103 = mask_3[1] ? byte_769 : _GEN_2835; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3104 = mask_3[2] ? byte_770 : _GEN_2836; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3105 = mask_3[3] ? byte_771 : _GEN_2837; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3106 = _GEN_4554 == 8'h3 ? _GEN_3102 : _GEN_2834; // @[executor.scala 473:84]
  wire [7:0] _GEN_3107 = _GEN_4554 == 8'h3 ? _GEN_3103 : _GEN_2835; // @[executor.scala 473:84]
  wire [7:0] _GEN_3108 = _GEN_4554 == 8'h3 ? _GEN_3104 : _GEN_2836; // @[executor.scala 473:84]
  wire [7:0] _GEN_3109 = _GEN_4554 == 8'h3 ? _GEN_3105 : _GEN_2837; // @[executor.scala 473:84]
  wire [7:0] _GEN_3110 = mask_3[0] ? byte_768 : _GEN_2838; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3111 = mask_3[1] ? byte_769 : _GEN_2839; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3112 = mask_3[2] ? byte_770 : _GEN_2840; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3113 = mask_3[3] ? byte_771 : _GEN_2841; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3114 = _GEN_4554 == 8'h4 ? _GEN_3110 : _GEN_2838; // @[executor.scala 473:84]
  wire [7:0] _GEN_3115 = _GEN_4554 == 8'h4 ? _GEN_3111 : _GEN_2839; // @[executor.scala 473:84]
  wire [7:0] _GEN_3116 = _GEN_4554 == 8'h4 ? _GEN_3112 : _GEN_2840; // @[executor.scala 473:84]
  wire [7:0] _GEN_3117 = _GEN_4554 == 8'h4 ? _GEN_3113 : _GEN_2841; // @[executor.scala 473:84]
  wire [7:0] _GEN_3118 = mask_3[0] ? byte_768 : _GEN_2842; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3119 = mask_3[1] ? byte_769 : _GEN_2843; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3120 = mask_3[2] ? byte_770 : _GEN_2844; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3121 = mask_3[3] ? byte_771 : _GEN_2845; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3122 = _GEN_4554 == 8'h5 ? _GEN_3118 : _GEN_2842; // @[executor.scala 473:84]
  wire [7:0] _GEN_3123 = _GEN_4554 == 8'h5 ? _GEN_3119 : _GEN_2843; // @[executor.scala 473:84]
  wire [7:0] _GEN_3124 = _GEN_4554 == 8'h5 ? _GEN_3120 : _GEN_2844; // @[executor.scala 473:84]
  wire [7:0] _GEN_3125 = _GEN_4554 == 8'h5 ? _GEN_3121 : _GEN_2845; // @[executor.scala 473:84]
  wire [7:0] _GEN_3126 = mask_3[0] ? byte_768 : _GEN_2846; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3127 = mask_3[1] ? byte_769 : _GEN_2847; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3128 = mask_3[2] ? byte_770 : _GEN_2848; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3129 = mask_3[3] ? byte_771 : _GEN_2849; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3130 = _GEN_4554 == 8'h6 ? _GEN_3126 : _GEN_2846; // @[executor.scala 473:84]
  wire [7:0] _GEN_3131 = _GEN_4554 == 8'h6 ? _GEN_3127 : _GEN_2847; // @[executor.scala 473:84]
  wire [7:0] _GEN_3132 = _GEN_4554 == 8'h6 ? _GEN_3128 : _GEN_2848; // @[executor.scala 473:84]
  wire [7:0] _GEN_3133 = _GEN_4554 == 8'h6 ? _GEN_3129 : _GEN_2849; // @[executor.scala 473:84]
  wire [7:0] _GEN_3134 = mask_3[0] ? byte_768 : _GEN_2850; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3135 = mask_3[1] ? byte_769 : _GEN_2851; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3136 = mask_3[2] ? byte_770 : _GEN_2852; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3137 = mask_3[3] ? byte_771 : _GEN_2853; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3138 = _GEN_4554 == 8'h7 ? _GEN_3134 : _GEN_2850; // @[executor.scala 473:84]
  wire [7:0] _GEN_3139 = _GEN_4554 == 8'h7 ? _GEN_3135 : _GEN_2851; // @[executor.scala 473:84]
  wire [7:0] _GEN_3140 = _GEN_4554 == 8'h7 ? _GEN_3136 : _GEN_2852; // @[executor.scala 473:84]
  wire [7:0] _GEN_3141 = _GEN_4554 == 8'h7 ? _GEN_3137 : _GEN_2853; // @[executor.scala 473:84]
  wire [7:0] _GEN_3142 = mask_3[0] ? byte_768 : _GEN_2854; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3143 = mask_3[1] ? byte_769 : _GEN_2855; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3144 = mask_3[2] ? byte_770 : _GEN_2856; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3145 = mask_3[3] ? byte_771 : _GEN_2857; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3146 = _GEN_4554 == 8'h8 ? _GEN_3142 : _GEN_2854; // @[executor.scala 473:84]
  wire [7:0] _GEN_3147 = _GEN_4554 == 8'h8 ? _GEN_3143 : _GEN_2855; // @[executor.scala 473:84]
  wire [7:0] _GEN_3148 = _GEN_4554 == 8'h8 ? _GEN_3144 : _GEN_2856; // @[executor.scala 473:84]
  wire [7:0] _GEN_3149 = _GEN_4554 == 8'h8 ? _GEN_3145 : _GEN_2857; // @[executor.scala 473:84]
  wire [7:0] _GEN_3150 = mask_3[0] ? byte_768 : _GEN_2858; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3151 = mask_3[1] ? byte_769 : _GEN_2859; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3152 = mask_3[2] ? byte_770 : _GEN_2860; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3153 = mask_3[3] ? byte_771 : _GEN_2861; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3154 = _GEN_4554 == 8'h9 ? _GEN_3150 : _GEN_2858; // @[executor.scala 473:84]
  wire [7:0] _GEN_3155 = _GEN_4554 == 8'h9 ? _GEN_3151 : _GEN_2859; // @[executor.scala 473:84]
  wire [7:0] _GEN_3156 = _GEN_4554 == 8'h9 ? _GEN_3152 : _GEN_2860; // @[executor.scala 473:84]
  wire [7:0] _GEN_3157 = _GEN_4554 == 8'h9 ? _GEN_3153 : _GEN_2861; // @[executor.scala 473:84]
  wire [7:0] _GEN_3158 = mask_3[0] ? byte_768 : _GEN_2862; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3159 = mask_3[1] ? byte_769 : _GEN_2863; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3160 = mask_3[2] ? byte_770 : _GEN_2864; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3161 = mask_3[3] ? byte_771 : _GEN_2865; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3162 = _GEN_4554 == 8'ha ? _GEN_3158 : _GEN_2862; // @[executor.scala 473:84]
  wire [7:0] _GEN_3163 = _GEN_4554 == 8'ha ? _GEN_3159 : _GEN_2863; // @[executor.scala 473:84]
  wire [7:0] _GEN_3164 = _GEN_4554 == 8'ha ? _GEN_3160 : _GEN_2864; // @[executor.scala 473:84]
  wire [7:0] _GEN_3165 = _GEN_4554 == 8'ha ? _GEN_3161 : _GEN_2865; // @[executor.scala 473:84]
  wire [7:0] _GEN_3166 = mask_3[0] ? byte_768 : _GEN_2866; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3167 = mask_3[1] ? byte_769 : _GEN_2867; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3168 = mask_3[2] ? byte_770 : _GEN_2868; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3169 = mask_3[3] ? byte_771 : _GEN_2869; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3170 = _GEN_4554 == 8'hb ? _GEN_3166 : _GEN_2866; // @[executor.scala 473:84]
  wire [7:0] _GEN_3171 = _GEN_4554 == 8'hb ? _GEN_3167 : _GEN_2867; // @[executor.scala 473:84]
  wire [7:0] _GEN_3172 = _GEN_4554 == 8'hb ? _GEN_3168 : _GEN_2868; // @[executor.scala 473:84]
  wire [7:0] _GEN_3173 = _GEN_4554 == 8'hb ? _GEN_3169 : _GEN_2869; // @[executor.scala 473:84]
  wire [7:0] _GEN_3174 = mask_3[0] ? byte_768 : _GEN_2870; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3175 = mask_3[1] ? byte_769 : _GEN_2871; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3176 = mask_3[2] ? byte_770 : _GEN_2872; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3177 = mask_3[3] ? byte_771 : _GEN_2873; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3178 = _GEN_4554 == 8'hc ? _GEN_3174 : _GEN_2870; // @[executor.scala 473:84]
  wire [7:0] _GEN_3179 = _GEN_4554 == 8'hc ? _GEN_3175 : _GEN_2871; // @[executor.scala 473:84]
  wire [7:0] _GEN_3180 = _GEN_4554 == 8'hc ? _GEN_3176 : _GEN_2872; // @[executor.scala 473:84]
  wire [7:0] _GEN_3181 = _GEN_4554 == 8'hc ? _GEN_3177 : _GEN_2873; // @[executor.scala 473:84]
  wire [7:0] _GEN_3182 = mask_3[0] ? byte_768 : _GEN_2874; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3183 = mask_3[1] ? byte_769 : _GEN_2875; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3184 = mask_3[2] ? byte_770 : _GEN_2876; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3185 = mask_3[3] ? byte_771 : _GEN_2877; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3186 = _GEN_4554 == 8'hd ? _GEN_3182 : _GEN_2874; // @[executor.scala 473:84]
  wire [7:0] _GEN_3187 = _GEN_4554 == 8'hd ? _GEN_3183 : _GEN_2875; // @[executor.scala 473:84]
  wire [7:0] _GEN_3188 = _GEN_4554 == 8'hd ? _GEN_3184 : _GEN_2876; // @[executor.scala 473:84]
  wire [7:0] _GEN_3189 = _GEN_4554 == 8'hd ? _GEN_3185 : _GEN_2877; // @[executor.scala 473:84]
  wire [7:0] _GEN_3190 = mask_3[0] ? byte_768 : _GEN_2878; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3191 = mask_3[1] ? byte_769 : _GEN_2879; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3192 = mask_3[2] ? byte_770 : _GEN_2880; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3193 = mask_3[3] ? byte_771 : _GEN_2881; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3194 = _GEN_4554 == 8'he ? _GEN_3190 : _GEN_2878; // @[executor.scala 473:84]
  wire [7:0] _GEN_3195 = _GEN_4554 == 8'he ? _GEN_3191 : _GEN_2879; // @[executor.scala 473:84]
  wire [7:0] _GEN_3196 = _GEN_4554 == 8'he ? _GEN_3192 : _GEN_2880; // @[executor.scala 473:84]
  wire [7:0] _GEN_3197 = _GEN_4554 == 8'he ? _GEN_3193 : _GEN_2881; // @[executor.scala 473:84]
  wire [7:0] _GEN_3198 = mask_3[0] ? byte_768 : _GEN_2882; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3199 = mask_3[1] ? byte_769 : _GEN_2883; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3200 = mask_3[2] ? byte_770 : _GEN_2884; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3201 = mask_3[3] ? byte_771 : _GEN_2885; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3202 = _GEN_4554 == 8'hf ? _GEN_3198 : _GEN_2882; // @[executor.scala 473:84]
  wire [7:0] _GEN_3203 = _GEN_4554 == 8'hf ? _GEN_3199 : _GEN_2883; // @[executor.scala 473:84]
  wire [7:0] _GEN_3204 = _GEN_4554 == 8'hf ? _GEN_3200 : _GEN_2884; // @[executor.scala 473:84]
  wire [7:0] _GEN_3205 = _GEN_4554 == 8'hf ? _GEN_3201 : _GEN_2885; // @[executor.scala 473:84]
  wire [7:0] _GEN_3206 = mask_3[0] ? byte_768 : _GEN_2886; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3207 = mask_3[1] ? byte_769 : _GEN_2887; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3208 = mask_3[2] ? byte_770 : _GEN_2888; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3209 = mask_3[3] ? byte_771 : _GEN_2889; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3210 = _GEN_4554 == 8'h10 ? _GEN_3206 : _GEN_2886; // @[executor.scala 473:84]
  wire [7:0] _GEN_3211 = _GEN_4554 == 8'h10 ? _GEN_3207 : _GEN_2887; // @[executor.scala 473:84]
  wire [7:0] _GEN_3212 = _GEN_4554 == 8'h10 ? _GEN_3208 : _GEN_2888; // @[executor.scala 473:84]
  wire [7:0] _GEN_3213 = _GEN_4554 == 8'h10 ? _GEN_3209 : _GEN_2889; // @[executor.scala 473:84]
  wire [7:0] _GEN_3214 = mask_3[0] ? byte_768 : _GEN_2890; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3215 = mask_3[1] ? byte_769 : _GEN_2891; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3216 = mask_3[2] ? byte_770 : _GEN_2892; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3217 = mask_3[3] ? byte_771 : _GEN_2893; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3218 = _GEN_4554 == 8'h11 ? _GEN_3214 : _GEN_2890; // @[executor.scala 473:84]
  wire [7:0] _GEN_3219 = _GEN_4554 == 8'h11 ? _GEN_3215 : _GEN_2891; // @[executor.scala 473:84]
  wire [7:0] _GEN_3220 = _GEN_4554 == 8'h11 ? _GEN_3216 : _GEN_2892; // @[executor.scala 473:84]
  wire [7:0] _GEN_3221 = _GEN_4554 == 8'h11 ? _GEN_3217 : _GEN_2893; // @[executor.scala 473:84]
  wire [7:0] _GEN_3222 = mask_3[0] ? byte_768 : _GEN_2894; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3223 = mask_3[1] ? byte_769 : _GEN_2895; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3224 = mask_3[2] ? byte_770 : _GEN_2896; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3225 = mask_3[3] ? byte_771 : _GEN_2897; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3226 = _GEN_4554 == 8'h12 ? _GEN_3222 : _GEN_2894; // @[executor.scala 473:84]
  wire [7:0] _GEN_3227 = _GEN_4554 == 8'h12 ? _GEN_3223 : _GEN_2895; // @[executor.scala 473:84]
  wire [7:0] _GEN_3228 = _GEN_4554 == 8'h12 ? _GEN_3224 : _GEN_2896; // @[executor.scala 473:84]
  wire [7:0] _GEN_3229 = _GEN_4554 == 8'h12 ? _GEN_3225 : _GEN_2897; // @[executor.scala 473:84]
  wire [7:0] _GEN_3230 = mask_3[0] ? byte_768 : _GEN_2898; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3231 = mask_3[1] ? byte_769 : _GEN_2899; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3232 = mask_3[2] ? byte_770 : _GEN_2900; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3233 = mask_3[3] ? byte_771 : _GEN_2901; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3234 = _GEN_4554 == 8'h13 ? _GEN_3230 : _GEN_2898; // @[executor.scala 473:84]
  wire [7:0] _GEN_3235 = _GEN_4554 == 8'h13 ? _GEN_3231 : _GEN_2899; // @[executor.scala 473:84]
  wire [7:0] _GEN_3236 = _GEN_4554 == 8'h13 ? _GEN_3232 : _GEN_2900; // @[executor.scala 473:84]
  wire [7:0] _GEN_3237 = _GEN_4554 == 8'h13 ? _GEN_3233 : _GEN_2901; // @[executor.scala 473:84]
  wire [7:0] _GEN_3238 = mask_3[0] ? byte_768 : _GEN_2902; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3239 = mask_3[1] ? byte_769 : _GEN_2903; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3240 = mask_3[2] ? byte_770 : _GEN_2904; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3241 = mask_3[3] ? byte_771 : _GEN_2905; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3242 = _GEN_4554 == 8'h14 ? _GEN_3238 : _GEN_2902; // @[executor.scala 473:84]
  wire [7:0] _GEN_3243 = _GEN_4554 == 8'h14 ? _GEN_3239 : _GEN_2903; // @[executor.scala 473:84]
  wire [7:0] _GEN_3244 = _GEN_4554 == 8'h14 ? _GEN_3240 : _GEN_2904; // @[executor.scala 473:84]
  wire [7:0] _GEN_3245 = _GEN_4554 == 8'h14 ? _GEN_3241 : _GEN_2905; // @[executor.scala 473:84]
  wire [7:0] _GEN_3246 = mask_3[0] ? byte_768 : _GEN_2906; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3247 = mask_3[1] ? byte_769 : _GEN_2907; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3248 = mask_3[2] ? byte_770 : _GEN_2908; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3249 = mask_3[3] ? byte_771 : _GEN_2909; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3250 = _GEN_4554 == 8'h15 ? _GEN_3246 : _GEN_2906; // @[executor.scala 473:84]
  wire [7:0] _GEN_3251 = _GEN_4554 == 8'h15 ? _GEN_3247 : _GEN_2907; // @[executor.scala 473:84]
  wire [7:0] _GEN_3252 = _GEN_4554 == 8'h15 ? _GEN_3248 : _GEN_2908; // @[executor.scala 473:84]
  wire [7:0] _GEN_3253 = _GEN_4554 == 8'h15 ? _GEN_3249 : _GEN_2909; // @[executor.scala 473:84]
  wire [7:0] _GEN_3254 = mask_3[0] ? byte_768 : _GEN_2910; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3255 = mask_3[1] ? byte_769 : _GEN_2911; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3256 = mask_3[2] ? byte_770 : _GEN_2912; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3257 = mask_3[3] ? byte_771 : _GEN_2913; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3258 = _GEN_4554 == 8'h16 ? _GEN_3254 : _GEN_2910; // @[executor.scala 473:84]
  wire [7:0] _GEN_3259 = _GEN_4554 == 8'h16 ? _GEN_3255 : _GEN_2911; // @[executor.scala 473:84]
  wire [7:0] _GEN_3260 = _GEN_4554 == 8'h16 ? _GEN_3256 : _GEN_2912; // @[executor.scala 473:84]
  wire [7:0] _GEN_3261 = _GEN_4554 == 8'h16 ? _GEN_3257 : _GEN_2913; // @[executor.scala 473:84]
  wire [7:0] _GEN_3262 = mask_3[0] ? byte_768 : _GEN_2914; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3263 = mask_3[1] ? byte_769 : _GEN_2915; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3264 = mask_3[2] ? byte_770 : _GEN_2916; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3265 = mask_3[3] ? byte_771 : _GEN_2917; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3266 = _GEN_4554 == 8'h17 ? _GEN_3262 : _GEN_2914; // @[executor.scala 473:84]
  wire [7:0] _GEN_3267 = _GEN_4554 == 8'h17 ? _GEN_3263 : _GEN_2915; // @[executor.scala 473:84]
  wire [7:0] _GEN_3268 = _GEN_4554 == 8'h17 ? _GEN_3264 : _GEN_2916; // @[executor.scala 473:84]
  wire [7:0] _GEN_3269 = _GEN_4554 == 8'h17 ? _GEN_3265 : _GEN_2917; // @[executor.scala 473:84]
  wire [7:0] _GEN_3270 = mask_3[0] ? byte_768 : _GEN_2918; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3271 = mask_3[1] ? byte_769 : _GEN_2919; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3272 = mask_3[2] ? byte_770 : _GEN_2920; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3273 = mask_3[3] ? byte_771 : _GEN_2921; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3274 = _GEN_4554 == 8'h18 ? _GEN_3270 : _GEN_2918; // @[executor.scala 473:84]
  wire [7:0] _GEN_3275 = _GEN_4554 == 8'h18 ? _GEN_3271 : _GEN_2919; // @[executor.scala 473:84]
  wire [7:0] _GEN_3276 = _GEN_4554 == 8'h18 ? _GEN_3272 : _GEN_2920; // @[executor.scala 473:84]
  wire [7:0] _GEN_3277 = _GEN_4554 == 8'h18 ? _GEN_3273 : _GEN_2921; // @[executor.scala 473:84]
  wire [7:0] _GEN_3278 = mask_3[0] ? byte_768 : _GEN_2922; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3279 = mask_3[1] ? byte_769 : _GEN_2923; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3280 = mask_3[2] ? byte_770 : _GEN_2924; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3281 = mask_3[3] ? byte_771 : _GEN_2925; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3282 = _GEN_4554 == 8'h19 ? _GEN_3278 : _GEN_2922; // @[executor.scala 473:84]
  wire [7:0] _GEN_3283 = _GEN_4554 == 8'h19 ? _GEN_3279 : _GEN_2923; // @[executor.scala 473:84]
  wire [7:0] _GEN_3284 = _GEN_4554 == 8'h19 ? _GEN_3280 : _GEN_2924; // @[executor.scala 473:84]
  wire [7:0] _GEN_3285 = _GEN_4554 == 8'h19 ? _GEN_3281 : _GEN_2925; // @[executor.scala 473:84]
  wire [7:0] _GEN_3286 = mask_3[0] ? byte_768 : _GEN_2926; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3287 = mask_3[1] ? byte_769 : _GEN_2927; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3288 = mask_3[2] ? byte_770 : _GEN_2928; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3289 = mask_3[3] ? byte_771 : _GEN_2929; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3290 = _GEN_4554 == 8'h1a ? _GEN_3286 : _GEN_2926; // @[executor.scala 473:84]
  wire [7:0] _GEN_3291 = _GEN_4554 == 8'h1a ? _GEN_3287 : _GEN_2927; // @[executor.scala 473:84]
  wire [7:0] _GEN_3292 = _GEN_4554 == 8'h1a ? _GEN_3288 : _GEN_2928; // @[executor.scala 473:84]
  wire [7:0] _GEN_3293 = _GEN_4554 == 8'h1a ? _GEN_3289 : _GEN_2929; // @[executor.scala 473:84]
  wire [7:0] _GEN_3294 = mask_3[0] ? byte_768 : _GEN_2930; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3295 = mask_3[1] ? byte_769 : _GEN_2931; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3296 = mask_3[2] ? byte_770 : _GEN_2932; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3297 = mask_3[3] ? byte_771 : _GEN_2933; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3298 = _GEN_4554 == 8'h1b ? _GEN_3294 : _GEN_2930; // @[executor.scala 473:84]
  wire [7:0] _GEN_3299 = _GEN_4554 == 8'h1b ? _GEN_3295 : _GEN_2931; // @[executor.scala 473:84]
  wire [7:0] _GEN_3300 = _GEN_4554 == 8'h1b ? _GEN_3296 : _GEN_2932; // @[executor.scala 473:84]
  wire [7:0] _GEN_3301 = _GEN_4554 == 8'h1b ? _GEN_3297 : _GEN_2933; // @[executor.scala 473:84]
  wire [7:0] _GEN_3302 = mask_3[0] ? byte_768 : _GEN_2934; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3303 = mask_3[1] ? byte_769 : _GEN_2935; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3304 = mask_3[2] ? byte_770 : _GEN_2936; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3305 = mask_3[3] ? byte_771 : _GEN_2937; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3306 = _GEN_4554 == 8'h1c ? _GEN_3302 : _GEN_2934; // @[executor.scala 473:84]
  wire [7:0] _GEN_3307 = _GEN_4554 == 8'h1c ? _GEN_3303 : _GEN_2935; // @[executor.scala 473:84]
  wire [7:0] _GEN_3308 = _GEN_4554 == 8'h1c ? _GEN_3304 : _GEN_2936; // @[executor.scala 473:84]
  wire [7:0] _GEN_3309 = _GEN_4554 == 8'h1c ? _GEN_3305 : _GEN_2937; // @[executor.scala 473:84]
  wire [7:0] _GEN_3310 = mask_3[0] ? byte_768 : _GEN_2938; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3311 = mask_3[1] ? byte_769 : _GEN_2939; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3312 = mask_3[2] ? byte_770 : _GEN_2940; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3313 = mask_3[3] ? byte_771 : _GEN_2941; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3314 = _GEN_4554 == 8'h1d ? _GEN_3310 : _GEN_2938; // @[executor.scala 473:84]
  wire [7:0] _GEN_3315 = _GEN_4554 == 8'h1d ? _GEN_3311 : _GEN_2939; // @[executor.scala 473:84]
  wire [7:0] _GEN_3316 = _GEN_4554 == 8'h1d ? _GEN_3312 : _GEN_2940; // @[executor.scala 473:84]
  wire [7:0] _GEN_3317 = _GEN_4554 == 8'h1d ? _GEN_3313 : _GEN_2941; // @[executor.scala 473:84]
  wire [7:0] _GEN_3318 = mask_3[0] ? byte_768 : _GEN_2942; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3319 = mask_3[1] ? byte_769 : _GEN_2943; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3320 = mask_3[2] ? byte_770 : _GEN_2944; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3321 = mask_3[3] ? byte_771 : _GEN_2945; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3322 = _GEN_4554 == 8'h1e ? _GEN_3318 : _GEN_2942; // @[executor.scala 473:84]
  wire [7:0] _GEN_3323 = _GEN_4554 == 8'h1e ? _GEN_3319 : _GEN_2943; // @[executor.scala 473:84]
  wire [7:0] _GEN_3324 = _GEN_4554 == 8'h1e ? _GEN_3320 : _GEN_2944; // @[executor.scala 473:84]
  wire [7:0] _GEN_3325 = _GEN_4554 == 8'h1e ? _GEN_3321 : _GEN_2945; // @[executor.scala 473:84]
  wire [7:0] _GEN_3326 = mask_3[0] ? byte_768 : _GEN_2946; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3327 = mask_3[1] ? byte_769 : _GEN_2947; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3328 = mask_3[2] ? byte_770 : _GEN_2948; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3329 = mask_3[3] ? byte_771 : _GEN_2949; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3330 = _GEN_4554 == 8'h1f ? _GEN_3326 : _GEN_2946; // @[executor.scala 473:84]
  wire [7:0] _GEN_3331 = _GEN_4554 == 8'h1f ? _GEN_3327 : _GEN_2947; // @[executor.scala 473:84]
  wire [7:0] _GEN_3332 = _GEN_4554 == 8'h1f ? _GEN_3328 : _GEN_2948; // @[executor.scala 473:84]
  wire [7:0] _GEN_3333 = _GEN_4554 == 8'h1f ? _GEN_3329 : _GEN_2949; // @[executor.scala 473:84]
  wire [7:0] _GEN_3334 = mask_3[0] ? byte_768 : _GEN_2950; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3335 = mask_3[1] ? byte_769 : _GEN_2951; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3336 = mask_3[2] ? byte_770 : _GEN_2952; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3337 = mask_3[3] ? byte_771 : _GEN_2953; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3338 = _GEN_4554 == 8'h20 ? _GEN_3334 : _GEN_2950; // @[executor.scala 473:84]
  wire [7:0] _GEN_3339 = _GEN_4554 == 8'h20 ? _GEN_3335 : _GEN_2951; // @[executor.scala 473:84]
  wire [7:0] _GEN_3340 = _GEN_4554 == 8'h20 ? _GEN_3336 : _GEN_2952; // @[executor.scala 473:84]
  wire [7:0] _GEN_3341 = _GEN_4554 == 8'h20 ? _GEN_3337 : _GEN_2953; // @[executor.scala 473:84]
  wire [7:0] _GEN_3342 = mask_3[0] ? byte_768 : _GEN_2954; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3343 = mask_3[1] ? byte_769 : _GEN_2955; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3344 = mask_3[2] ? byte_770 : _GEN_2956; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3345 = mask_3[3] ? byte_771 : _GEN_2957; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3346 = _GEN_4554 == 8'h21 ? _GEN_3342 : _GEN_2954; // @[executor.scala 473:84]
  wire [7:0] _GEN_3347 = _GEN_4554 == 8'h21 ? _GEN_3343 : _GEN_2955; // @[executor.scala 473:84]
  wire [7:0] _GEN_3348 = _GEN_4554 == 8'h21 ? _GEN_3344 : _GEN_2956; // @[executor.scala 473:84]
  wire [7:0] _GEN_3349 = _GEN_4554 == 8'h21 ? _GEN_3345 : _GEN_2957; // @[executor.scala 473:84]
  wire [7:0] _GEN_3350 = mask_3[0] ? byte_768 : _GEN_2958; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3351 = mask_3[1] ? byte_769 : _GEN_2959; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3352 = mask_3[2] ? byte_770 : _GEN_2960; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3353 = mask_3[3] ? byte_771 : _GEN_2961; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3354 = _GEN_4554 == 8'h22 ? _GEN_3350 : _GEN_2958; // @[executor.scala 473:84]
  wire [7:0] _GEN_3355 = _GEN_4554 == 8'h22 ? _GEN_3351 : _GEN_2959; // @[executor.scala 473:84]
  wire [7:0] _GEN_3356 = _GEN_4554 == 8'h22 ? _GEN_3352 : _GEN_2960; // @[executor.scala 473:84]
  wire [7:0] _GEN_3357 = _GEN_4554 == 8'h22 ? _GEN_3353 : _GEN_2961; // @[executor.scala 473:84]
  wire [7:0] _GEN_3358 = mask_3[0] ? byte_768 : _GEN_2962; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3359 = mask_3[1] ? byte_769 : _GEN_2963; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3360 = mask_3[2] ? byte_770 : _GEN_2964; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3361 = mask_3[3] ? byte_771 : _GEN_2965; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3362 = _GEN_4554 == 8'h23 ? _GEN_3358 : _GEN_2962; // @[executor.scala 473:84]
  wire [7:0] _GEN_3363 = _GEN_4554 == 8'h23 ? _GEN_3359 : _GEN_2963; // @[executor.scala 473:84]
  wire [7:0] _GEN_3364 = _GEN_4554 == 8'h23 ? _GEN_3360 : _GEN_2964; // @[executor.scala 473:84]
  wire [7:0] _GEN_3365 = _GEN_4554 == 8'h23 ? _GEN_3361 : _GEN_2965; // @[executor.scala 473:84]
  wire [7:0] _GEN_3366 = mask_3[0] ? byte_768 : _GEN_2966; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3367 = mask_3[1] ? byte_769 : _GEN_2967; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3368 = mask_3[2] ? byte_770 : _GEN_2968; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3369 = mask_3[3] ? byte_771 : _GEN_2969; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3370 = _GEN_4554 == 8'h24 ? _GEN_3366 : _GEN_2966; // @[executor.scala 473:84]
  wire [7:0] _GEN_3371 = _GEN_4554 == 8'h24 ? _GEN_3367 : _GEN_2967; // @[executor.scala 473:84]
  wire [7:0] _GEN_3372 = _GEN_4554 == 8'h24 ? _GEN_3368 : _GEN_2968; // @[executor.scala 473:84]
  wire [7:0] _GEN_3373 = _GEN_4554 == 8'h24 ? _GEN_3369 : _GEN_2969; // @[executor.scala 473:84]
  wire [7:0] _GEN_3374 = mask_3[0] ? byte_768 : _GEN_2970; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3375 = mask_3[1] ? byte_769 : _GEN_2971; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3376 = mask_3[2] ? byte_770 : _GEN_2972; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3377 = mask_3[3] ? byte_771 : _GEN_2973; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3378 = _GEN_4554 == 8'h25 ? _GEN_3374 : _GEN_2970; // @[executor.scala 473:84]
  wire [7:0] _GEN_3379 = _GEN_4554 == 8'h25 ? _GEN_3375 : _GEN_2971; // @[executor.scala 473:84]
  wire [7:0] _GEN_3380 = _GEN_4554 == 8'h25 ? _GEN_3376 : _GEN_2972; // @[executor.scala 473:84]
  wire [7:0] _GEN_3381 = _GEN_4554 == 8'h25 ? _GEN_3377 : _GEN_2973; // @[executor.scala 473:84]
  wire [7:0] _GEN_3382 = mask_3[0] ? byte_768 : _GEN_2974; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3383 = mask_3[1] ? byte_769 : _GEN_2975; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3384 = mask_3[2] ? byte_770 : _GEN_2976; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3385 = mask_3[3] ? byte_771 : _GEN_2977; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3386 = _GEN_4554 == 8'h26 ? _GEN_3382 : _GEN_2974; // @[executor.scala 473:84]
  wire [7:0] _GEN_3387 = _GEN_4554 == 8'h26 ? _GEN_3383 : _GEN_2975; // @[executor.scala 473:84]
  wire [7:0] _GEN_3388 = _GEN_4554 == 8'h26 ? _GEN_3384 : _GEN_2976; // @[executor.scala 473:84]
  wire [7:0] _GEN_3389 = _GEN_4554 == 8'h26 ? _GEN_3385 : _GEN_2977; // @[executor.scala 473:84]
  wire [7:0] _GEN_3390 = mask_3[0] ? byte_768 : _GEN_2978; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3391 = mask_3[1] ? byte_769 : _GEN_2979; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3392 = mask_3[2] ? byte_770 : _GEN_2980; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3393 = mask_3[3] ? byte_771 : _GEN_2981; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3394 = _GEN_4554 == 8'h27 ? _GEN_3390 : _GEN_2978; // @[executor.scala 473:84]
  wire [7:0] _GEN_3395 = _GEN_4554 == 8'h27 ? _GEN_3391 : _GEN_2979; // @[executor.scala 473:84]
  wire [7:0] _GEN_3396 = _GEN_4554 == 8'h27 ? _GEN_3392 : _GEN_2980; // @[executor.scala 473:84]
  wire [7:0] _GEN_3397 = _GEN_4554 == 8'h27 ? _GEN_3393 : _GEN_2981; // @[executor.scala 473:84]
  wire [7:0] _GEN_3398 = mask_3[0] ? byte_768 : _GEN_2982; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3399 = mask_3[1] ? byte_769 : _GEN_2983; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3400 = mask_3[2] ? byte_770 : _GEN_2984; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3401 = mask_3[3] ? byte_771 : _GEN_2985; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3402 = _GEN_4554 == 8'h28 ? _GEN_3398 : _GEN_2982; // @[executor.scala 473:84]
  wire [7:0] _GEN_3403 = _GEN_4554 == 8'h28 ? _GEN_3399 : _GEN_2983; // @[executor.scala 473:84]
  wire [7:0] _GEN_3404 = _GEN_4554 == 8'h28 ? _GEN_3400 : _GEN_2984; // @[executor.scala 473:84]
  wire [7:0] _GEN_3405 = _GEN_4554 == 8'h28 ? _GEN_3401 : _GEN_2985; // @[executor.scala 473:84]
  wire [7:0] _GEN_3406 = mask_3[0] ? byte_768 : _GEN_2986; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3407 = mask_3[1] ? byte_769 : _GEN_2987; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3408 = mask_3[2] ? byte_770 : _GEN_2988; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3409 = mask_3[3] ? byte_771 : _GEN_2989; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3410 = _GEN_4554 == 8'h29 ? _GEN_3406 : _GEN_2986; // @[executor.scala 473:84]
  wire [7:0] _GEN_3411 = _GEN_4554 == 8'h29 ? _GEN_3407 : _GEN_2987; // @[executor.scala 473:84]
  wire [7:0] _GEN_3412 = _GEN_4554 == 8'h29 ? _GEN_3408 : _GEN_2988; // @[executor.scala 473:84]
  wire [7:0] _GEN_3413 = _GEN_4554 == 8'h29 ? _GEN_3409 : _GEN_2989; // @[executor.scala 473:84]
  wire [7:0] _GEN_3414 = mask_3[0] ? byte_768 : _GEN_2990; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3415 = mask_3[1] ? byte_769 : _GEN_2991; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3416 = mask_3[2] ? byte_770 : _GEN_2992; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3417 = mask_3[3] ? byte_771 : _GEN_2993; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3418 = _GEN_4554 == 8'h2a ? _GEN_3414 : _GEN_2990; // @[executor.scala 473:84]
  wire [7:0] _GEN_3419 = _GEN_4554 == 8'h2a ? _GEN_3415 : _GEN_2991; // @[executor.scala 473:84]
  wire [7:0] _GEN_3420 = _GEN_4554 == 8'h2a ? _GEN_3416 : _GEN_2992; // @[executor.scala 473:84]
  wire [7:0] _GEN_3421 = _GEN_4554 == 8'h2a ? _GEN_3417 : _GEN_2993; // @[executor.scala 473:84]
  wire [7:0] _GEN_3422 = mask_3[0] ? byte_768 : _GEN_2994; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3423 = mask_3[1] ? byte_769 : _GEN_2995; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3424 = mask_3[2] ? byte_770 : _GEN_2996; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3425 = mask_3[3] ? byte_771 : _GEN_2997; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3426 = _GEN_4554 == 8'h2b ? _GEN_3422 : _GEN_2994; // @[executor.scala 473:84]
  wire [7:0] _GEN_3427 = _GEN_4554 == 8'h2b ? _GEN_3423 : _GEN_2995; // @[executor.scala 473:84]
  wire [7:0] _GEN_3428 = _GEN_4554 == 8'h2b ? _GEN_3424 : _GEN_2996; // @[executor.scala 473:84]
  wire [7:0] _GEN_3429 = _GEN_4554 == 8'h2b ? _GEN_3425 : _GEN_2997; // @[executor.scala 473:84]
  wire [7:0] _GEN_3430 = mask_3[0] ? byte_768 : _GEN_2998; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3431 = mask_3[1] ? byte_769 : _GEN_2999; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3432 = mask_3[2] ? byte_770 : _GEN_3000; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3433 = mask_3[3] ? byte_771 : _GEN_3001; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3434 = _GEN_4554 == 8'h2c ? _GEN_3430 : _GEN_2998; // @[executor.scala 473:84]
  wire [7:0] _GEN_3435 = _GEN_4554 == 8'h2c ? _GEN_3431 : _GEN_2999; // @[executor.scala 473:84]
  wire [7:0] _GEN_3436 = _GEN_4554 == 8'h2c ? _GEN_3432 : _GEN_3000; // @[executor.scala 473:84]
  wire [7:0] _GEN_3437 = _GEN_4554 == 8'h2c ? _GEN_3433 : _GEN_3001; // @[executor.scala 473:84]
  wire [7:0] _GEN_3438 = mask_3[0] ? byte_768 : _GEN_3002; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3439 = mask_3[1] ? byte_769 : _GEN_3003; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3440 = mask_3[2] ? byte_770 : _GEN_3004; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3441 = mask_3[3] ? byte_771 : _GEN_3005; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3442 = _GEN_4554 == 8'h2d ? _GEN_3438 : _GEN_3002; // @[executor.scala 473:84]
  wire [7:0] _GEN_3443 = _GEN_4554 == 8'h2d ? _GEN_3439 : _GEN_3003; // @[executor.scala 473:84]
  wire [7:0] _GEN_3444 = _GEN_4554 == 8'h2d ? _GEN_3440 : _GEN_3004; // @[executor.scala 473:84]
  wire [7:0] _GEN_3445 = _GEN_4554 == 8'h2d ? _GEN_3441 : _GEN_3005; // @[executor.scala 473:84]
  wire [7:0] _GEN_3446 = mask_3[0] ? byte_768 : _GEN_3006; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3447 = mask_3[1] ? byte_769 : _GEN_3007; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3448 = mask_3[2] ? byte_770 : _GEN_3008; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3449 = mask_3[3] ? byte_771 : _GEN_3009; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3450 = _GEN_4554 == 8'h2e ? _GEN_3446 : _GEN_3006; // @[executor.scala 473:84]
  wire [7:0] _GEN_3451 = _GEN_4554 == 8'h2e ? _GEN_3447 : _GEN_3007; // @[executor.scala 473:84]
  wire [7:0] _GEN_3452 = _GEN_4554 == 8'h2e ? _GEN_3448 : _GEN_3008; // @[executor.scala 473:84]
  wire [7:0] _GEN_3453 = _GEN_4554 == 8'h2e ? _GEN_3449 : _GEN_3009; // @[executor.scala 473:84]
  wire [7:0] _GEN_3454 = mask_3[0] ? byte_768 : _GEN_3010; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3455 = mask_3[1] ? byte_769 : _GEN_3011; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3456 = mask_3[2] ? byte_770 : _GEN_3012; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3457 = mask_3[3] ? byte_771 : _GEN_3013; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3458 = _GEN_4554 == 8'h2f ? _GEN_3454 : _GEN_3010; // @[executor.scala 473:84]
  wire [7:0] _GEN_3459 = _GEN_4554 == 8'h2f ? _GEN_3455 : _GEN_3011; // @[executor.scala 473:84]
  wire [7:0] _GEN_3460 = _GEN_4554 == 8'h2f ? _GEN_3456 : _GEN_3012; // @[executor.scala 473:84]
  wire [7:0] _GEN_3461 = _GEN_4554 == 8'h2f ? _GEN_3457 : _GEN_3013; // @[executor.scala 473:84]
  wire [7:0] _GEN_3462 = mask_3[0] ? byte_768 : _GEN_3014; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3463 = mask_3[1] ? byte_769 : _GEN_3015; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3464 = mask_3[2] ? byte_770 : _GEN_3016; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3465 = mask_3[3] ? byte_771 : _GEN_3017; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3466 = _GEN_4554 == 8'h30 ? _GEN_3462 : _GEN_3014; // @[executor.scala 473:84]
  wire [7:0] _GEN_3467 = _GEN_4554 == 8'h30 ? _GEN_3463 : _GEN_3015; // @[executor.scala 473:84]
  wire [7:0] _GEN_3468 = _GEN_4554 == 8'h30 ? _GEN_3464 : _GEN_3016; // @[executor.scala 473:84]
  wire [7:0] _GEN_3469 = _GEN_4554 == 8'h30 ? _GEN_3465 : _GEN_3017; // @[executor.scala 473:84]
  wire [7:0] _GEN_3470 = mask_3[0] ? byte_768 : _GEN_3018; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3471 = mask_3[1] ? byte_769 : _GEN_3019; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3472 = mask_3[2] ? byte_770 : _GEN_3020; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3473 = mask_3[3] ? byte_771 : _GEN_3021; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3474 = _GEN_4554 == 8'h31 ? _GEN_3470 : _GEN_3018; // @[executor.scala 473:84]
  wire [7:0] _GEN_3475 = _GEN_4554 == 8'h31 ? _GEN_3471 : _GEN_3019; // @[executor.scala 473:84]
  wire [7:0] _GEN_3476 = _GEN_4554 == 8'h31 ? _GEN_3472 : _GEN_3020; // @[executor.scala 473:84]
  wire [7:0] _GEN_3477 = _GEN_4554 == 8'h31 ? _GEN_3473 : _GEN_3021; // @[executor.scala 473:84]
  wire [7:0] _GEN_3478 = mask_3[0] ? byte_768 : _GEN_3022; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3479 = mask_3[1] ? byte_769 : _GEN_3023; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3480 = mask_3[2] ? byte_770 : _GEN_3024; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3481 = mask_3[3] ? byte_771 : _GEN_3025; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3482 = _GEN_4554 == 8'h32 ? _GEN_3478 : _GEN_3022; // @[executor.scala 473:84]
  wire [7:0] _GEN_3483 = _GEN_4554 == 8'h32 ? _GEN_3479 : _GEN_3023; // @[executor.scala 473:84]
  wire [7:0] _GEN_3484 = _GEN_4554 == 8'h32 ? _GEN_3480 : _GEN_3024; // @[executor.scala 473:84]
  wire [7:0] _GEN_3485 = _GEN_4554 == 8'h32 ? _GEN_3481 : _GEN_3025; // @[executor.scala 473:84]
  wire [7:0] _GEN_3486 = mask_3[0] ? byte_768 : _GEN_3026; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3487 = mask_3[1] ? byte_769 : _GEN_3027; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3488 = mask_3[2] ? byte_770 : _GEN_3028; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3489 = mask_3[3] ? byte_771 : _GEN_3029; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3490 = _GEN_4554 == 8'h33 ? _GEN_3486 : _GEN_3026; // @[executor.scala 473:84]
  wire [7:0] _GEN_3491 = _GEN_4554 == 8'h33 ? _GEN_3487 : _GEN_3027; // @[executor.scala 473:84]
  wire [7:0] _GEN_3492 = _GEN_4554 == 8'h33 ? _GEN_3488 : _GEN_3028; // @[executor.scala 473:84]
  wire [7:0] _GEN_3493 = _GEN_4554 == 8'h33 ? _GEN_3489 : _GEN_3029; // @[executor.scala 473:84]
  wire [7:0] _GEN_3494 = mask_3[0] ? byte_768 : _GEN_3030; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3495 = mask_3[1] ? byte_769 : _GEN_3031; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3496 = mask_3[2] ? byte_770 : _GEN_3032; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3497 = mask_3[3] ? byte_771 : _GEN_3033; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3498 = _GEN_4554 == 8'h34 ? _GEN_3494 : _GEN_3030; // @[executor.scala 473:84]
  wire [7:0] _GEN_3499 = _GEN_4554 == 8'h34 ? _GEN_3495 : _GEN_3031; // @[executor.scala 473:84]
  wire [7:0] _GEN_3500 = _GEN_4554 == 8'h34 ? _GEN_3496 : _GEN_3032; // @[executor.scala 473:84]
  wire [7:0] _GEN_3501 = _GEN_4554 == 8'h34 ? _GEN_3497 : _GEN_3033; // @[executor.scala 473:84]
  wire [7:0] _GEN_3502 = mask_3[0] ? byte_768 : _GEN_3034; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3503 = mask_3[1] ? byte_769 : _GEN_3035; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3504 = mask_3[2] ? byte_770 : _GEN_3036; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3505 = mask_3[3] ? byte_771 : _GEN_3037; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3506 = _GEN_4554 == 8'h35 ? _GEN_3502 : _GEN_3034; // @[executor.scala 473:84]
  wire [7:0] _GEN_3507 = _GEN_4554 == 8'h35 ? _GEN_3503 : _GEN_3035; // @[executor.scala 473:84]
  wire [7:0] _GEN_3508 = _GEN_4554 == 8'h35 ? _GEN_3504 : _GEN_3036; // @[executor.scala 473:84]
  wire [7:0] _GEN_3509 = _GEN_4554 == 8'h35 ? _GEN_3505 : _GEN_3037; // @[executor.scala 473:84]
  wire [7:0] _GEN_3510 = mask_3[0] ? byte_768 : _GEN_3038; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3511 = mask_3[1] ? byte_769 : _GEN_3039; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3512 = mask_3[2] ? byte_770 : _GEN_3040; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3513 = mask_3[3] ? byte_771 : _GEN_3041; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3514 = _GEN_4554 == 8'h36 ? _GEN_3510 : _GEN_3038; // @[executor.scala 473:84]
  wire [7:0] _GEN_3515 = _GEN_4554 == 8'h36 ? _GEN_3511 : _GEN_3039; // @[executor.scala 473:84]
  wire [7:0] _GEN_3516 = _GEN_4554 == 8'h36 ? _GEN_3512 : _GEN_3040; // @[executor.scala 473:84]
  wire [7:0] _GEN_3517 = _GEN_4554 == 8'h36 ? _GEN_3513 : _GEN_3041; // @[executor.scala 473:84]
  wire [7:0] _GEN_3518 = mask_3[0] ? byte_768 : _GEN_3042; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3519 = mask_3[1] ? byte_769 : _GEN_3043; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3520 = mask_3[2] ? byte_770 : _GEN_3044; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3521 = mask_3[3] ? byte_771 : _GEN_3045; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3522 = _GEN_4554 == 8'h37 ? _GEN_3518 : _GEN_3042; // @[executor.scala 473:84]
  wire [7:0] _GEN_3523 = _GEN_4554 == 8'h37 ? _GEN_3519 : _GEN_3043; // @[executor.scala 473:84]
  wire [7:0] _GEN_3524 = _GEN_4554 == 8'h37 ? _GEN_3520 : _GEN_3044; // @[executor.scala 473:84]
  wire [7:0] _GEN_3525 = _GEN_4554 == 8'h37 ? _GEN_3521 : _GEN_3045; // @[executor.scala 473:84]
  wire [7:0] _GEN_3526 = mask_3[0] ? byte_768 : _GEN_3046; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3527 = mask_3[1] ? byte_769 : _GEN_3047; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3528 = mask_3[2] ? byte_770 : _GEN_3048; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3529 = mask_3[3] ? byte_771 : _GEN_3049; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3530 = _GEN_4554 == 8'h38 ? _GEN_3526 : _GEN_3046; // @[executor.scala 473:84]
  wire [7:0] _GEN_3531 = _GEN_4554 == 8'h38 ? _GEN_3527 : _GEN_3047; // @[executor.scala 473:84]
  wire [7:0] _GEN_3532 = _GEN_4554 == 8'h38 ? _GEN_3528 : _GEN_3048; // @[executor.scala 473:84]
  wire [7:0] _GEN_3533 = _GEN_4554 == 8'h38 ? _GEN_3529 : _GEN_3049; // @[executor.scala 473:84]
  wire [7:0] _GEN_3534 = mask_3[0] ? byte_768 : _GEN_3050; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3535 = mask_3[1] ? byte_769 : _GEN_3051; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3536 = mask_3[2] ? byte_770 : _GEN_3052; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3537 = mask_3[3] ? byte_771 : _GEN_3053; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3538 = _GEN_4554 == 8'h39 ? _GEN_3534 : _GEN_3050; // @[executor.scala 473:84]
  wire [7:0] _GEN_3539 = _GEN_4554 == 8'h39 ? _GEN_3535 : _GEN_3051; // @[executor.scala 473:84]
  wire [7:0] _GEN_3540 = _GEN_4554 == 8'h39 ? _GEN_3536 : _GEN_3052; // @[executor.scala 473:84]
  wire [7:0] _GEN_3541 = _GEN_4554 == 8'h39 ? _GEN_3537 : _GEN_3053; // @[executor.scala 473:84]
  wire [7:0] _GEN_3542 = mask_3[0] ? byte_768 : _GEN_3054; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3543 = mask_3[1] ? byte_769 : _GEN_3055; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3544 = mask_3[2] ? byte_770 : _GEN_3056; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3545 = mask_3[3] ? byte_771 : _GEN_3057; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3546 = _GEN_4554 == 8'h3a ? _GEN_3542 : _GEN_3054; // @[executor.scala 473:84]
  wire [7:0] _GEN_3547 = _GEN_4554 == 8'h3a ? _GEN_3543 : _GEN_3055; // @[executor.scala 473:84]
  wire [7:0] _GEN_3548 = _GEN_4554 == 8'h3a ? _GEN_3544 : _GEN_3056; // @[executor.scala 473:84]
  wire [7:0] _GEN_3549 = _GEN_4554 == 8'h3a ? _GEN_3545 : _GEN_3057; // @[executor.scala 473:84]
  wire [7:0] _GEN_3550 = mask_3[0] ? byte_768 : _GEN_3058; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3551 = mask_3[1] ? byte_769 : _GEN_3059; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3552 = mask_3[2] ? byte_770 : _GEN_3060; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3553 = mask_3[3] ? byte_771 : _GEN_3061; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3554 = _GEN_4554 == 8'h3b ? _GEN_3550 : _GEN_3058; // @[executor.scala 473:84]
  wire [7:0] _GEN_3555 = _GEN_4554 == 8'h3b ? _GEN_3551 : _GEN_3059; // @[executor.scala 473:84]
  wire [7:0] _GEN_3556 = _GEN_4554 == 8'h3b ? _GEN_3552 : _GEN_3060; // @[executor.scala 473:84]
  wire [7:0] _GEN_3557 = _GEN_4554 == 8'h3b ? _GEN_3553 : _GEN_3061; // @[executor.scala 473:84]
  wire [7:0] _GEN_3558 = mask_3[0] ? byte_768 : _GEN_3062; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3559 = mask_3[1] ? byte_769 : _GEN_3063; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3560 = mask_3[2] ? byte_770 : _GEN_3064; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3561 = mask_3[3] ? byte_771 : _GEN_3065; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3562 = _GEN_4554 == 8'h3c ? _GEN_3558 : _GEN_3062; // @[executor.scala 473:84]
  wire [7:0] _GEN_3563 = _GEN_4554 == 8'h3c ? _GEN_3559 : _GEN_3063; // @[executor.scala 473:84]
  wire [7:0] _GEN_3564 = _GEN_4554 == 8'h3c ? _GEN_3560 : _GEN_3064; // @[executor.scala 473:84]
  wire [7:0] _GEN_3565 = _GEN_4554 == 8'h3c ? _GEN_3561 : _GEN_3065; // @[executor.scala 473:84]
  wire [7:0] _GEN_3566 = mask_3[0] ? byte_768 : _GEN_3066; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3567 = mask_3[1] ? byte_769 : _GEN_3067; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3568 = mask_3[2] ? byte_770 : _GEN_3068; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3569 = mask_3[3] ? byte_771 : _GEN_3069; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3570 = _GEN_4554 == 8'h3d ? _GEN_3566 : _GEN_3066; // @[executor.scala 473:84]
  wire [7:0] _GEN_3571 = _GEN_4554 == 8'h3d ? _GEN_3567 : _GEN_3067; // @[executor.scala 473:84]
  wire [7:0] _GEN_3572 = _GEN_4554 == 8'h3d ? _GEN_3568 : _GEN_3068; // @[executor.scala 473:84]
  wire [7:0] _GEN_3573 = _GEN_4554 == 8'h3d ? _GEN_3569 : _GEN_3069; // @[executor.scala 473:84]
  wire [7:0] _GEN_3574 = mask_3[0] ? byte_768 : _GEN_3070; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3575 = mask_3[1] ? byte_769 : _GEN_3071; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3576 = mask_3[2] ? byte_770 : _GEN_3072; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3577 = mask_3[3] ? byte_771 : _GEN_3073; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3578 = _GEN_4554 == 8'h3e ? _GEN_3574 : _GEN_3070; // @[executor.scala 473:84]
  wire [7:0] _GEN_3579 = _GEN_4554 == 8'h3e ? _GEN_3575 : _GEN_3071; // @[executor.scala 473:84]
  wire [7:0] _GEN_3580 = _GEN_4554 == 8'h3e ? _GEN_3576 : _GEN_3072; // @[executor.scala 473:84]
  wire [7:0] _GEN_3581 = _GEN_4554 == 8'h3e ? _GEN_3577 : _GEN_3073; // @[executor.scala 473:84]
  wire [7:0] _GEN_3582 = mask_3[0] ? byte_768 : _GEN_3074; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3583 = mask_3[1] ? byte_769 : _GEN_3075; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3584 = mask_3[2] ? byte_770 : _GEN_3076; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3585 = mask_3[3] ? byte_771 : _GEN_3077; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3586 = _GEN_4554 == 8'h3f ? _GEN_3582 : _GEN_3074; // @[executor.scala 473:84]
  wire [7:0] _GEN_3587 = _GEN_4554 == 8'h3f ? _GEN_3583 : _GEN_3075; // @[executor.scala 473:84]
  wire [7:0] _GEN_3588 = _GEN_4554 == 8'h3f ? _GEN_3584 : _GEN_3076; // @[executor.scala 473:84]
  wire [7:0] _GEN_3589 = _GEN_4554 == 8'h3f ? _GEN_3585 : _GEN_3077; // @[executor.scala 473:84]
  wire [7:0] _GEN_3590 = opcode_3 != 4'h0 ? _GEN_3082 : _GEN_2822; // @[executor.scala 470:55]
  wire [7:0] _GEN_3591 = opcode_3 != 4'h0 ? _GEN_3083 : _GEN_2823; // @[executor.scala 470:55]
  wire [7:0] _GEN_3592 = opcode_3 != 4'h0 ? _GEN_3084 : _GEN_2824; // @[executor.scala 470:55]
  wire [7:0] _GEN_3593 = opcode_3 != 4'h0 ? _GEN_3085 : _GEN_2825; // @[executor.scala 470:55]
  wire [7:0] _GEN_3594 = opcode_3 != 4'h0 ? _GEN_3090 : _GEN_2826; // @[executor.scala 470:55]
  wire [7:0] _GEN_3595 = opcode_3 != 4'h0 ? _GEN_3091 : _GEN_2827; // @[executor.scala 470:55]
  wire [7:0] _GEN_3596 = opcode_3 != 4'h0 ? _GEN_3092 : _GEN_2828; // @[executor.scala 470:55]
  wire [7:0] _GEN_3597 = opcode_3 != 4'h0 ? _GEN_3093 : _GEN_2829; // @[executor.scala 470:55]
  wire [7:0] _GEN_3598 = opcode_3 != 4'h0 ? _GEN_3098 : _GEN_2830; // @[executor.scala 470:55]
  wire [7:0] _GEN_3599 = opcode_3 != 4'h0 ? _GEN_3099 : _GEN_2831; // @[executor.scala 470:55]
  wire [7:0] _GEN_3600 = opcode_3 != 4'h0 ? _GEN_3100 : _GEN_2832; // @[executor.scala 470:55]
  wire [7:0] _GEN_3601 = opcode_3 != 4'h0 ? _GEN_3101 : _GEN_2833; // @[executor.scala 470:55]
  wire [7:0] _GEN_3602 = opcode_3 != 4'h0 ? _GEN_3106 : _GEN_2834; // @[executor.scala 470:55]
  wire [7:0] _GEN_3603 = opcode_3 != 4'h0 ? _GEN_3107 : _GEN_2835; // @[executor.scala 470:55]
  wire [7:0] _GEN_3604 = opcode_3 != 4'h0 ? _GEN_3108 : _GEN_2836; // @[executor.scala 470:55]
  wire [7:0] _GEN_3605 = opcode_3 != 4'h0 ? _GEN_3109 : _GEN_2837; // @[executor.scala 470:55]
  wire [7:0] _GEN_3606 = opcode_3 != 4'h0 ? _GEN_3114 : _GEN_2838; // @[executor.scala 470:55]
  wire [7:0] _GEN_3607 = opcode_3 != 4'h0 ? _GEN_3115 : _GEN_2839; // @[executor.scala 470:55]
  wire [7:0] _GEN_3608 = opcode_3 != 4'h0 ? _GEN_3116 : _GEN_2840; // @[executor.scala 470:55]
  wire [7:0] _GEN_3609 = opcode_3 != 4'h0 ? _GEN_3117 : _GEN_2841; // @[executor.scala 470:55]
  wire [7:0] _GEN_3610 = opcode_3 != 4'h0 ? _GEN_3122 : _GEN_2842; // @[executor.scala 470:55]
  wire [7:0] _GEN_3611 = opcode_3 != 4'h0 ? _GEN_3123 : _GEN_2843; // @[executor.scala 470:55]
  wire [7:0] _GEN_3612 = opcode_3 != 4'h0 ? _GEN_3124 : _GEN_2844; // @[executor.scala 470:55]
  wire [7:0] _GEN_3613 = opcode_3 != 4'h0 ? _GEN_3125 : _GEN_2845; // @[executor.scala 470:55]
  wire [7:0] _GEN_3614 = opcode_3 != 4'h0 ? _GEN_3130 : _GEN_2846; // @[executor.scala 470:55]
  wire [7:0] _GEN_3615 = opcode_3 != 4'h0 ? _GEN_3131 : _GEN_2847; // @[executor.scala 470:55]
  wire [7:0] _GEN_3616 = opcode_3 != 4'h0 ? _GEN_3132 : _GEN_2848; // @[executor.scala 470:55]
  wire [7:0] _GEN_3617 = opcode_3 != 4'h0 ? _GEN_3133 : _GEN_2849; // @[executor.scala 470:55]
  wire [7:0] _GEN_3618 = opcode_3 != 4'h0 ? _GEN_3138 : _GEN_2850; // @[executor.scala 470:55]
  wire [7:0] _GEN_3619 = opcode_3 != 4'h0 ? _GEN_3139 : _GEN_2851; // @[executor.scala 470:55]
  wire [7:0] _GEN_3620 = opcode_3 != 4'h0 ? _GEN_3140 : _GEN_2852; // @[executor.scala 470:55]
  wire [7:0] _GEN_3621 = opcode_3 != 4'h0 ? _GEN_3141 : _GEN_2853; // @[executor.scala 470:55]
  wire [7:0] _GEN_3622 = opcode_3 != 4'h0 ? _GEN_3146 : _GEN_2854; // @[executor.scala 470:55]
  wire [7:0] _GEN_3623 = opcode_3 != 4'h0 ? _GEN_3147 : _GEN_2855; // @[executor.scala 470:55]
  wire [7:0] _GEN_3624 = opcode_3 != 4'h0 ? _GEN_3148 : _GEN_2856; // @[executor.scala 470:55]
  wire [7:0] _GEN_3625 = opcode_3 != 4'h0 ? _GEN_3149 : _GEN_2857; // @[executor.scala 470:55]
  wire [7:0] _GEN_3626 = opcode_3 != 4'h0 ? _GEN_3154 : _GEN_2858; // @[executor.scala 470:55]
  wire [7:0] _GEN_3627 = opcode_3 != 4'h0 ? _GEN_3155 : _GEN_2859; // @[executor.scala 470:55]
  wire [7:0] _GEN_3628 = opcode_3 != 4'h0 ? _GEN_3156 : _GEN_2860; // @[executor.scala 470:55]
  wire [7:0] _GEN_3629 = opcode_3 != 4'h0 ? _GEN_3157 : _GEN_2861; // @[executor.scala 470:55]
  wire [7:0] _GEN_3630 = opcode_3 != 4'h0 ? _GEN_3162 : _GEN_2862; // @[executor.scala 470:55]
  wire [7:0] _GEN_3631 = opcode_3 != 4'h0 ? _GEN_3163 : _GEN_2863; // @[executor.scala 470:55]
  wire [7:0] _GEN_3632 = opcode_3 != 4'h0 ? _GEN_3164 : _GEN_2864; // @[executor.scala 470:55]
  wire [7:0] _GEN_3633 = opcode_3 != 4'h0 ? _GEN_3165 : _GEN_2865; // @[executor.scala 470:55]
  wire [7:0] _GEN_3634 = opcode_3 != 4'h0 ? _GEN_3170 : _GEN_2866; // @[executor.scala 470:55]
  wire [7:0] _GEN_3635 = opcode_3 != 4'h0 ? _GEN_3171 : _GEN_2867; // @[executor.scala 470:55]
  wire [7:0] _GEN_3636 = opcode_3 != 4'h0 ? _GEN_3172 : _GEN_2868; // @[executor.scala 470:55]
  wire [7:0] _GEN_3637 = opcode_3 != 4'h0 ? _GEN_3173 : _GEN_2869; // @[executor.scala 470:55]
  wire [7:0] _GEN_3638 = opcode_3 != 4'h0 ? _GEN_3178 : _GEN_2870; // @[executor.scala 470:55]
  wire [7:0] _GEN_3639 = opcode_3 != 4'h0 ? _GEN_3179 : _GEN_2871; // @[executor.scala 470:55]
  wire [7:0] _GEN_3640 = opcode_3 != 4'h0 ? _GEN_3180 : _GEN_2872; // @[executor.scala 470:55]
  wire [7:0] _GEN_3641 = opcode_3 != 4'h0 ? _GEN_3181 : _GEN_2873; // @[executor.scala 470:55]
  wire [7:0] _GEN_3642 = opcode_3 != 4'h0 ? _GEN_3186 : _GEN_2874; // @[executor.scala 470:55]
  wire [7:0] _GEN_3643 = opcode_3 != 4'h0 ? _GEN_3187 : _GEN_2875; // @[executor.scala 470:55]
  wire [7:0] _GEN_3644 = opcode_3 != 4'h0 ? _GEN_3188 : _GEN_2876; // @[executor.scala 470:55]
  wire [7:0] _GEN_3645 = opcode_3 != 4'h0 ? _GEN_3189 : _GEN_2877; // @[executor.scala 470:55]
  wire [7:0] _GEN_3646 = opcode_3 != 4'h0 ? _GEN_3194 : _GEN_2878; // @[executor.scala 470:55]
  wire [7:0] _GEN_3647 = opcode_3 != 4'h0 ? _GEN_3195 : _GEN_2879; // @[executor.scala 470:55]
  wire [7:0] _GEN_3648 = opcode_3 != 4'h0 ? _GEN_3196 : _GEN_2880; // @[executor.scala 470:55]
  wire [7:0] _GEN_3649 = opcode_3 != 4'h0 ? _GEN_3197 : _GEN_2881; // @[executor.scala 470:55]
  wire [7:0] _GEN_3650 = opcode_3 != 4'h0 ? _GEN_3202 : _GEN_2882; // @[executor.scala 470:55]
  wire [7:0] _GEN_3651 = opcode_3 != 4'h0 ? _GEN_3203 : _GEN_2883; // @[executor.scala 470:55]
  wire [7:0] _GEN_3652 = opcode_3 != 4'h0 ? _GEN_3204 : _GEN_2884; // @[executor.scala 470:55]
  wire [7:0] _GEN_3653 = opcode_3 != 4'h0 ? _GEN_3205 : _GEN_2885; // @[executor.scala 470:55]
  wire [7:0] _GEN_3654 = opcode_3 != 4'h0 ? _GEN_3210 : _GEN_2886; // @[executor.scala 470:55]
  wire [7:0] _GEN_3655 = opcode_3 != 4'h0 ? _GEN_3211 : _GEN_2887; // @[executor.scala 470:55]
  wire [7:0] _GEN_3656 = opcode_3 != 4'h0 ? _GEN_3212 : _GEN_2888; // @[executor.scala 470:55]
  wire [7:0] _GEN_3657 = opcode_3 != 4'h0 ? _GEN_3213 : _GEN_2889; // @[executor.scala 470:55]
  wire [7:0] _GEN_3658 = opcode_3 != 4'h0 ? _GEN_3218 : _GEN_2890; // @[executor.scala 470:55]
  wire [7:0] _GEN_3659 = opcode_3 != 4'h0 ? _GEN_3219 : _GEN_2891; // @[executor.scala 470:55]
  wire [7:0] _GEN_3660 = opcode_3 != 4'h0 ? _GEN_3220 : _GEN_2892; // @[executor.scala 470:55]
  wire [7:0] _GEN_3661 = opcode_3 != 4'h0 ? _GEN_3221 : _GEN_2893; // @[executor.scala 470:55]
  wire [7:0] _GEN_3662 = opcode_3 != 4'h0 ? _GEN_3226 : _GEN_2894; // @[executor.scala 470:55]
  wire [7:0] _GEN_3663 = opcode_3 != 4'h0 ? _GEN_3227 : _GEN_2895; // @[executor.scala 470:55]
  wire [7:0] _GEN_3664 = opcode_3 != 4'h0 ? _GEN_3228 : _GEN_2896; // @[executor.scala 470:55]
  wire [7:0] _GEN_3665 = opcode_3 != 4'h0 ? _GEN_3229 : _GEN_2897; // @[executor.scala 470:55]
  wire [7:0] _GEN_3666 = opcode_3 != 4'h0 ? _GEN_3234 : _GEN_2898; // @[executor.scala 470:55]
  wire [7:0] _GEN_3667 = opcode_3 != 4'h0 ? _GEN_3235 : _GEN_2899; // @[executor.scala 470:55]
  wire [7:0] _GEN_3668 = opcode_3 != 4'h0 ? _GEN_3236 : _GEN_2900; // @[executor.scala 470:55]
  wire [7:0] _GEN_3669 = opcode_3 != 4'h0 ? _GEN_3237 : _GEN_2901; // @[executor.scala 470:55]
  wire [7:0] _GEN_3670 = opcode_3 != 4'h0 ? _GEN_3242 : _GEN_2902; // @[executor.scala 470:55]
  wire [7:0] _GEN_3671 = opcode_3 != 4'h0 ? _GEN_3243 : _GEN_2903; // @[executor.scala 470:55]
  wire [7:0] _GEN_3672 = opcode_3 != 4'h0 ? _GEN_3244 : _GEN_2904; // @[executor.scala 470:55]
  wire [7:0] _GEN_3673 = opcode_3 != 4'h0 ? _GEN_3245 : _GEN_2905; // @[executor.scala 470:55]
  wire [7:0] _GEN_3674 = opcode_3 != 4'h0 ? _GEN_3250 : _GEN_2906; // @[executor.scala 470:55]
  wire [7:0] _GEN_3675 = opcode_3 != 4'h0 ? _GEN_3251 : _GEN_2907; // @[executor.scala 470:55]
  wire [7:0] _GEN_3676 = opcode_3 != 4'h0 ? _GEN_3252 : _GEN_2908; // @[executor.scala 470:55]
  wire [7:0] _GEN_3677 = opcode_3 != 4'h0 ? _GEN_3253 : _GEN_2909; // @[executor.scala 470:55]
  wire [7:0] _GEN_3678 = opcode_3 != 4'h0 ? _GEN_3258 : _GEN_2910; // @[executor.scala 470:55]
  wire [7:0] _GEN_3679 = opcode_3 != 4'h0 ? _GEN_3259 : _GEN_2911; // @[executor.scala 470:55]
  wire [7:0] _GEN_3680 = opcode_3 != 4'h0 ? _GEN_3260 : _GEN_2912; // @[executor.scala 470:55]
  wire [7:0] _GEN_3681 = opcode_3 != 4'h0 ? _GEN_3261 : _GEN_2913; // @[executor.scala 470:55]
  wire [7:0] _GEN_3682 = opcode_3 != 4'h0 ? _GEN_3266 : _GEN_2914; // @[executor.scala 470:55]
  wire [7:0] _GEN_3683 = opcode_3 != 4'h0 ? _GEN_3267 : _GEN_2915; // @[executor.scala 470:55]
  wire [7:0] _GEN_3684 = opcode_3 != 4'h0 ? _GEN_3268 : _GEN_2916; // @[executor.scala 470:55]
  wire [7:0] _GEN_3685 = opcode_3 != 4'h0 ? _GEN_3269 : _GEN_2917; // @[executor.scala 470:55]
  wire [7:0] _GEN_3686 = opcode_3 != 4'h0 ? _GEN_3274 : _GEN_2918; // @[executor.scala 470:55]
  wire [7:0] _GEN_3687 = opcode_3 != 4'h0 ? _GEN_3275 : _GEN_2919; // @[executor.scala 470:55]
  wire [7:0] _GEN_3688 = opcode_3 != 4'h0 ? _GEN_3276 : _GEN_2920; // @[executor.scala 470:55]
  wire [7:0] _GEN_3689 = opcode_3 != 4'h0 ? _GEN_3277 : _GEN_2921; // @[executor.scala 470:55]
  wire [7:0] _GEN_3690 = opcode_3 != 4'h0 ? _GEN_3282 : _GEN_2922; // @[executor.scala 470:55]
  wire [7:0] _GEN_3691 = opcode_3 != 4'h0 ? _GEN_3283 : _GEN_2923; // @[executor.scala 470:55]
  wire [7:0] _GEN_3692 = opcode_3 != 4'h0 ? _GEN_3284 : _GEN_2924; // @[executor.scala 470:55]
  wire [7:0] _GEN_3693 = opcode_3 != 4'h0 ? _GEN_3285 : _GEN_2925; // @[executor.scala 470:55]
  wire [7:0] _GEN_3694 = opcode_3 != 4'h0 ? _GEN_3290 : _GEN_2926; // @[executor.scala 470:55]
  wire [7:0] _GEN_3695 = opcode_3 != 4'h0 ? _GEN_3291 : _GEN_2927; // @[executor.scala 470:55]
  wire [7:0] _GEN_3696 = opcode_3 != 4'h0 ? _GEN_3292 : _GEN_2928; // @[executor.scala 470:55]
  wire [7:0] _GEN_3697 = opcode_3 != 4'h0 ? _GEN_3293 : _GEN_2929; // @[executor.scala 470:55]
  wire [7:0] _GEN_3698 = opcode_3 != 4'h0 ? _GEN_3298 : _GEN_2930; // @[executor.scala 470:55]
  wire [7:0] _GEN_3699 = opcode_3 != 4'h0 ? _GEN_3299 : _GEN_2931; // @[executor.scala 470:55]
  wire [7:0] _GEN_3700 = opcode_3 != 4'h0 ? _GEN_3300 : _GEN_2932; // @[executor.scala 470:55]
  wire [7:0] _GEN_3701 = opcode_3 != 4'h0 ? _GEN_3301 : _GEN_2933; // @[executor.scala 470:55]
  wire [7:0] _GEN_3702 = opcode_3 != 4'h0 ? _GEN_3306 : _GEN_2934; // @[executor.scala 470:55]
  wire [7:0] _GEN_3703 = opcode_3 != 4'h0 ? _GEN_3307 : _GEN_2935; // @[executor.scala 470:55]
  wire [7:0] _GEN_3704 = opcode_3 != 4'h0 ? _GEN_3308 : _GEN_2936; // @[executor.scala 470:55]
  wire [7:0] _GEN_3705 = opcode_3 != 4'h0 ? _GEN_3309 : _GEN_2937; // @[executor.scala 470:55]
  wire [7:0] _GEN_3706 = opcode_3 != 4'h0 ? _GEN_3314 : _GEN_2938; // @[executor.scala 470:55]
  wire [7:0] _GEN_3707 = opcode_3 != 4'h0 ? _GEN_3315 : _GEN_2939; // @[executor.scala 470:55]
  wire [7:0] _GEN_3708 = opcode_3 != 4'h0 ? _GEN_3316 : _GEN_2940; // @[executor.scala 470:55]
  wire [7:0] _GEN_3709 = opcode_3 != 4'h0 ? _GEN_3317 : _GEN_2941; // @[executor.scala 470:55]
  wire [7:0] _GEN_3710 = opcode_3 != 4'h0 ? _GEN_3322 : _GEN_2942; // @[executor.scala 470:55]
  wire [7:0] _GEN_3711 = opcode_3 != 4'h0 ? _GEN_3323 : _GEN_2943; // @[executor.scala 470:55]
  wire [7:0] _GEN_3712 = opcode_3 != 4'h0 ? _GEN_3324 : _GEN_2944; // @[executor.scala 470:55]
  wire [7:0] _GEN_3713 = opcode_3 != 4'h0 ? _GEN_3325 : _GEN_2945; // @[executor.scala 470:55]
  wire [7:0] _GEN_3714 = opcode_3 != 4'h0 ? _GEN_3330 : _GEN_2946; // @[executor.scala 470:55]
  wire [7:0] _GEN_3715 = opcode_3 != 4'h0 ? _GEN_3331 : _GEN_2947; // @[executor.scala 470:55]
  wire [7:0] _GEN_3716 = opcode_3 != 4'h0 ? _GEN_3332 : _GEN_2948; // @[executor.scala 470:55]
  wire [7:0] _GEN_3717 = opcode_3 != 4'h0 ? _GEN_3333 : _GEN_2949; // @[executor.scala 470:55]
  wire [7:0] _GEN_3718 = opcode_3 != 4'h0 ? _GEN_3338 : _GEN_2950; // @[executor.scala 470:55]
  wire [7:0] _GEN_3719 = opcode_3 != 4'h0 ? _GEN_3339 : _GEN_2951; // @[executor.scala 470:55]
  wire [7:0] _GEN_3720 = opcode_3 != 4'h0 ? _GEN_3340 : _GEN_2952; // @[executor.scala 470:55]
  wire [7:0] _GEN_3721 = opcode_3 != 4'h0 ? _GEN_3341 : _GEN_2953; // @[executor.scala 470:55]
  wire [7:0] _GEN_3722 = opcode_3 != 4'h0 ? _GEN_3346 : _GEN_2954; // @[executor.scala 470:55]
  wire [7:0] _GEN_3723 = opcode_3 != 4'h0 ? _GEN_3347 : _GEN_2955; // @[executor.scala 470:55]
  wire [7:0] _GEN_3724 = opcode_3 != 4'h0 ? _GEN_3348 : _GEN_2956; // @[executor.scala 470:55]
  wire [7:0] _GEN_3725 = opcode_3 != 4'h0 ? _GEN_3349 : _GEN_2957; // @[executor.scala 470:55]
  wire [7:0] _GEN_3726 = opcode_3 != 4'h0 ? _GEN_3354 : _GEN_2958; // @[executor.scala 470:55]
  wire [7:0] _GEN_3727 = opcode_3 != 4'h0 ? _GEN_3355 : _GEN_2959; // @[executor.scala 470:55]
  wire [7:0] _GEN_3728 = opcode_3 != 4'h0 ? _GEN_3356 : _GEN_2960; // @[executor.scala 470:55]
  wire [7:0] _GEN_3729 = opcode_3 != 4'h0 ? _GEN_3357 : _GEN_2961; // @[executor.scala 470:55]
  wire [7:0] _GEN_3730 = opcode_3 != 4'h0 ? _GEN_3362 : _GEN_2962; // @[executor.scala 470:55]
  wire [7:0] _GEN_3731 = opcode_3 != 4'h0 ? _GEN_3363 : _GEN_2963; // @[executor.scala 470:55]
  wire [7:0] _GEN_3732 = opcode_3 != 4'h0 ? _GEN_3364 : _GEN_2964; // @[executor.scala 470:55]
  wire [7:0] _GEN_3733 = opcode_3 != 4'h0 ? _GEN_3365 : _GEN_2965; // @[executor.scala 470:55]
  wire [7:0] _GEN_3734 = opcode_3 != 4'h0 ? _GEN_3370 : _GEN_2966; // @[executor.scala 470:55]
  wire [7:0] _GEN_3735 = opcode_3 != 4'h0 ? _GEN_3371 : _GEN_2967; // @[executor.scala 470:55]
  wire [7:0] _GEN_3736 = opcode_3 != 4'h0 ? _GEN_3372 : _GEN_2968; // @[executor.scala 470:55]
  wire [7:0] _GEN_3737 = opcode_3 != 4'h0 ? _GEN_3373 : _GEN_2969; // @[executor.scala 470:55]
  wire [7:0] _GEN_3738 = opcode_3 != 4'h0 ? _GEN_3378 : _GEN_2970; // @[executor.scala 470:55]
  wire [7:0] _GEN_3739 = opcode_3 != 4'h0 ? _GEN_3379 : _GEN_2971; // @[executor.scala 470:55]
  wire [7:0] _GEN_3740 = opcode_3 != 4'h0 ? _GEN_3380 : _GEN_2972; // @[executor.scala 470:55]
  wire [7:0] _GEN_3741 = opcode_3 != 4'h0 ? _GEN_3381 : _GEN_2973; // @[executor.scala 470:55]
  wire [7:0] _GEN_3742 = opcode_3 != 4'h0 ? _GEN_3386 : _GEN_2974; // @[executor.scala 470:55]
  wire [7:0] _GEN_3743 = opcode_3 != 4'h0 ? _GEN_3387 : _GEN_2975; // @[executor.scala 470:55]
  wire [7:0] _GEN_3744 = opcode_3 != 4'h0 ? _GEN_3388 : _GEN_2976; // @[executor.scala 470:55]
  wire [7:0] _GEN_3745 = opcode_3 != 4'h0 ? _GEN_3389 : _GEN_2977; // @[executor.scala 470:55]
  wire [7:0] _GEN_3746 = opcode_3 != 4'h0 ? _GEN_3394 : _GEN_2978; // @[executor.scala 470:55]
  wire [7:0] _GEN_3747 = opcode_3 != 4'h0 ? _GEN_3395 : _GEN_2979; // @[executor.scala 470:55]
  wire [7:0] _GEN_3748 = opcode_3 != 4'h0 ? _GEN_3396 : _GEN_2980; // @[executor.scala 470:55]
  wire [7:0] _GEN_3749 = opcode_3 != 4'h0 ? _GEN_3397 : _GEN_2981; // @[executor.scala 470:55]
  wire [7:0] _GEN_3750 = opcode_3 != 4'h0 ? _GEN_3402 : _GEN_2982; // @[executor.scala 470:55]
  wire [7:0] _GEN_3751 = opcode_3 != 4'h0 ? _GEN_3403 : _GEN_2983; // @[executor.scala 470:55]
  wire [7:0] _GEN_3752 = opcode_3 != 4'h0 ? _GEN_3404 : _GEN_2984; // @[executor.scala 470:55]
  wire [7:0] _GEN_3753 = opcode_3 != 4'h0 ? _GEN_3405 : _GEN_2985; // @[executor.scala 470:55]
  wire [7:0] _GEN_3754 = opcode_3 != 4'h0 ? _GEN_3410 : _GEN_2986; // @[executor.scala 470:55]
  wire [7:0] _GEN_3755 = opcode_3 != 4'h0 ? _GEN_3411 : _GEN_2987; // @[executor.scala 470:55]
  wire [7:0] _GEN_3756 = opcode_3 != 4'h0 ? _GEN_3412 : _GEN_2988; // @[executor.scala 470:55]
  wire [7:0] _GEN_3757 = opcode_3 != 4'h0 ? _GEN_3413 : _GEN_2989; // @[executor.scala 470:55]
  wire [7:0] _GEN_3758 = opcode_3 != 4'h0 ? _GEN_3418 : _GEN_2990; // @[executor.scala 470:55]
  wire [7:0] _GEN_3759 = opcode_3 != 4'h0 ? _GEN_3419 : _GEN_2991; // @[executor.scala 470:55]
  wire [7:0] _GEN_3760 = opcode_3 != 4'h0 ? _GEN_3420 : _GEN_2992; // @[executor.scala 470:55]
  wire [7:0] _GEN_3761 = opcode_3 != 4'h0 ? _GEN_3421 : _GEN_2993; // @[executor.scala 470:55]
  wire [7:0] _GEN_3762 = opcode_3 != 4'h0 ? _GEN_3426 : _GEN_2994; // @[executor.scala 470:55]
  wire [7:0] _GEN_3763 = opcode_3 != 4'h0 ? _GEN_3427 : _GEN_2995; // @[executor.scala 470:55]
  wire [7:0] _GEN_3764 = opcode_3 != 4'h0 ? _GEN_3428 : _GEN_2996; // @[executor.scala 470:55]
  wire [7:0] _GEN_3765 = opcode_3 != 4'h0 ? _GEN_3429 : _GEN_2997; // @[executor.scala 470:55]
  wire [7:0] _GEN_3766 = opcode_3 != 4'h0 ? _GEN_3434 : _GEN_2998; // @[executor.scala 470:55]
  wire [7:0] _GEN_3767 = opcode_3 != 4'h0 ? _GEN_3435 : _GEN_2999; // @[executor.scala 470:55]
  wire [7:0] _GEN_3768 = opcode_3 != 4'h0 ? _GEN_3436 : _GEN_3000; // @[executor.scala 470:55]
  wire [7:0] _GEN_3769 = opcode_3 != 4'h0 ? _GEN_3437 : _GEN_3001; // @[executor.scala 470:55]
  wire [7:0] _GEN_3770 = opcode_3 != 4'h0 ? _GEN_3442 : _GEN_3002; // @[executor.scala 470:55]
  wire [7:0] _GEN_3771 = opcode_3 != 4'h0 ? _GEN_3443 : _GEN_3003; // @[executor.scala 470:55]
  wire [7:0] _GEN_3772 = opcode_3 != 4'h0 ? _GEN_3444 : _GEN_3004; // @[executor.scala 470:55]
  wire [7:0] _GEN_3773 = opcode_3 != 4'h0 ? _GEN_3445 : _GEN_3005; // @[executor.scala 470:55]
  wire [7:0] _GEN_3774 = opcode_3 != 4'h0 ? _GEN_3450 : _GEN_3006; // @[executor.scala 470:55]
  wire [7:0] _GEN_3775 = opcode_3 != 4'h0 ? _GEN_3451 : _GEN_3007; // @[executor.scala 470:55]
  wire [7:0] _GEN_3776 = opcode_3 != 4'h0 ? _GEN_3452 : _GEN_3008; // @[executor.scala 470:55]
  wire [7:0] _GEN_3777 = opcode_3 != 4'h0 ? _GEN_3453 : _GEN_3009; // @[executor.scala 470:55]
  wire [7:0] _GEN_3778 = opcode_3 != 4'h0 ? _GEN_3458 : _GEN_3010; // @[executor.scala 470:55]
  wire [7:0] _GEN_3779 = opcode_3 != 4'h0 ? _GEN_3459 : _GEN_3011; // @[executor.scala 470:55]
  wire [7:0] _GEN_3780 = opcode_3 != 4'h0 ? _GEN_3460 : _GEN_3012; // @[executor.scala 470:55]
  wire [7:0] _GEN_3781 = opcode_3 != 4'h0 ? _GEN_3461 : _GEN_3013; // @[executor.scala 470:55]
  wire [7:0] _GEN_3782 = opcode_3 != 4'h0 ? _GEN_3466 : _GEN_3014; // @[executor.scala 470:55]
  wire [7:0] _GEN_3783 = opcode_3 != 4'h0 ? _GEN_3467 : _GEN_3015; // @[executor.scala 470:55]
  wire [7:0] _GEN_3784 = opcode_3 != 4'h0 ? _GEN_3468 : _GEN_3016; // @[executor.scala 470:55]
  wire [7:0] _GEN_3785 = opcode_3 != 4'h0 ? _GEN_3469 : _GEN_3017; // @[executor.scala 470:55]
  wire [7:0] _GEN_3786 = opcode_3 != 4'h0 ? _GEN_3474 : _GEN_3018; // @[executor.scala 470:55]
  wire [7:0] _GEN_3787 = opcode_3 != 4'h0 ? _GEN_3475 : _GEN_3019; // @[executor.scala 470:55]
  wire [7:0] _GEN_3788 = opcode_3 != 4'h0 ? _GEN_3476 : _GEN_3020; // @[executor.scala 470:55]
  wire [7:0] _GEN_3789 = opcode_3 != 4'h0 ? _GEN_3477 : _GEN_3021; // @[executor.scala 470:55]
  wire [7:0] _GEN_3790 = opcode_3 != 4'h0 ? _GEN_3482 : _GEN_3022; // @[executor.scala 470:55]
  wire [7:0] _GEN_3791 = opcode_3 != 4'h0 ? _GEN_3483 : _GEN_3023; // @[executor.scala 470:55]
  wire [7:0] _GEN_3792 = opcode_3 != 4'h0 ? _GEN_3484 : _GEN_3024; // @[executor.scala 470:55]
  wire [7:0] _GEN_3793 = opcode_3 != 4'h0 ? _GEN_3485 : _GEN_3025; // @[executor.scala 470:55]
  wire [7:0] _GEN_3794 = opcode_3 != 4'h0 ? _GEN_3490 : _GEN_3026; // @[executor.scala 470:55]
  wire [7:0] _GEN_3795 = opcode_3 != 4'h0 ? _GEN_3491 : _GEN_3027; // @[executor.scala 470:55]
  wire [7:0] _GEN_3796 = opcode_3 != 4'h0 ? _GEN_3492 : _GEN_3028; // @[executor.scala 470:55]
  wire [7:0] _GEN_3797 = opcode_3 != 4'h0 ? _GEN_3493 : _GEN_3029; // @[executor.scala 470:55]
  wire [7:0] _GEN_3798 = opcode_3 != 4'h0 ? _GEN_3498 : _GEN_3030; // @[executor.scala 470:55]
  wire [7:0] _GEN_3799 = opcode_3 != 4'h0 ? _GEN_3499 : _GEN_3031; // @[executor.scala 470:55]
  wire [7:0] _GEN_3800 = opcode_3 != 4'h0 ? _GEN_3500 : _GEN_3032; // @[executor.scala 470:55]
  wire [7:0] _GEN_3801 = opcode_3 != 4'h0 ? _GEN_3501 : _GEN_3033; // @[executor.scala 470:55]
  wire [7:0] _GEN_3802 = opcode_3 != 4'h0 ? _GEN_3506 : _GEN_3034; // @[executor.scala 470:55]
  wire [7:0] _GEN_3803 = opcode_3 != 4'h0 ? _GEN_3507 : _GEN_3035; // @[executor.scala 470:55]
  wire [7:0] _GEN_3804 = opcode_3 != 4'h0 ? _GEN_3508 : _GEN_3036; // @[executor.scala 470:55]
  wire [7:0] _GEN_3805 = opcode_3 != 4'h0 ? _GEN_3509 : _GEN_3037; // @[executor.scala 470:55]
  wire [7:0] _GEN_3806 = opcode_3 != 4'h0 ? _GEN_3514 : _GEN_3038; // @[executor.scala 470:55]
  wire [7:0] _GEN_3807 = opcode_3 != 4'h0 ? _GEN_3515 : _GEN_3039; // @[executor.scala 470:55]
  wire [7:0] _GEN_3808 = opcode_3 != 4'h0 ? _GEN_3516 : _GEN_3040; // @[executor.scala 470:55]
  wire [7:0] _GEN_3809 = opcode_3 != 4'h0 ? _GEN_3517 : _GEN_3041; // @[executor.scala 470:55]
  wire [7:0] _GEN_3810 = opcode_3 != 4'h0 ? _GEN_3522 : _GEN_3042; // @[executor.scala 470:55]
  wire [7:0] _GEN_3811 = opcode_3 != 4'h0 ? _GEN_3523 : _GEN_3043; // @[executor.scala 470:55]
  wire [7:0] _GEN_3812 = opcode_3 != 4'h0 ? _GEN_3524 : _GEN_3044; // @[executor.scala 470:55]
  wire [7:0] _GEN_3813 = opcode_3 != 4'h0 ? _GEN_3525 : _GEN_3045; // @[executor.scala 470:55]
  wire [7:0] _GEN_3814 = opcode_3 != 4'h0 ? _GEN_3530 : _GEN_3046; // @[executor.scala 470:55]
  wire [7:0] _GEN_3815 = opcode_3 != 4'h0 ? _GEN_3531 : _GEN_3047; // @[executor.scala 470:55]
  wire [7:0] _GEN_3816 = opcode_3 != 4'h0 ? _GEN_3532 : _GEN_3048; // @[executor.scala 470:55]
  wire [7:0] _GEN_3817 = opcode_3 != 4'h0 ? _GEN_3533 : _GEN_3049; // @[executor.scala 470:55]
  wire [7:0] _GEN_3818 = opcode_3 != 4'h0 ? _GEN_3538 : _GEN_3050; // @[executor.scala 470:55]
  wire [7:0] _GEN_3819 = opcode_3 != 4'h0 ? _GEN_3539 : _GEN_3051; // @[executor.scala 470:55]
  wire [7:0] _GEN_3820 = opcode_3 != 4'h0 ? _GEN_3540 : _GEN_3052; // @[executor.scala 470:55]
  wire [7:0] _GEN_3821 = opcode_3 != 4'h0 ? _GEN_3541 : _GEN_3053; // @[executor.scala 470:55]
  wire [7:0] _GEN_3822 = opcode_3 != 4'h0 ? _GEN_3546 : _GEN_3054; // @[executor.scala 470:55]
  wire [7:0] _GEN_3823 = opcode_3 != 4'h0 ? _GEN_3547 : _GEN_3055; // @[executor.scala 470:55]
  wire [7:0] _GEN_3824 = opcode_3 != 4'h0 ? _GEN_3548 : _GEN_3056; // @[executor.scala 470:55]
  wire [7:0] _GEN_3825 = opcode_3 != 4'h0 ? _GEN_3549 : _GEN_3057; // @[executor.scala 470:55]
  wire [7:0] _GEN_3826 = opcode_3 != 4'h0 ? _GEN_3554 : _GEN_3058; // @[executor.scala 470:55]
  wire [7:0] _GEN_3827 = opcode_3 != 4'h0 ? _GEN_3555 : _GEN_3059; // @[executor.scala 470:55]
  wire [7:0] _GEN_3828 = opcode_3 != 4'h0 ? _GEN_3556 : _GEN_3060; // @[executor.scala 470:55]
  wire [7:0] _GEN_3829 = opcode_3 != 4'h0 ? _GEN_3557 : _GEN_3061; // @[executor.scala 470:55]
  wire [7:0] _GEN_3830 = opcode_3 != 4'h0 ? _GEN_3562 : _GEN_3062; // @[executor.scala 470:55]
  wire [7:0] _GEN_3831 = opcode_3 != 4'h0 ? _GEN_3563 : _GEN_3063; // @[executor.scala 470:55]
  wire [7:0] _GEN_3832 = opcode_3 != 4'h0 ? _GEN_3564 : _GEN_3064; // @[executor.scala 470:55]
  wire [7:0] _GEN_3833 = opcode_3 != 4'h0 ? _GEN_3565 : _GEN_3065; // @[executor.scala 470:55]
  wire [7:0] _GEN_3834 = opcode_3 != 4'h0 ? _GEN_3570 : _GEN_3066; // @[executor.scala 470:55]
  wire [7:0] _GEN_3835 = opcode_3 != 4'h0 ? _GEN_3571 : _GEN_3067; // @[executor.scala 470:55]
  wire [7:0] _GEN_3836 = opcode_3 != 4'h0 ? _GEN_3572 : _GEN_3068; // @[executor.scala 470:55]
  wire [7:0] _GEN_3837 = opcode_3 != 4'h0 ? _GEN_3573 : _GEN_3069; // @[executor.scala 470:55]
  wire [7:0] _GEN_3838 = opcode_3 != 4'h0 ? _GEN_3578 : _GEN_3070; // @[executor.scala 470:55]
  wire [7:0] _GEN_3839 = opcode_3 != 4'h0 ? _GEN_3579 : _GEN_3071; // @[executor.scala 470:55]
  wire [7:0] _GEN_3840 = opcode_3 != 4'h0 ? _GEN_3580 : _GEN_3072; // @[executor.scala 470:55]
  wire [7:0] _GEN_3841 = opcode_3 != 4'h0 ? _GEN_3581 : _GEN_3073; // @[executor.scala 470:55]
  wire [7:0] _GEN_3842 = opcode_3 != 4'h0 ? _GEN_3586 : _GEN_3074; // @[executor.scala 470:55]
  wire [7:0] _GEN_3843 = opcode_3 != 4'h0 ? _GEN_3587 : _GEN_3075; // @[executor.scala 470:55]
  wire [7:0] _GEN_3844 = opcode_3 != 4'h0 ? _GEN_3588 : _GEN_3076; // @[executor.scala 470:55]
  wire [7:0] _GEN_3845 = opcode_3 != 4'h0 ? _GEN_3589 : _GEN_3077; // @[executor.scala 470:55]
  wire [7:0] _GEN_3848 = opcode_3 == 4'hf ? _GEN_2822 : _GEN_3590; // @[executor.scala 466:52]
  wire [7:0] _GEN_3849 = opcode_3 == 4'hf ? _GEN_2823 : _GEN_3591; // @[executor.scala 466:52]
  wire [7:0] _GEN_3850 = opcode_3 == 4'hf ? _GEN_2824 : _GEN_3592; // @[executor.scala 466:52]
  wire [7:0] _GEN_3851 = opcode_3 == 4'hf ? _GEN_2825 : _GEN_3593; // @[executor.scala 466:52]
  wire [7:0] _GEN_3852 = opcode_3 == 4'hf ? _GEN_2826 : _GEN_3594; // @[executor.scala 466:52]
  wire [7:0] _GEN_3853 = opcode_3 == 4'hf ? _GEN_2827 : _GEN_3595; // @[executor.scala 466:52]
  wire [7:0] _GEN_3854 = opcode_3 == 4'hf ? _GEN_2828 : _GEN_3596; // @[executor.scala 466:52]
  wire [7:0] _GEN_3855 = opcode_3 == 4'hf ? _GEN_2829 : _GEN_3597; // @[executor.scala 466:52]
  wire [7:0] _GEN_3856 = opcode_3 == 4'hf ? _GEN_2830 : _GEN_3598; // @[executor.scala 466:52]
  wire [7:0] _GEN_3857 = opcode_3 == 4'hf ? _GEN_2831 : _GEN_3599; // @[executor.scala 466:52]
  wire [7:0] _GEN_3858 = opcode_3 == 4'hf ? _GEN_2832 : _GEN_3600; // @[executor.scala 466:52]
  wire [7:0] _GEN_3859 = opcode_3 == 4'hf ? _GEN_2833 : _GEN_3601; // @[executor.scala 466:52]
  wire [7:0] _GEN_3860 = opcode_3 == 4'hf ? _GEN_2834 : _GEN_3602; // @[executor.scala 466:52]
  wire [7:0] _GEN_3861 = opcode_3 == 4'hf ? _GEN_2835 : _GEN_3603; // @[executor.scala 466:52]
  wire [7:0] _GEN_3862 = opcode_3 == 4'hf ? _GEN_2836 : _GEN_3604; // @[executor.scala 466:52]
  wire [7:0] _GEN_3863 = opcode_3 == 4'hf ? _GEN_2837 : _GEN_3605; // @[executor.scala 466:52]
  wire [7:0] _GEN_3864 = opcode_3 == 4'hf ? _GEN_2838 : _GEN_3606; // @[executor.scala 466:52]
  wire [7:0] _GEN_3865 = opcode_3 == 4'hf ? _GEN_2839 : _GEN_3607; // @[executor.scala 466:52]
  wire [7:0] _GEN_3866 = opcode_3 == 4'hf ? _GEN_2840 : _GEN_3608; // @[executor.scala 466:52]
  wire [7:0] _GEN_3867 = opcode_3 == 4'hf ? _GEN_2841 : _GEN_3609; // @[executor.scala 466:52]
  wire [7:0] _GEN_3868 = opcode_3 == 4'hf ? _GEN_2842 : _GEN_3610; // @[executor.scala 466:52]
  wire [7:0] _GEN_3869 = opcode_3 == 4'hf ? _GEN_2843 : _GEN_3611; // @[executor.scala 466:52]
  wire [7:0] _GEN_3870 = opcode_3 == 4'hf ? _GEN_2844 : _GEN_3612; // @[executor.scala 466:52]
  wire [7:0] _GEN_3871 = opcode_3 == 4'hf ? _GEN_2845 : _GEN_3613; // @[executor.scala 466:52]
  wire [7:0] _GEN_3872 = opcode_3 == 4'hf ? _GEN_2846 : _GEN_3614; // @[executor.scala 466:52]
  wire [7:0] _GEN_3873 = opcode_3 == 4'hf ? _GEN_2847 : _GEN_3615; // @[executor.scala 466:52]
  wire [7:0] _GEN_3874 = opcode_3 == 4'hf ? _GEN_2848 : _GEN_3616; // @[executor.scala 466:52]
  wire [7:0] _GEN_3875 = opcode_3 == 4'hf ? _GEN_2849 : _GEN_3617; // @[executor.scala 466:52]
  wire [7:0] _GEN_3876 = opcode_3 == 4'hf ? _GEN_2850 : _GEN_3618; // @[executor.scala 466:52]
  wire [7:0] _GEN_3877 = opcode_3 == 4'hf ? _GEN_2851 : _GEN_3619; // @[executor.scala 466:52]
  wire [7:0] _GEN_3878 = opcode_3 == 4'hf ? _GEN_2852 : _GEN_3620; // @[executor.scala 466:52]
  wire [7:0] _GEN_3879 = opcode_3 == 4'hf ? _GEN_2853 : _GEN_3621; // @[executor.scala 466:52]
  wire [7:0] _GEN_3880 = opcode_3 == 4'hf ? _GEN_2854 : _GEN_3622; // @[executor.scala 466:52]
  wire [7:0] _GEN_3881 = opcode_3 == 4'hf ? _GEN_2855 : _GEN_3623; // @[executor.scala 466:52]
  wire [7:0] _GEN_3882 = opcode_3 == 4'hf ? _GEN_2856 : _GEN_3624; // @[executor.scala 466:52]
  wire [7:0] _GEN_3883 = opcode_3 == 4'hf ? _GEN_2857 : _GEN_3625; // @[executor.scala 466:52]
  wire [7:0] _GEN_3884 = opcode_3 == 4'hf ? _GEN_2858 : _GEN_3626; // @[executor.scala 466:52]
  wire [7:0] _GEN_3885 = opcode_3 == 4'hf ? _GEN_2859 : _GEN_3627; // @[executor.scala 466:52]
  wire [7:0] _GEN_3886 = opcode_3 == 4'hf ? _GEN_2860 : _GEN_3628; // @[executor.scala 466:52]
  wire [7:0] _GEN_3887 = opcode_3 == 4'hf ? _GEN_2861 : _GEN_3629; // @[executor.scala 466:52]
  wire [7:0] _GEN_3888 = opcode_3 == 4'hf ? _GEN_2862 : _GEN_3630; // @[executor.scala 466:52]
  wire [7:0] _GEN_3889 = opcode_3 == 4'hf ? _GEN_2863 : _GEN_3631; // @[executor.scala 466:52]
  wire [7:0] _GEN_3890 = opcode_3 == 4'hf ? _GEN_2864 : _GEN_3632; // @[executor.scala 466:52]
  wire [7:0] _GEN_3891 = opcode_3 == 4'hf ? _GEN_2865 : _GEN_3633; // @[executor.scala 466:52]
  wire [7:0] _GEN_3892 = opcode_3 == 4'hf ? _GEN_2866 : _GEN_3634; // @[executor.scala 466:52]
  wire [7:0] _GEN_3893 = opcode_3 == 4'hf ? _GEN_2867 : _GEN_3635; // @[executor.scala 466:52]
  wire [7:0] _GEN_3894 = opcode_3 == 4'hf ? _GEN_2868 : _GEN_3636; // @[executor.scala 466:52]
  wire [7:0] _GEN_3895 = opcode_3 == 4'hf ? _GEN_2869 : _GEN_3637; // @[executor.scala 466:52]
  wire [7:0] _GEN_3896 = opcode_3 == 4'hf ? _GEN_2870 : _GEN_3638; // @[executor.scala 466:52]
  wire [7:0] _GEN_3897 = opcode_3 == 4'hf ? _GEN_2871 : _GEN_3639; // @[executor.scala 466:52]
  wire [7:0] _GEN_3898 = opcode_3 == 4'hf ? _GEN_2872 : _GEN_3640; // @[executor.scala 466:52]
  wire [7:0] _GEN_3899 = opcode_3 == 4'hf ? _GEN_2873 : _GEN_3641; // @[executor.scala 466:52]
  wire [7:0] _GEN_3900 = opcode_3 == 4'hf ? _GEN_2874 : _GEN_3642; // @[executor.scala 466:52]
  wire [7:0] _GEN_3901 = opcode_3 == 4'hf ? _GEN_2875 : _GEN_3643; // @[executor.scala 466:52]
  wire [7:0] _GEN_3902 = opcode_3 == 4'hf ? _GEN_2876 : _GEN_3644; // @[executor.scala 466:52]
  wire [7:0] _GEN_3903 = opcode_3 == 4'hf ? _GEN_2877 : _GEN_3645; // @[executor.scala 466:52]
  wire [7:0] _GEN_3904 = opcode_3 == 4'hf ? _GEN_2878 : _GEN_3646; // @[executor.scala 466:52]
  wire [7:0] _GEN_3905 = opcode_3 == 4'hf ? _GEN_2879 : _GEN_3647; // @[executor.scala 466:52]
  wire [7:0] _GEN_3906 = opcode_3 == 4'hf ? _GEN_2880 : _GEN_3648; // @[executor.scala 466:52]
  wire [7:0] _GEN_3907 = opcode_3 == 4'hf ? _GEN_2881 : _GEN_3649; // @[executor.scala 466:52]
  wire [7:0] _GEN_3908 = opcode_3 == 4'hf ? _GEN_2882 : _GEN_3650; // @[executor.scala 466:52]
  wire [7:0] _GEN_3909 = opcode_3 == 4'hf ? _GEN_2883 : _GEN_3651; // @[executor.scala 466:52]
  wire [7:0] _GEN_3910 = opcode_3 == 4'hf ? _GEN_2884 : _GEN_3652; // @[executor.scala 466:52]
  wire [7:0] _GEN_3911 = opcode_3 == 4'hf ? _GEN_2885 : _GEN_3653; // @[executor.scala 466:52]
  wire [7:0] _GEN_3912 = opcode_3 == 4'hf ? _GEN_2886 : _GEN_3654; // @[executor.scala 466:52]
  wire [7:0] _GEN_3913 = opcode_3 == 4'hf ? _GEN_2887 : _GEN_3655; // @[executor.scala 466:52]
  wire [7:0] _GEN_3914 = opcode_3 == 4'hf ? _GEN_2888 : _GEN_3656; // @[executor.scala 466:52]
  wire [7:0] _GEN_3915 = opcode_3 == 4'hf ? _GEN_2889 : _GEN_3657; // @[executor.scala 466:52]
  wire [7:0] _GEN_3916 = opcode_3 == 4'hf ? _GEN_2890 : _GEN_3658; // @[executor.scala 466:52]
  wire [7:0] _GEN_3917 = opcode_3 == 4'hf ? _GEN_2891 : _GEN_3659; // @[executor.scala 466:52]
  wire [7:0] _GEN_3918 = opcode_3 == 4'hf ? _GEN_2892 : _GEN_3660; // @[executor.scala 466:52]
  wire [7:0] _GEN_3919 = opcode_3 == 4'hf ? _GEN_2893 : _GEN_3661; // @[executor.scala 466:52]
  wire [7:0] _GEN_3920 = opcode_3 == 4'hf ? _GEN_2894 : _GEN_3662; // @[executor.scala 466:52]
  wire [7:0] _GEN_3921 = opcode_3 == 4'hf ? _GEN_2895 : _GEN_3663; // @[executor.scala 466:52]
  wire [7:0] _GEN_3922 = opcode_3 == 4'hf ? _GEN_2896 : _GEN_3664; // @[executor.scala 466:52]
  wire [7:0] _GEN_3923 = opcode_3 == 4'hf ? _GEN_2897 : _GEN_3665; // @[executor.scala 466:52]
  wire [7:0] _GEN_3924 = opcode_3 == 4'hf ? _GEN_2898 : _GEN_3666; // @[executor.scala 466:52]
  wire [7:0] _GEN_3925 = opcode_3 == 4'hf ? _GEN_2899 : _GEN_3667; // @[executor.scala 466:52]
  wire [7:0] _GEN_3926 = opcode_3 == 4'hf ? _GEN_2900 : _GEN_3668; // @[executor.scala 466:52]
  wire [7:0] _GEN_3927 = opcode_3 == 4'hf ? _GEN_2901 : _GEN_3669; // @[executor.scala 466:52]
  wire [7:0] _GEN_3928 = opcode_3 == 4'hf ? _GEN_2902 : _GEN_3670; // @[executor.scala 466:52]
  wire [7:0] _GEN_3929 = opcode_3 == 4'hf ? _GEN_2903 : _GEN_3671; // @[executor.scala 466:52]
  wire [7:0] _GEN_3930 = opcode_3 == 4'hf ? _GEN_2904 : _GEN_3672; // @[executor.scala 466:52]
  wire [7:0] _GEN_3931 = opcode_3 == 4'hf ? _GEN_2905 : _GEN_3673; // @[executor.scala 466:52]
  wire [7:0] _GEN_3932 = opcode_3 == 4'hf ? _GEN_2906 : _GEN_3674; // @[executor.scala 466:52]
  wire [7:0] _GEN_3933 = opcode_3 == 4'hf ? _GEN_2907 : _GEN_3675; // @[executor.scala 466:52]
  wire [7:0] _GEN_3934 = opcode_3 == 4'hf ? _GEN_2908 : _GEN_3676; // @[executor.scala 466:52]
  wire [7:0] _GEN_3935 = opcode_3 == 4'hf ? _GEN_2909 : _GEN_3677; // @[executor.scala 466:52]
  wire [7:0] _GEN_3936 = opcode_3 == 4'hf ? _GEN_2910 : _GEN_3678; // @[executor.scala 466:52]
  wire [7:0] _GEN_3937 = opcode_3 == 4'hf ? _GEN_2911 : _GEN_3679; // @[executor.scala 466:52]
  wire [7:0] _GEN_3938 = opcode_3 == 4'hf ? _GEN_2912 : _GEN_3680; // @[executor.scala 466:52]
  wire [7:0] _GEN_3939 = opcode_3 == 4'hf ? _GEN_2913 : _GEN_3681; // @[executor.scala 466:52]
  wire [7:0] _GEN_3940 = opcode_3 == 4'hf ? _GEN_2914 : _GEN_3682; // @[executor.scala 466:52]
  wire [7:0] _GEN_3941 = opcode_3 == 4'hf ? _GEN_2915 : _GEN_3683; // @[executor.scala 466:52]
  wire [7:0] _GEN_3942 = opcode_3 == 4'hf ? _GEN_2916 : _GEN_3684; // @[executor.scala 466:52]
  wire [7:0] _GEN_3943 = opcode_3 == 4'hf ? _GEN_2917 : _GEN_3685; // @[executor.scala 466:52]
  wire [7:0] _GEN_3944 = opcode_3 == 4'hf ? _GEN_2918 : _GEN_3686; // @[executor.scala 466:52]
  wire [7:0] _GEN_3945 = opcode_3 == 4'hf ? _GEN_2919 : _GEN_3687; // @[executor.scala 466:52]
  wire [7:0] _GEN_3946 = opcode_3 == 4'hf ? _GEN_2920 : _GEN_3688; // @[executor.scala 466:52]
  wire [7:0] _GEN_3947 = opcode_3 == 4'hf ? _GEN_2921 : _GEN_3689; // @[executor.scala 466:52]
  wire [7:0] _GEN_3948 = opcode_3 == 4'hf ? _GEN_2922 : _GEN_3690; // @[executor.scala 466:52]
  wire [7:0] _GEN_3949 = opcode_3 == 4'hf ? _GEN_2923 : _GEN_3691; // @[executor.scala 466:52]
  wire [7:0] _GEN_3950 = opcode_3 == 4'hf ? _GEN_2924 : _GEN_3692; // @[executor.scala 466:52]
  wire [7:0] _GEN_3951 = opcode_3 == 4'hf ? _GEN_2925 : _GEN_3693; // @[executor.scala 466:52]
  wire [7:0] _GEN_3952 = opcode_3 == 4'hf ? _GEN_2926 : _GEN_3694; // @[executor.scala 466:52]
  wire [7:0] _GEN_3953 = opcode_3 == 4'hf ? _GEN_2927 : _GEN_3695; // @[executor.scala 466:52]
  wire [7:0] _GEN_3954 = opcode_3 == 4'hf ? _GEN_2928 : _GEN_3696; // @[executor.scala 466:52]
  wire [7:0] _GEN_3955 = opcode_3 == 4'hf ? _GEN_2929 : _GEN_3697; // @[executor.scala 466:52]
  wire [7:0] _GEN_3956 = opcode_3 == 4'hf ? _GEN_2930 : _GEN_3698; // @[executor.scala 466:52]
  wire [7:0] _GEN_3957 = opcode_3 == 4'hf ? _GEN_2931 : _GEN_3699; // @[executor.scala 466:52]
  wire [7:0] _GEN_3958 = opcode_3 == 4'hf ? _GEN_2932 : _GEN_3700; // @[executor.scala 466:52]
  wire [7:0] _GEN_3959 = opcode_3 == 4'hf ? _GEN_2933 : _GEN_3701; // @[executor.scala 466:52]
  wire [7:0] _GEN_3960 = opcode_3 == 4'hf ? _GEN_2934 : _GEN_3702; // @[executor.scala 466:52]
  wire [7:0] _GEN_3961 = opcode_3 == 4'hf ? _GEN_2935 : _GEN_3703; // @[executor.scala 466:52]
  wire [7:0] _GEN_3962 = opcode_3 == 4'hf ? _GEN_2936 : _GEN_3704; // @[executor.scala 466:52]
  wire [7:0] _GEN_3963 = opcode_3 == 4'hf ? _GEN_2937 : _GEN_3705; // @[executor.scala 466:52]
  wire [7:0] _GEN_3964 = opcode_3 == 4'hf ? _GEN_2938 : _GEN_3706; // @[executor.scala 466:52]
  wire [7:0] _GEN_3965 = opcode_3 == 4'hf ? _GEN_2939 : _GEN_3707; // @[executor.scala 466:52]
  wire [7:0] _GEN_3966 = opcode_3 == 4'hf ? _GEN_2940 : _GEN_3708; // @[executor.scala 466:52]
  wire [7:0] _GEN_3967 = opcode_3 == 4'hf ? _GEN_2941 : _GEN_3709; // @[executor.scala 466:52]
  wire [7:0] _GEN_3968 = opcode_3 == 4'hf ? _GEN_2942 : _GEN_3710; // @[executor.scala 466:52]
  wire [7:0] _GEN_3969 = opcode_3 == 4'hf ? _GEN_2943 : _GEN_3711; // @[executor.scala 466:52]
  wire [7:0] _GEN_3970 = opcode_3 == 4'hf ? _GEN_2944 : _GEN_3712; // @[executor.scala 466:52]
  wire [7:0] _GEN_3971 = opcode_3 == 4'hf ? _GEN_2945 : _GEN_3713; // @[executor.scala 466:52]
  wire [7:0] _GEN_3972 = opcode_3 == 4'hf ? _GEN_2946 : _GEN_3714; // @[executor.scala 466:52]
  wire [7:0] _GEN_3973 = opcode_3 == 4'hf ? _GEN_2947 : _GEN_3715; // @[executor.scala 466:52]
  wire [7:0] _GEN_3974 = opcode_3 == 4'hf ? _GEN_2948 : _GEN_3716; // @[executor.scala 466:52]
  wire [7:0] _GEN_3975 = opcode_3 == 4'hf ? _GEN_2949 : _GEN_3717; // @[executor.scala 466:52]
  wire [7:0] _GEN_3976 = opcode_3 == 4'hf ? _GEN_2950 : _GEN_3718; // @[executor.scala 466:52]
  wire [7:0] _GEN_3977 = opcode_3 == 4'hf ? _GEN_2951 : _GEN_3719; // @[executor.scala 466:52]
  wire [7:0] _GEN_3978 = opcode_3 == 4'hf ? _GEN_2952 : _GEN_3720; // @[executor.scala 466:52]
  wire [7:0] _GEN_3979 = opcode_3 == 4'hf ? _GEN_2953 : _GEN_3721; // @[executor.scala 466:52]
  wire [7:0] _GEN_3980 = opcode_3 == 4'hf ? _GEN_2954 : _GEN_3722; // @[executor.scala 466:52]
  wire [7:0] _GEN_3981 = opcode_3 == 4'hf ? _GEN_2955 : _GEN_3723; // @[executor.scala 466:52]
  wire [7:0] _GEN_3982 = opcode_3 == 4'hf ? _GEN_2956 : _GEN_3724; // @[executor.scala 466:52]
  wire [7:0] _GEN_3983 = opcode_3 == 4'hf ? _GEN_2957 : _GEN_3725; // @[executor.scala 466:52]
  wire [7:0] _GEN_3984 = opcode_3 == 4'hf ? _GEN_2958 : _GEN_3726; // @[executor.scala 466:52]
  wire [7:0] _GEN_3985 = opcode_3 == 4'hf ? _GEN_2959 : _GEN_3727; // @[executor.scala 466:52]
  wire [7:0] _GEN_3986 = opcode_3 == 4'hf ? _GEN_2960 : _GEN_3728; // @[executor.scala 466:52]
  wire [7:0] _GEN_3987 = opcode_3 == 4'hf ? _GEN_2961 : _GEN_3729; // @[executor.scala 466:52]
  wire [7:0] _GEN_3988 = opcode_3 == 4'hf ? _GEN_2962 : _GEN_3730; // @[executor.scala 466:52]
  wire [7:0] _GEN_3989 = opcode_3 == 4'hf ? _GEN_2963 : _GEN_3731; // @[executor.scala 466:52]
  wire [7:0] _GEN_3990 = opcode_3 == 4'hf ? _GEN_2964 : _GEN_3732; // @[executor.scala 466:52]
  wire [7:0] _GEN_3991 = opcode_3 == 4'hf ? _GEN_2965 : _GEN_3733; // @[executor.scala 466:52]
  wire [7:0] _GEN_3992 = opcode_3 == 4'hf ? _GEN_2966 : _GEN_3734; // @[executor.scala 466:52]
  wire [7:0] _GEN_3993 = opcode_3 == 4'hf ? _GEN_2967 : _GEN_3735; // @[executor.scala 466:52]
  wire [7:0] _GEN_3994 = opcode_3 == 4'hf ? _GEN_2968 : _GEN_3736; // @[executor.scala 466:52]
  wire [7:0] _GEN_3995 = opcode_3 == 4'hf ? _GEN_2969 : _GEN_3737; // @[executor.scala 466:52]
  wire [7:0] _GEN_3996 = opcode_3 == 4'hf ? _GEN_2970 : _GEN_3738; // @[executor.scala 466:52]
  wire [7:0] _GEN_3997 = opcode_3 == 4'hf ? _GEN_2971 : _GEN_3739; // @[executor.scala 466:52]
  wire [7:0] _GEN_3998 = opcode_3 == 4'hf ? _GEN_2972 : _GEN_3740; // @[executor.scala 466:52]
  wire [7:0] _GEN_3999 = opcode_3 == 4'hf ? _GEN_2973 : _GEN_3741; // @[executor.scala 466:52]
  wire [7:0] _GEN_4000 = opcode_3 == 4'hf ? _GEN_2974 : _GEN_3742; // @[executor.scala 466:52]
  wire [7:0] _GEN_4001 = opcode_3 == 4'hf ? _GEN_2975 : _GEN_3743; // @[executor.scala 466:52]
  wire [7:0] _GEN_4002 = opcode_3 == 4'hf ? _GEN_2976 : _GEN_3744; // @[executor.scala 466:52]
  wire [7:0] _GEN_4003 = opcode_3 == 4'hf ? _GEN_2977 : _GEN_3745; // @[executor.scala 466:52]
  wire [7:0] _GEN_4004 = opcode_3 == 4'hf ? _GEN_2978 : _GEN_3746; // @[executor.scala 466:52]
  wire [7:0] _GEN_4005 = opcode_3 == 4'hf ? _GEN_2979 : _GEN_3747; // @[executor.scala 466:52]
  wire [7:0] _GEN_4006 = opcode_3 == 4'hf ? _GEN_2980 : _GEN_3748; // @[executor.scala 466:52]
  wire [7:0] _GEN_4007 = opcode_3 == 4'hf ? _GEN_2981 : _GEN_3749; // @[executor.scala 466:52]
  wire [7:0] _GEN_4008 = opcode_3 == 4'hf ? _GEN_2982 : _GEN_3750; // @[executor.scala 466:52]
  wire [7:0] _GEN_4009 = opcode_3 == 4'hf ? _GEN_2983 : _GEN_3751; // @[executor.scala 466:52]
  wire [7:0] _GEN_4010 = opcode_3 == 4'hf ? _GEN_2984 : _GEN_3752; // @[executor.scala 466:52]
  wire [7:0] _GEN_4011 = opcode_3 == 4'hf ? _GEN_2985 : _GEN_3753; // @[executor.scala 466:52]
  wire [7:0] _GEN_4012 = opcode_3 == 4'hf ? _GEN_2986 : _GEN_3754; // @[executor.scala 466:52]
  wire [7:0] _GEN_4013 = opcode_3 == 4'hf ? _GEN_2987 : _GEN_3755; // @[executor.scala 466:52]
  wire [7:0] _GEN_4014 = opcode_3 == 4'hf ? _GEN_2988 : _GEN_3756; // @[executor.scala 466:52]
  wire [7:0] _GEN_4015 = opcode_3 == 4'hf ? _GEN_2989 : _GEN_3757; // @[executor.scala 466:52]
  wire [7:0] _GEN_4016 = opcode_3 == 4'hf ? _GEN_2990 : _GEN_3758; // @[executor.scala 466:52]
  wire [7:0] _GEN_4017 = opcode_3 == 4'hf ? _GEN_2991 : _GEN_3759; // @[executor.scala 466:52]
  wire [7:0] _GEN_4018 = opcode_3 == 4'hf ? _GEN_2992 : _GEN_3760; // @[executor.scala 466:52]
  wire [7:0] _GEN_4019 = opcode_3 == 4'hf ? _GEN_2993 : _GEN_3761; // @[executor.scala 466:52]
  wire [7:0] _GEN_4020 = opcode_3 == 4'hf ? _GEN_2994 : _GEN_3762; // @[executor.scala 466:52]
  wire [7:0] _GEN_4021 = opcode_3 == 4'hf ? _GEN_2995 : _GEN_3763; // @[executor.scala 466:52]
  wire [7:0] _GEN_4022 = opcode_3 == 4'hf ? _GEN_2996 : _GEN_3764; // @[executor.scala 466:52]
  wire [7:0] _GEN_4023 = opcode_3 == 4'hf ? _GEN_2997 : _GEN_3765; // @[executor.scala 466:52]
  wire [7:0] _GEN_4024 = opcode_3 == 4'hf ? _GEN_2998 : _GEN_3766; // @[executor.scala 466:52]
  wire [7:0] _GEN_4025 = opcode_3 == 4'hf ? _GEN_2999 : _GEN_3767; // @[executor.scala 466:52]
  wire [7:0] _GEN_4026 = opcode_3 == 4'hf ? _GEN_3000 : _GEN_3768; // @[executor.scala 466:52]
  wire [7:0] _GEN_4027 = opcode_3 == 4'hf ? _GEN_3001 : _GEN_3769; // @[executor.scala 466:52]
  wire [7:0] _GEN_4028 = opcode_3 == 4'hf ? _GEN_3002 : _GEN_3770; // @[executor.scala 466:52]
  wire [7:0] _GEN_4029 = opcode_3 == 4'hf ? _GEN_3003 : _GEN_3771; // @[executor.scala 466:52]
  wire [7:0] _GEN_4030 = opcode_3 == 4'hf ? _GEN_3004 : _GEN_3772; // @[executor.scala 466:52]
  wire [7:0] _GEN_4031 = opcode_3 == 4'hf ? _GEN_3005 : _GEN_3773; // @[executor.scala 466:52]
  wire [7:0] _GEN_4032 = opcode_3 == 4'hf ? _GEN_3006 : _GEN_3774; // @[executor.scala 466:52]
  wire [7:0] _GEN_4033 = opcode_3 == 4'hf ? _GEN_3007 : _GEN_3775; // @[executor.scala 466:52]
  wire [7:0] _GEN_4034 = opcode_3 == 4'hf ? _GEN_3008 : _GEN_3776; // @[executor.scala 466:52]
  wire [7:0] _GEN_4035 = opcode_3 == 4'hf ? _GEN_3009 : _GEN_3777; // @[executor.scala 466:52]
  wire [7:0] _GEN_4036 = opcode_3 == 4'hf ? _GEN_3010 : _GEN_3778; // @[executor.scala 466:52]
  wire [7:0] _GEN_4037 = opcode_3 == 4'hf ? _GEN_3011 : _GEN_3779; // @[executor.scala 466:52]
  wire [7:0] _GEN_4038 = opcode_3 == 4'hf ? _GEN_3012 : _GEN_3780; // @[executor.scala 466:52]
  wire [7:0] _GEN_4039 = opcode_3 == 4'hf ? _GEN_3013 : _GEN_3781; // @[executor.scala 466:52]
  wire [7:0] _GEN_4040 = opcode_3 == 4'hf ? _GEN_3014 : _GEN_3782; // @[executor.scala 466:52]
  wire [7:0] _GEN_4041 = opcode_3 == 4'hf ? _GEN_3015 : _GEN_3783; // @[executor.scala 466:52]
  wire [7:0] _GEN_4042 = opcode_3 == 4'hf ? _GEN_3016 : _GEN_3784; // @[executor.scala 466:52]
  wire [7:0] _GEN_4043 = opcode_3 == 4'hf ? _GEN_3017 : _GEN_3785; // @[executor.scala 466:52]
  wire [7:0] _GEN_4044 = opcode_3 == 4'hf ? _GEN_3018 : _GEN_3786; // @[executor.scala 466:52]
  wire [7:0] _GEN_4045 = opcode_3 == 4'hf ? _GEN_3019 : _GEN_3787; // @[executor.scala 466:52]
  wire [7:0] _GEN_4046 = opcode_3 == 4'hf ? _GEN_3020 : _GEN_3788; // @[executor.scala 466:52]
  wire [7:0] _GEN_4047 = opcode_3 == 4'hf ? _GEN_3021 : _GEN_3789; // @[executor.scala 466:52]
  wire [7:0] _GEN_4048 = opcode_3 == 4'hf ? _GEN_3022 : _GEN_3790; // @[executor.scala 466:52]
  wire [7:0] _GEN_4049 = opcode_3 == 4'hf ? _GEN_3023 : _GEN_3791; // @[executor.scala 466:52]
  wire [7:0] _GEN_4050 = opcode_3 == 4'hf ? _GEN_3024 : _GEN_3792; // @[executor.scala 466:52]
  wire [7:0] _GEN_4051 = opcode_3 == 4'hf ? _GEN_3025 : _GEN_3793; // @[executor.scala 466:52]
  wire [7:0] _GEN_4052 = opcode_3 == 4'hf ? _GEN_3026 : _GEN_3794; // @[executor.scala 466:52]
  wire [7:0] _GEN_4053 = opcode_3 == 4'hf ? _GEN_3027 : _GEN_3795; // @[executor.scala 466:52]
  wire [7:0] _GEN_4054 = opcode_3 == 4'hf ? _GEN_3028 : _GEN_3796; // @[executor.scala 466:52]
  wire [7:0] _GEN_4055 = opcode_3 == 4'hf ? _GEN_3029 : _GEN_3797; // @[executor.scala 466:52]
  wire [7:0] _GEN_4056 = opcode_3 == 4'hf ? _GEN_3030 : _GEN_3798; // @[executor.scala 466:52]
  wire [7:0] _GEN_4057 = opcode_3 == 4'hf ? _GEN_3031 : _GEN_3799; // @[executor.scala 466:52]
  wire [7:0] _GEN_4058 = opcode_3 == 4'hf ? _GEN_3032 : _GEN_3800; // @[executor.scala 466:52]
  wire [7:0] _GEN_4059 = opcode_3 == 4'hf ? _GEN_3033 : _GEN_3801; // @[executor.scala 466:52]
  wire [7:0] _GEN_4060 = opcode_3 == 4'hf ? _GEN_3034 : _GEN_3802; // @[executor.scala 466:52]
  wire [7:0] _GEN_4061 = opcode_3 == 4'hf ? _GEN_3035 : _GEN_3803; // @[executor.scala 466:52]
  wire [7:0] _GEN_4062 = opcode_3 == 4'hf ? _GEN_3036 : _GEN_3804; // @[executor.scala 466:52]
  wire [7:0] _GEN_4063 = opcode_3 == 4'hf ? _GEN_3037 : _GEN_3805; // @[executor.scala 466:52]
  wire [7:0] _GEN_4064 = opcode_3 == 4'hf ? _GEN_3038 : _GEN_3806; // @[executor.scala 466:52]
  wire [7:0] _GEN_4065 = opcode_3 == 4'hf ? _GEN_3039 : _GEN_3807; // @[executor.scala 466:52]
  wire [7:0] _GEN_4066 = opcode_3 == 4'hf ? _GEN_3040 : _GEN_3808; // @[executor.scala 466:52]
  wire [7:0] _GEN_4067 = opcode_3 == 4'hf ? _GEN_3041 : _GEN_3809; // @[executor.scala 466:52]
  wire [7:0] _GEN_4068 = opcode_3 == 4'hf ? _GEN_3042 : _GEN_3810; // @[executor.scala 466:52]
  wire [7:0] _GEN_4069 = opcode_3 == 4'hf ? _GEN_3043 : _GEN_3811; // @[executor.scala 466:52]
  wire [7:0] _GEN_4070 = opcode_3 == 4'hf ? _GEN_3044 : _GEN_3812; // @[executor.scala 466:52]
  wire [7:0] _GEN_4071 = opcode_3 == 4'hf ? _GEN_3045 : _GEN_3813; // @[executor.scala 466:52]
  wire [7:0] _GEN_4072 = opcode_3 == 4'hf ? _GEN_3046 : _GEN_3814; // @[executor.scala 466:52]
  wire [7:0] _GEN_4073 = opcode_3 == 4'hf ? _GEN_3047 : _GEN_3815; // @[executor.scala 466:52]
  wire [7:0] _GEN_4074 = opcode_3 == 4'hf ? _GEN_3048 : _GEN_3816; // @[executor.scala 466:52]
  wire [7:0] _GEN_4075 = opcode_3 == 4'hf ? _GEN_3049 : _GEN_3817; // @[executor.scala 466:52]
  wire [7:0] _GEN_4076 = opcode_3 == 4'hf ? _GEN_3050 : _GEN_3818; // @[executor.scala 466:52]
  wire [7:0] _GEN_4077 = opcode_3 == 4'hf ? _GEN_3051 : _GEN_3819; // @[executor.scala 466:52]
  wire [7:0] _GEN_4078 = opcode_3 == 4'hf ? _GEN_3052 : _GEN_3820; // @[executor.scala 466:52]
  wire [7:0] _GEN_4079 = opcode_3 == 4'hf ? _GEN_3053 : _GEN_3821; // @[executor.scala 466:52]
  wire [7:0] _GEN_4080 = opcode_3 == 4'hf ? _GEN_3054 : _GEN_3822; // @[executor.scala 466:52]
  wire [7:0] _GEN_4081 = opcode_3 == 4'hf ? _GEN_3055 : _GEN_3823; // @[executor.scala 466:52]
  wire [7:0] _GEN_4082 = opcode_3 == 4'hf ? _GEN_3056 : _GEN_3824; // @[executor.scala 466:52]
  wire [7:0] _GEN_4083 = opcode_3 == 4'hf ? _GEN_3057 : _GEN_3825; // @[executor.scala 466:52]
  wire [7:0] _GEN_4084 = opcode_3 == 4'hf ? _GEN_3058 : _GEN_3826; // @[executor.scala 466:52]
  wire [7:0] _GEN_4085 = opcode_3 == 4'hf ? _GEN_3059 : _GEN_3827; // @[executor.scala 466:52]
  wire [7:0] _GEN_4086 = opcode_3 == 4'hf ? _GEN_3060 : _GEN_3828; // @[executor.scala 466:52]
  wire [7:0] _GEN_4087 = opcode_3 == 4'hf ? _GEN_3061 : _GEN_3829; // @[executor.scala 466:52]
  wire [7:0] _GEN_4088 = opcode_3 == 4'hf ? _GEN_3062 : _GEN_3830; // @[executor.scala 466:52]
  wire [7:0] _GEN_4089 = opcode_3 == 4'hf ? _GEN_3063 : _GEN_3831; // @[executor.scala 466:52]
  wire [7:0] _GEN_4090 = opcode_3 == 4'hf ? _GEN_3064 : _GEN_3832; // @[executor.scala 466:52]
  wire [7:0] _GEN_4091 = opcode_3 == 4'hf ? _GEN_3065 : _GEN_3833; // @[executor.scala 466:52]
  wire [7:0] _GEN_4092 = opcode_3 == 4'hf ? _GEN_3066 : _GEN_3834; // @[executor.scala 466:52]
  wire [7:0] _GEN_4093 = opcode_3 == 4'hf ? _GEN_3067 : _GEN_3835; // @[executor.scala 466:52]
  wire [7:0] _GEN_4094 = opcode_3 == 4'hf ? _GEN_3068 : _GEN_3836; // @[executor.scala 466:52]
  wire [7:0] _GEN_4095 = opcode_3 == 4'hf ? _GEN_3069 : _GEN_3837; // @[executor.scala 466:52]
  wire [7:0] _GEN_4096 = opcode_3 == 4'hf ? _GEN_3070 : _GEN_3838; // @[executor.scala 466:52]
  wire [7:0] _GEN_4097 = opcode_3 == 4'hf ? _GEN_3071 : _GEN_3839; // @[executor.scala 466:52]
  wire [7:0] _GEN_4098 = opcode_3 == 4'hf ? _GEN_3072 : _GEN_3840; // @[executor.scala 466:52]
  wire [7:0] _GEN_4099 = opcode_3 == 4'hf ? _GEN_3073 : _GEN_3841; // @[executor.scala 466:52]
  wire [7:0] _GEN_4100 = opcode_3 == 4'hf ? _GEN_3074 : _GEN_3842; // @[executor.scala 466:52]
  wire [7:0] _GEN_4101 = opcode_3 == 4'hf ? _GEN_3075 : _GEN_3843; // @[executor.scala 466:52]
  wire [7:0] _GEN_4102 = opcode_3 == 4'hf ? _GEN_3076 : _GEN_3844; // @[executor.scala 466:52]
  wire [7:0] _GEN_4103 = opcode_3 == 4'hf ? _GEN_3077 : _GEN_3845; // @[executor.scala 466:52]
  assign io_pipe_phv_out_data_0 = phv_is_valid_processor ? _GEN_3851 : phv_data_0; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_1 = phv_is_valid_processor ? _GEN_3850 : phv_data_1; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_2 = phv_is_valid_processor ? _GEN_3849 : phv_data_2; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_3 = phv_is_valid_processor ? _GEN_3848 : phv_data_3; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_4 = phv_is_valid_processor ? _GEN_3855 : phv_data_4; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_5 = phv_is_valid_processor ? _GEN_3854 : phv_data_5; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_6 = phv_is_valid_processor ? _GEN_3853 : phv_data_6; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_7 = phv_is_valid_processor ? _GEN_3852 : phv_data_7; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_8 = phv_is_valid_processor ? _GEN_3859 : phv_data_8; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_9 = phv_is_valid_processor ? _GEN_3858 : phv_data_9; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_10 = phv_is_valid_processor ? _GEN_3857 : phv_data_10; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_11 = phv_is_valid_processor ? _GEN_3856 : phv_data_11; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_12 = phv_is_valid_processor ? _GEN_3863 : phv_data_12; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_13 = phv_is_valid_processor ? _GEN_3862 : phv_data_13; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_14 = phv_is_valid_processor ? _GEN_3861 : phv_data_14; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_15 = phv_is_valid_processor ? _GEN_3860 : phv_data_15; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_16 = phv_is_valid_processor ? _GEN_3867 : phv_data_16; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_17 = phv_is_valid_processor ? _GEN_3866 : phv_data_17; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_18 = phv_is_valid_processor ? _GEN_3865 : phv_data_18; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_19 = phv_is_valid_processor ? _GEN_3864 : phv_data_19; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_20 = phv_is_valid_processor ? _GEN_3871 : phv_data_20; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_21 = phv_is_valid_processor ? _GEN_3870 : phv_data_21; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_22 = phv_is_valid_processor ? _GEN_3869 : phv_data_22; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_23 = phv_is_valid_processor ? _GEN_3868 : phv_data_23; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_24 = phv_is_valid_processor ? _GEN_3875 : phv_data_24; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_25 = phv_is_valid_processor ? _GEN_3874 : phv_data_25; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_26 = phv_is_valid_processor ? _GEN_3873 : phv_data_26; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_27 = phv_is_valid_processor ? _GEN_3872 : phv_data_27; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_28 = phv_is_valid_processor ? _GEN_3879 : phv_data_28; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_29 = phv_is_valid_processor ? _GEN_3878 : phv_data_29; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_30 = phv_is_valid_processor ? _GEN_3877 : phv_data_30; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_31 = phv_is_valid_processor ? _GEN_3876 : phv_data_31; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_32 = phv_is_valid_processor ? _GEN_3883 : phv_data_32; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_33 = phv_is_valid_processor ? _GEN_3882 : phv_data_33; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_34 = phv_is_valid_processor ? _GEN_3881 : phv_data_34; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_35 = phv_is_valid_processor ? _GEN_3880 : phv_data_35; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_36 = phv_is_valid_processor ? _GEN_3887 : phv_data_36; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_37 = phv_is_valid_processor ? _GEN_3886 : phv_data_37; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_38 = phv_is_valid_processor ? _GEN_3885 : phv_data_38; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_39 = phv_is_valid_processor ? _GEN_3884 : phv_data_39; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_40 = phv_is_valid_processor ? _GEN_3891 : phv_data_40; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_41 = phv_is_valid_processor ? _GEN_3890 : phv_data_41; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_42 = phv_is_valid_processor ? _GEN_3889 : phv_data_42; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_43 = phv_is_valid_processor ? _GEN_3888 : phv_data_43; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_44 = phv_is_valid_processor ? _GEN_3895 : phv_data_44; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_45 = phv_is_valid_processor ? _GEN_3894 : phv_data_45; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_46 = phv_is_valid_processor ? _GEN_3893 : phv_data_46; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_47 = phv_is_valid_processor ? _GEN_3892 : phv_data_47; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_48 = phv_is_valid_processor ? _GEN_3899 : phv_data_48; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_49 = phv_is_valid_processor ? _GEN_3898 : phv_data_49; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_50 = phv_is_valid_processor ? _GEN_3897 : phv_data_50; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_51 = phv_is_valid_processor ? _GEN_3896 : phv_data_51; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_52 = phv_is_valid_processor ? _GEN_3903 : phv_data_52; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_53 = phv_is_valid_processor ? _GEN_3902 : phv_data_53; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_54 = phv_is_valid_processor ? _GEN_3901 : phv_data_54; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_55 = phv_is_valid_processor ? _GEN_3900 : phv_data_55; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_56 = phv_is_valid_processor ? _GEN_3907 : phv_data_56; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_57 = phv_is_valid_processor ? _GEN_3906 : phv_data_57; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_58 = phv_is_valid_processor ? _GEN_3905 : phv_data_58; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_59 = phv_is_valid_processor ? _GEN_3904 : phv_data_59; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_60 = phv_is_valid_processor ? _GEN_3911 : phv_data_60; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_61 = phv_is_valid_processor ? _GEN_3910 : phv_data_61; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_62 = phv_is_valid_processor ? _GEN_3909 : phv_data_62; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_63 = phv_is_valid_processor ? _GEN_3908 : phv_data_63; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_64 = phv_is_valid_processor ? _GEN_3915 : phv_data_64; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_65 = phv_is_valid_processor ? _GEN_3914 : phv_data_65; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_66 = phv_is_valid_processor ? _GEN_3913 : phv_data_66; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_67 = phv_is_valid_processor ? _GEN_3912 : phv_data_67; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_68 = phv_is_valid_processor ? _GEN_3919 : phv_data_68; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_69 = phv_is_valid_processor ? _GEN_3918 : phv_data_69; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_70 = phv_is_valid_processor ? _GEN_3917 : phv_data_70; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_71 = phv_is_valid_processor ? _GEN_3916 : phv_data_71; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_72 = phv_is_valid_processor ? _GEN_3923 : phv_data_72; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_73 = phv_is_valid_processor ? _GEN_3922 : phv_data_73; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_74 = phv_is_valid_processor ? _GEN_3921 : phv_data_74; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_75 = phv_is_valid_processor ? _GEN_3920 : phv_data_75; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_76 = phv_is_valid_processor ? _GEN_3927 : phv_data_76; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_77 = phv_is_valid_processor ? _GEN_3926 : phv_data_77; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_78 = phv_is_valid_processor ? _GEN_3925 : phv_data_78; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_79 = phv_is_valid_processor ? _GEN_3924 : phv_data_79; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_80 = phv_is_valid_processor ? _GEN_3931 : phv_data_80; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_81 = phv_is_valid_processor ? _GEN_3930 : phv_data_81; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_82 = phv_is_valid_processor ? _GEN_3929 : phv_data_82; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_83 = phv_is_valid_processor ? _GEN_3928 : phv_data_83; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_84 = phv_is_valid_processor ? _GEN_3935 : phv_data_84; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_85 = phv_is_valid_processor ? _GEN_3934 : phv_data_85; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_86 = phv_is_valid_processor ? _GEN_3933 : phv_data_86; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_87 = phv_is_valid_processor ? _GEN_3932 : phv_data_87; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_88 = phv_is_valid_processor ? _GEN_3939 : phv_data_88; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_89 = phv_is_valid_processor ? _GEN_3938 : phv_data_89; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_90 = phv_is_valid_processor ? _GEN_3937 : phv_data_90; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_91 = phv_is_valid_processor ? _GEN_3936 : phv_data_91; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_92 = phv_is_valid_processor ? _GEN_3943 : phv_data_92; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_93 = phv_is_valid_processor ? _GEN_3942 : phv_data_93; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_94 = phv_is_valid_processor ? _GEN_3941 : phv_data_94; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_95 = phv_is_valid_processor ? _GEN_3940 : phv_data_95; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_96 = phv_is_valid_processor ? _GEN_3947 : phv_data_96; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_97 = phv_is_valid_processor ? _GEN_3946 : phv_data_97; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_98 = phv_is_valid_processor ? _GEN_3945 : phv_data_98; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_99 = phv_is_valid_processor ? _GEN_3944 : phv_data_99; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_100 = phv_is_valid_processor ? _GEN_3951 : phv_data_100; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_101 = phv_is_valid_processor ? _GEN_3950 : phv_data_101; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_102 = phv_is_valid_processor ? _GEN_3949 : phv_data_102; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_103 = phv_is_valid_processor ? _GEN_3948 : phv_data_103; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_104 = phv_is_valid_processor ? _GEN_3955 : phv_data_104; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_105 = phv_is_valid_processor ? _GEN_3954 : phv_data_105; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_106 = phv_is_valid_processor ? _GEN_3953 : phv_data_106; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_107 = phv_is_valid_processor ? _GEN_3952 : phv_data_107; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_108 = phv_is_valid_processor ? _GEN_3959 : phv_data_108; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_109 = phv_is_valid_processor ? _GEN_3958 : phv_data_109; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_110 = phv_is_valid_processor ? _GEN_3957 : phv_data_110; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_111 = phv_is_valid_processor ? _GEN_3956 : phv_data_111; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_112 = phv_is_valid_processor ? _GEN_3963 : phv_data_112; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_113 = phv_is_valid_processor ? _GEN_3962 : phv_data_113; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_114 = phv_is_valid_processor ? _GEN_3961 : phv_data_114; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_115 = phv_is_valid_processor ? _GEN_3960 : phv_data_115; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_116 = phv_is_valid_processor ? _GEN_3967 : phv_data_116; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_117 = phv_is_valid_processor ? _GEN_3966 : phv_data_117; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_118 = phv_is_valid_processor ? _GEN_3965 : phv_data_118; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_119 = phv_is_valid_processor ? _GEN_3964 : phv_data_119; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_120 = phv_is_valid_processor ? _GEN_3971 : phv_data_120; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_121 = phv_is_valid_processor ? _GEN_3970 : phv_data_121; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_122 = phv_is_valid_processor ? _GEN_3969 : phv_data_122; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_123 = phv_is_valid_processor ? _GEN_3968 : phv_data_123; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_124 = phv_is_valid_processor ? _GEN_3975 : phv_data_124; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_125 = phv_is_valid_processor ? _GEN_3974 : phv_data_125; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_126 = phv_is_valid_processor ? _GEN_3973 : phv_data_126; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_127 = phv_is_valid_processor ? _GEN_3972 : phv_data_127; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_128 = phv_is_valid_processor ? _GEN_3979 : phv_data_128; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_129 = phv_is_valid_processor ? _GEN_3978 : phv_data_129; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_130 = phv_is_valid_processor ? _GEN_3977 : phv_data_130; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_131 = phv_is_valid_processor ? _GEN_3976 : phv_data_131; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_132 = phv_is_valid_processor ? _GEN_3983 : phv_data_132; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_133 = phv_is_valid_processor ? _GEN_3982 : phv_data_133; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_134 = phv_is_valid_processor ? _GEN_3981 : phv_data_134; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_135 = phv_is_valid_processor ? _GEN_3980 : phv_data_135; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_136 = phv_is_valid_processor ? _GEN_3987 : phv_data_136; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_137 = phv_is_valid_processor ? _GEN_3986 : phv_data_137; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_138 = phv_is_valid_processor ? _GEN_3985 : phv_data_138; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_139 = phv_is_valid_processor ? _GEN_3984 : phv_data_139; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_140 = phv_is_valid_processor ? _GEN_3991 : phv_data_140; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_141 = phv_is_valid_processor ? _GEN_3990 : phv_data_141; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_142 = phv_is_valid_processor ? _GEN_3989 : phv_data_142; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_143 = phv_is_valid_processor ? _GEN_3988 : phv_data_143; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_144 = phv_is_valid_processor ? _GEN_3995 : phv_data_144; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_145 = phv_is_valid_processor ? _GEN_3994 : phv_data_145; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_146 = phv_is_valid_processor ? _GEN_3993 : phv_data_146; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_147 = phv_is_valid_processor ? _GEN_3992 : phv_data_147; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_148 = phv_is_valid_processor ? _GEN_3999 : phv_data_148; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_149 = phv_is_valid_processor ? _GEN_3998 : phv_data_149; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_150 = phv_is_valid_processor ? _GEN_3997 : phv_data_150; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_151 = phv_is_valid_processor ? _GEN_3996 : phv_data_151; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_152 = phv_is_valid_processor ? _GEN_4003 : phv_data_152; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_153 = phv_is_valid_processor ? _GEN_4002 : phv_data_153; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_154 = phv_is_valid_processor ? _GEN_4001 : phv_data_154; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_155 = phv_is_valid_processor ? _GEN_4000 : phv_data_155; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_156 = phv_is_valid_processor ? _GEN_4007 : phv_data_156; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_157 = phv_is_valid_processor ? _GEN_4006 : phv_data_157; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_158 = phv_is_valid_processor ? _GEN_4005 : phv_data_158; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_159 = phv_is_valid_processor ? _GEN_4004 : phv_data_159; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_160 = phv_is_valid_processor ? _GEN_4011 : phv_data_160; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_161 = phv_is_valid_processor ? _GEN_4010 : phv_data_161; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_162 = phv_is_valid_processor ? _GEN_4009 : phv_data_162; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_163 = phv_is_valid_processor ? _GEN_4008 : phv_data_163; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_164 = phv_is_valid_processor ? _GEN_4015 : phv_data_164; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_165 = phv_is_valid_processor ? _GEN_4014 : phv_data_165; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_166 = phv_is_valid_processor ? _GEN_4013 : phv_data_166; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_167 = phv_is_valid_processor ? _GEN_4012 : phv_data_167; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_168 = phv_is_valid_processor ? _GEN_4019 : phv_data_168; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_169 = phv_is_valid_processor ? _GEN_4018 : phv_data_169; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_170 = phv_is_valid_processor ? _GEN_4017 : phv_data_170; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_171 = phv_is_valid_processor ? _GEN_4016 : phv_data_171; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_172 = phv_is_valid_processor ? _GEN_4023 : phv_data_172; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_173 = phv_is_valid_processor ? _GEN_4022 : phv_data_173; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_174 = phv_is_valid_processor ? _GEN_4021 : phv_data_174; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_175 = phv_is_valid_processor ? _GEN_4020 : phv_data_175; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_176 = phv_is_valid_processor ? _GEN_4027 : phv_data_176; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_177 = phv_is_valid_processor ? _GEN_4026 : phv_data_177; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_178 = phv_is_valid_processor ? _GEN_4025 : phv_data_178; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_179 = phv_is_valid_processor ? _GEN_4024 : phv_data_179; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_180 = phv_is_valid_processor ? _GEN_4031 : phv_data_180; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_181 = phv_is_valid_processor ? _GEN_4030 : phv_data_181; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_182 = phv_is_valid_processor ? _GEN_4029 : phv_data_182; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_183 = phv_is_valid_processor ? _GEN_4028 : phv_data_183; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_184 = phv_is_valid_processor ? _GEN_4035 : phv_data_184; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_185 = phv_is_valid_processor ? _GEN_4034 : phv_data_185; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_186 = phv_is_valid_processor ? _GEN_4033 : phv_data_186; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_187 = phv_is_valid_processor ? _GEN_4032 : phv_data_187; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_188 = phv_is_valid_processor ? _GEN_4039 : phv_data_188; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_189 = phv_is_valid_processor ? _GEN_4038 : phv_data_189; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_190 = phv_is_valid_processor ? _GEN_4037 : phv_data_190; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_191 = phv_is_valid_processor ? _GEN_4036 : phv_data_191; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_192 = phv_is_valid_processor ? _GEN_4043 : phv_data_192; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_193 = phv_is_valid_processor ? _GEN_4042 : phv_data_193; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_194 = phv_is_valid_processor ? _GEN_4041 : phv_data_194; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_195 = phv_is_valid_processor ? _GEN_4040 : phv_data_195; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_196 = phv_is_valid_processor ? _GEN_4047 : phv_data_196; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_197 = phv_is_valid_processor ? _GEN_4046 : phv_data_197; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_198 = phv_is_valid_processor ? _GEN_4045 : phv_data_198; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_199 = phv_is_valid_processor ? _GEN_4044 : phv_data_199; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_200 = phv_is_valid_processor ? _GEN_4051 : phv_data_200; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_201 = phv_is_valid_processor ? _GEN_4050 : phv_data_201; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_202 = phv_is_valid_processor ? _GEN_4049 : phv_data_202; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_203 = phv_is_valid_processor ? _GEN_4048 : phv_data_203; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_204 = phv_is_valid_processor ? _GEN_4055 : phv_data_204; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_205 = phv_is_valid_processor ? _GEN_4054 : phv_data_205; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_206 = phv_is_valid_processor ? _GEN_4053 : phv_data_206; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_207 = phv_is_valid_processor ? _GEN_4052 : phv_data_207; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_208 = phv_is_valid_processor ? _GEN_4059 : phv_data_208; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_209 = phv_is_valid_processor ? _GEN_4058 : phv_data_209; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_210 = phv_is_valid_processor ? _GEN_4057 : phv_data_210; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_211 = phv_is_valid_processor ? _GEN_4056 : phv_data_211; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_212 = phv_is_valid_processor ? _GEN_4063 : phv_data_212; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_213 = phv_is_valid_processor ? _GEN_4062 : phv_data_213; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_214 = phv_is_valid_processor ? _GEN_4061 : phv_data_214; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_215 = phv_is_valid_processor ? _GEN_4060 : phv_data_215; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_216 = phv_is_valid_processor ? _GEN_4067 : phv_data_216; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_217 = phv_is_valid_processor ? _GEN_4066 : phv_data_217; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_218 = phv_is_valid_processor ? _GEN_4065 : phv_data_218; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_219 = phv_is_valid_processor ? _GEN_4064 : phv_data_219; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_220 = phv_is_valid_processor ? _GEN_4071 : phv_data_220; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_221 = phv_is_valid_processor ? _GEN_4070 : phv_data_221; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_222 = phv_is_valid_processor ? _GEN_4069 : phv_data_222; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_223 = phv_is_valid_processor ? _GEN_4068 : phv_data_223; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_224 = phv_is_valid_processor ? _GEN_4075 : phv_data_224; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_225 = phv_is_valid_processor ? _GEN_4074 : phv_data_225; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_226 = phv_is_valid_processor ? _GEN_4073 : phv_data_226; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_227 = phv_is_valid_processor ? _GEN_4072 : phv_data_227; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_228 = phv_is_valid_processor ? _GEN_4079 : phv_data_228; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_229 = phv_is_valid_processor ? _GEN_4078 : phv_data_229; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_230 = phv_is_valid_processor ? _GEN_4077 : phv_data_230; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_231 = phv_is_valid_processor ? _GEN_4076 : phv_data_231; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_232 = phv_is_valid_processor ? _GEN_4083 : phv_data_232; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_233 = phv_is_valid_processor ? _GEN_4082 : phv_data_233; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_234 = phv_is_valid_processor ? _GEN_4081 : phv_data_234; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_235 = phv_is_valid_processor ? _GEN_4080 : phv_data_235; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_236 = phv_is_valid_processor ? _GEN_4087 : phv_data_236; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_237 = phv_is_valid_processor ? _GEN_4086 : phv_data_237; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_238 = phv_is_valid_processor ? _GEN_4085 : phv_data_238; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_239 = phv_is_valid_processor ? _GEN_4084 : phv_data_239; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_240 = phv_is_valid_processor ? _GEN_4091 : phv_data_240; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_241 = phv_is_valid_processor ? _GEN_4090 : phv_data_241; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_242 = phv_is_valid_processor ? _GEN_4089 : phv_data_242; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_243 = phv_is_valid_processor ? _GEN_4088 : phv_data_243; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_244 = phv_is_valid_processor ? _GEN_4095 : phv_data_244; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_245 = phv_is_valid_processor ? _GEN_4094 : phv_data_245; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_246 = phv_is_valid_processor ? _GEN_4093 : phv_data_246; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_247 = phv_is_valid_processor ? _GEN_4092 : phv_data_247; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_248 = phv_is_valid_processor ? _GEN_4099 : phv_data_248; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_249 = phv_is_valid_processor ? _GEN_4098 : phv_data_249; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_250 = phv_is_valid_processor ? _GEN_4097 : phv_data_250; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_251 = phv_is_valid_processor ? _GEN_4096 : phv_data_251; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_252 = phv_is_valid_processor ? _GEN_4103 : phv_data_252; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_253 = phv_is_valid_processor ? _GEN_4102 : phv_data_253; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_254 = phv_is_valid_processor ? _GEN_4101 : phv_data_254; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_255 = phv_is_valid_processor ? _GEN_4100 : phv_data_255; // @[executor.scala 461:39 executor.scala 450:25]
  always @(posedge clock) begin
    phv_data_0 <= io_pipe_phv_in_data_0; // @[executor.scala 449:13]
    phv_data_1 <= io_pipe_phv_in_data_1; // @[executor.scala 449:13]
    phv_data_2 <= io_pipe_phv_in_data_2; // @[executor.scala 449:13]
    phv_data_3 <= io_pipe_phv_in_data_3; // @[executor.scala 449:13]
    phv_data_4 <= io_pipe_phv_in_data_4; // @[executor.scala 449:13]
    phv_data_5 <= io_pipe_phv_in_data_5; // @[executor.scala 449:13]
    phv_data_6 <= io_pipe_phv_in_data_6; // @[executor.scala 449:13]
    phv_data_7 <= io_pipe_phv_in_data_7; // @[executor.scala 449:13]
    phv_data_8 <= io_pipe_phv_in_data_8; // @[executor.scala 449:13]
    phv_data_9 <= io_pipe_phv_in_data_9; // @[executor.scala 449:13]
    phv_data_10 <= io_pipe_phv_in_data_10; // @[executor.scala 449:13]
    phv_data_11 <= io_pipe_phv_in_data_11; // @[executor.scala 449:13]
    phv_data_12 <= io_pipe_phv_in_data_12; // @[executor.scala 449:13]
    phv_data_13 <= io_pipe_phv_in_data_13; // @[executor.scala 449:13]
    phv_data_14 <= io_pipe_phv_in_data_14; // @[executor.scala 449:13]
    phv_data_15 <= io_pipe_phv_in_data_15; // @[executor.scala 449:13]
    phv_data_16 <= io_pipe_phv_in_data_16; // @[executor.scala 449:13]
    phv_data_17 <= io_pipe_phv_in_data_17; // @[executor.scala 449:13]
    phv_data_18 <= io_pipe_phv_in_data_18; // @[executor.scala 449:13]
    phv_data_19 <= io_pipe_phv_in_data_19; // @[executor.scala 449:13]
    phv_data_20 <= io_pipe_phv_in_data_20; // @[executor.scala 449:13]
    phv_data_21 <= io_pipe_phv_in_data_21; // @[executor.scala 449:13]
    phv_data_22 <= io_pipe_phv_in_data_22; // @[executor.scala 449:13]
    phv_data_23 <= io_pipe_phv_in_data_23; // @[executor.scala 449:13]
    phv_data_24 <= io_pipe_phv_in_data_24; // @[executor.scala 449:13]
    phv_data_25 <= io_pipe_phv_in_data_25; // @[executor.scala 449:13]
    phv_data_26 <= io_pipe_phv_in_data_26; // @[executor.scala 449:13]
    phv_data_27 <= io_pipe_phv_in_data_27; // @[executor.scala 449:13]
    phv_data_28 <= io_pipe_phv_in_data_28; // @[executor.scala 449:13]
    phv_data_29 <= io_pipe_phv_in_data_29; // @[executor.scala 449:13]
    phv_data_30 <= io_pipe_phv_in_data_30; // @[executor.scala 449:13]
    phv_data_31 <= io_pipe_phv_in_data_31; // @[executor.scala 449:13]
    phv_data_32 <= io_pipe_phv_in_data_32; // @[executor.scala 449:13]
    phv_data_33 <= io_pipe_phv_in_data_33; // @[executor.scala 449:13]
    phv_data_34 <= io_pipe_phv_in_data_34; // @[executor.scala 449:13]
    phv_data_35 <= io_pipe_phv_in_data_35; // @[executor.scala 449:13]
    phv_data_36 <= io_pipe_phv_in_data_36; // @[executor.scala 449:13]
    phv_data_37 <= io_pipe_phv_in_data_37; // @[executor.scala 449:13]
    phv_data_38 <= io_pipe_phv_in_data_38; // @[executor.scala 449:13]
    phv_data_39 <= io_pipe_phv_in_data_39; // @[executor.scala 449:13]
    phv_data_40 <= io_pipe_phv_in_data_40; // @[executor.scala 449:13]
    phv_data_41 <= io_pipe_phv_in_data_41; // @[executor.scala 449:13]
    phv_data_42 <= io_pipe_phv_in_data_42; // @[executor.scala 449:13]
    phv_data_43 <= io_pipe_phv_in_data_43; // @[executor.scala 449:13]
    phv_data_44 <= io_pipe_phv_in_data_44; // @[executor.scala 449:13]
    phv_data_45 <= io_pipe_phv_in_data_45; // @[executor.scala 449:13]
    phv_data_46 <= io_pipe_phv_in_data_46; // @[executor.scala 449:13]
    phv_data_47 <= io_pipe_phv_in_data_47; // @[executor.scala 449:13]
    phv_data_48 <= io_pipe_phv_in_data_48; // @[executor.scala 449:13]
    phv_data_49 <= io_pipe_phv_in_data_49; // @[executor.scala 449:13]
    phv_data_50 <= io_pipe_phv_in_data_50; // @[executor.scala 449:13]
    phv_data_51 <= io_pipe_phv_in_data_51; // @[executor.scala 449:13]
    phv_data_52 <= io_pipe_phv_in_data_52; // @[executor.scala 449:13]
    phv_data_53 <= io_pipe_phv_in_data_53; // @[executor.scala 449:13]
    phv_data_54 <= io_pipe_phv_in_data_54; // @[executor.scala 449:13]
    phv_data_55 <= io_pipe_phv_in_data_55; // @[executor.scala 449:13]
    phv_data_56 <= io_pipe_phv_in_data_56; // @[executor.scala 449:13]
    phv_data_57 <= io_pipe_phv_in_data_57; // @[executor.scala 449:13]
    phv_data_58 <= io_pipe_phv_in_data_58; // @[executor.scala 449:13]
    phv_data_59 <= io_pipe_phv_in_data_59; // @[executor.scala 449:13]
    phv_data_60 <= io_pipe_phv_in_data_60; // @[executor.scala 449:13]
    phv_data_61 <= io_pipe_phv_in_data_61; // @[executor.scala 449:13]
    phv_data_62 <= io_pipe_phv_in_data_62; // @[executor.scala 449:13]
    phv_data_63 <= io_pipe_phv_in_data_63; // @[executor.scala 449:13]
    phv_data_64 <= io_pipe_phv_in_data_64; // @[executor.scala 449:13]
    phv_data_65 <= io_pipe_phv_in_data_65; // @[executor.scala 449:13]
    phv_data_66 <= io_pipe_phv_in_data_66; // @[executor.scala 449:13]
    phv_data_67 <= io_pipe_phv_in_data_67; // @[executor.scala 449:13]
    phv_data_68 <= io_pipe_phv_in_data_68; // @[executor.scala 449:13]
    phv_data_69 <= io_pipe_phv_in_data_69; // @[executor.scala 449:13]
    phv_data_70 <= io_pipe_phv_in_data_70; // @[executor.scala 449:13]
    phv_data_71 <= io_pipe_phv_in_data_71; // @[executor.scala 449:13]
    phv_data_72 <= io_pipe_phv_in_data_72; // @[executor.scala 449:13]
    phv_data_73 <= io_pipe_phv_in_data_73; // @[executor.scala 449:13]
    phv_data_74 <= io_pipe_phv_in_data_74; // @[executor.scala 449:13]
    phv_data_75 <= io_pipe_phv_in_data_75; // @[executor.scala 449:13]
    phv_data_76 <= io_pipe_phv_in_data_76; // @[executor.scala 449:13]
    phv_data_77 <= io_pipe_phv_in_data_77; // @[executor.scala 449:13]
    phv_data_78 <= io_pipe_phv_in_data_78; // @[executor.scala 449:13]
    phv_data_79 <= io_pipe_phv_in_data_79; // @[executor.scala 449:13]
    phv_data_80 <= io_pipe_phv_in_data_80; // @[executor.scala 449:13]
    phv_data_81 <= io_pipe_phv_in_data_81; // @[executor.scala 449:13]
    phv_data_82 <= io_pipe_phv_in_data_82; // @[executor.scala 449:13]
    phv_data_83 <= io_pipe_phv_in_data_83; // @[executor.scala 449:13]
    phv_data_84 <= io_pipe_phv_in_data_84; // @[executor.scala 449:13]
    phv_data_85 <= io_pipe_phv_in_data_85; // @[executor.scala 449:13]
    phv_data_86 <= io_pipe_phv_in_data_86; // @[executor.scala 449:13]
    phv_data_87 <= io_pipe_phv_in_data_87; // @[executor.scala 449:13]
    phv_data_88 <= io_pipe_phv_in_data_88; // @[executor.scala 449:13]
    phv_data_89 <= io_pipe_phv_in_data_89; // @[executor.scala 449:13]
    phv_data_90 <= io_pipe_phv_in_data_90; // @[executor.scala 449:13]
    phv_data_91 <= io_pipe_phv_in_data_91; // @[executor.scala 449:13]
    phv_data_92 <= io_pipe_phv_in_data_92; // @[executor.scala 449:13]
    phv_data_93 <= io_pipe_phv_in_data_93; // @[executor.scala 449:13]
    phv_data_94 <= io_pipe_phv_in_data_94; // @[executor.scala 449:13]
    phv_data_95 <= io_pipe_phv_in_data_95; // @[executor.scala 449:13]
    phv_data_96 <= io_pipe_phv_in_data_96; // @[executor.scala 449:13]
    phv_data_97 <= io_pipe_phv_in_data_97; // @[executor.scala 449:13]
    phv_data_98 <= io_pipe_phv_in_data_98; // @[executor.scala 449:13]
    phv_data_99 <= io_pipe_phv_in_data_99; // @[executor.scala 449:13]
    phv_data_100 <= io_pipe_phv_in_data_100; // @[executor.scala 449:13]
    phv_data_101 <= io_pipe_phv_in_data_101; // @[executor.scala 449:13]
    phv_data_102 <= io_pipe_phv_in_data_102; // @[executor.scala 449:13]
    phv_data_103 <= io_pipe_phv_in_data_103; // @[executor.scala 449:13]
    phv_data_104 <= io_pipe_phv_in_data_104; // @[executor.scala 449:13]
    phv_data_105 <= io_pipe_phv_in_data_105; // @[executor.scala 449:13]
    phv_data_106 <= io_pipe_phv_in_data_106; // @[executor.scala 449:13]
    phv_data_107 <= io_pipe_phv_in_data_107; // @[executor.scala 449:13]
    phv_data_108 <= io_pipe_phv_in_data_108; // @[executor.scala 449:13]
    phv_data_109 <= io_pipe_phv_in_data_109; // @[executor.scala 449:13]
    phv_data_110 <= io_pipe_phv_in_data_110; // @[executor.scala 449:13]
    phv_data_111 <= io_pipe_phv_in_data_111; // @[executor.scala 449:13]
    phv_data_112 <= io_pipe_phv_in_data_112; // @[executor.scala 449:13]
    phv_data_113 <= io_pipe_phv_in_data_113; // @[executor.scala 449:13]
    phv_data_114 <= io_pipe_phv_in_data_114; // @[executor.scala 449:13]
    phv_data_115 <= io_pipe_phv_in_data_115; // @[executor.scala 449:13]
    phv_data_116 <= io_pipe_phv_in_data_116; // @[executor.scala 449:13]
    phv_data_117 <= io_pipe_phv_in_data_117; // @[executor.scala 449:13]
    phv_data_118 <= io_pipe_phv_in_data_118; // @[executor.scala 449:13]
    phv_data_119 <= io_pipe_phv_in_data_119; // @[executor.scala 449:13]
    phv_data_120 <= io_pipe_phv_in_data_120; // @[executor.scala 449:13]
    phv_data_121 <= io_pipe_phv_in_data_121; // @[executor.scala 449:13]
    phv_data_122 <= io_pipe_phv_in_data_122; // @[executor.scala 449:13]
    phv_data_123 <= io_pipe_phv_in_data_123; // @[executor.scala 449:13]
    phv_data_124 <= io_pipe_phv_in_data_124; // @[executor.scala 449:13]
    phv_data_125 <= io_pipe_phv_in_data_125; // @[executor.scala 449:13]
    phv_data_126 <= io_pipe_phv_in_data_126; // @[executor.scala 449:13]
    phv_data_127 <= io_pipe_phv_in_data_127; // @[executor.scala 449:13]
    phv_data_128 <= io_pipe_phv_in_data_128; // @[executor.scala 449:13]
    phv_data_129 <= io_pipe_phv_in_data_129; // @[executor.scala 449:13]
    phv_data_130 <= io_pipe_phv_in_data_130; // @[executor.scala 449:13]
    phv_data_131 <= io_pipe_phv_in_data_131; // @[executor.scala 449:13]
    phv_data_132 <= io_pipe_phv_in_data_132; // @[executor.scala 449:13]
    phv_data_133 <= io_pipe_phv_in_data_133; // @[executor.scala 449:13]
    phv_data_134 <= io_pipe_phv_in_data_134; // @[executor.scala 449:13]
    phv_data_135 <= io_pipe_phv_in_data_135; // @[executor.scala 449:13]
    phv_data_136 <= io_pipe_phv_in_data_136; // @[executor.scala 449:13]
    phv_data_137 <= io_pipe_phv_in_data_137; // @[executor.scala 449:13]
    phv_data_138 <= io_pipe_phv_in_data_138; // @[executor.scala 449:13]
    phv_data_139 <= io_pipe_phv_in_data_139; // @[executor.scala 449:13]
    phv_data_140 <= io_pipe_phv_in_data_140; // @[executor.scala 449:13]
    phv_data_141 <= io_pipe_phv_in_data_141; // @[executor.scala 449:13]
    phv_data_142 <= io_pipe_phv_in_data_142; // @[executor.scala 449:13]
    phv_data_143 <= io_pipe_phv_in_data_143; // @[executor.scala 449:13]
    phv_data_144 <= io_pipe_phv_in_data_144; // @[executor.scala 449:13]
    phv_data_145 <= io_pipe_phv_in_data_145; // @[executor.scala 449:13]
    phv_data_146 <= io_pipe_phv_in_data_146; // @[executor.scala 449:13]
    phv_data_147 <= io_pipe_phv_in_data_147; // @[executor.scala 449:13]
    phv_data_148 <= io_pipe_phv_in_data_148; // @[executor.scala 449:13]
    phv_data_149 <= io_pipe_phv_in_data_149; // @[executor.scala 449:13]
    phv_data_150 <= io_pipe_phv_in_data_150; // @[executor.scala 449:13]
    phv_data_151 <= io_pipe_phv_in_data_151; // @[executor.scala 449:13]
    phv_data_152 <= io_pipe_phv_in_data_152; // @[executor.scala 449:13]
    phv_data_153 <= io_pipe_phv_in_data_153; // @[executor.scala 449:13]
    phv_data_154 <= io_pipe_phv_in_data_154; // @[executor.scala 449:13]
    phv_data_155 <= io_pipe_phv_in_data_155; // @[executor.scala 449:13]
    phv_data_156 <= io_pipe_phv_in_data_156; // @[executor.scala 449:13]
    phv_data_157 <= io_pipe_phv_in_data_157; // @[executor.scala 449:13]
    phv_data_158 <= io_pipe_phv_in_data_158; // @[executor.scala 449:13]
    phv_data_159 <= io_pipe_phv_in_data_159; // @[executor.scala 449:13]
    phv_data_160 <= io_pipe_phv_in_data_160; // @[executor.scala 449:13]
    phv_data_161 <= io_pipe_phv_in_data_161; // @[executor.scala 449:13]
    phv_data_162 <= io_pipe_phv_in_data_162; // @[executor.scala 449:13]
    phv_data_163 <= io_pipe_phv_in_data_163; // @[executor.scala 449:13]
    phv_data_164 <= io_pipe_phv_in_data_164; // @[executor.scala 449:13]
    phv_data_165 <= io_pipe_phv_in_data_165; // @[executor.scala 449:13]
    phv_data_166 <= io_pipe_phv_in_data_166; // @[executor.scala 449:13]
    phv_data_167 <= io_pipe_phv_in_data_167; // @[executor.scala 449:13]
    phv_data_168 <= io_pipe_phv_in_data_168; // @[executor.scala 449:13]
    phv_data_169 <= io_pipe_phv_in_data_169; // @[executor.scala 449:13]
    phv_data_170 <= io_pipe_phv_in_data_170; // @[executor.scala 449:13]
    phv_data_171 <= io_pipe_phv_in_data_171; // @[executor.scala 449:13]
    phv_data_172 <= io_pipe_phv_in_data_172; // @[executor.scala 449:13]
    phv_data_173 <= io_pipe_phv_in_data_173; // @[executor.scala 449:13]
    phv_data_174 <= io_pipe_phv_in_data_174; // @[executor.scala 449:13]
    phv_data_175 <= io_pipe_phv_in_data_175; // @[executor.scala 449:13]
    phv_data_176 <= io_pipe_phv_in_data_176; // @[executor.scala 449:13]
    phv_data_177 <= io_pipe_phv_in_data_177; // @[executor.scala 449:13]
    phv_data_178 <= io_pipe_phv_in_data_178; // @[executor.scala 449:13]
    phv_data_179 <= io_pipe_phv_in_data_179; // @[executor.scala 449:13]
    phv_data_180 <= io_pipe_phv_in_data_180; // @[executor.scala 449:13]
    phv_data_181 <= io_pipe_phv_in_data_181; // @[executor.scala 449:13]
    phv_data_182 <= io_pipe_phv_in_data_182; // @[executor.scala 449:13]
    phv_data_183 <= io_pipe_phv_in_data_183; // @[executor.scala 449:13]
    phv_data_184 <= io_pipe_phv_in_data_184; // @[executor.scala 449:13]
    phv_data_185 <= io_pipe_phv_in_data_185; // @[executor.scala 449:13]
    phv_data_186 <= io_pipe_phv_in_data_186; // @[executor.scala 449:13]
    phv_data_187 <= io_pipe_phv_in_data_187; // @[executor.scala 449:13]
    phv_data_188 <= io_pipe_phv_in_data_188; // @[executor.scala 449:13]
    phv_data_189 <= io_pipe_phv_in_data_189; // @[executor.scala 449:13]
    phv_data_190 <= io_pipe_phv_in_data_190; // @[executor.scala 449:13]
    phv_data_191 <= io_pipe_phv_in_data_191; // @[executor.scala 449:13]
    phv_data_192 <= io_pipe_phv_in_data_192; // @[executor.scala 449:13]
    phv_data_193 <= io_pipe_phv_in_data_193; // @[executor.scala 449:13]
    phv_data_194 <= io_pipe_phv_in_data_194; // @[executor.scala 449:13]
    phv_data_195 <= io_pipe_phv_in_data_195; // @[executor.scala 449:13]
    phv_data_196 <= io_pipe_phv_in_data_196; // @[executor.scala 449:13]
    phv_data_197 <= io_pipe_phv_in_data_197; // @[executor.scala 449:13]
    phv_data_198 <= io_pipe_phv_in_data_198; // @[executor.scala 449:13]
    phv_data_199 <= io_pipe_phv_in_data_199; // @[executor.scala 449:13]
    phv_data_200 <= io_pipe_phv_in_data_200; // @[executor.scala 449:13]
    phv_data_201 <= io_pipe_phv_in_data_201; // @[executor.scala 449:13]
    phv_data_202 <= io_pipe_phv_in_data_202; // @[executor.scala 449:13]
    phv_data_203 <= io_pipe_phv_in_data_203; // @[executor.scala 449:13]
    phv_data_204 <= io_pipe_phv_in_data_204; // @[executor.scala 449:13]
    phv_data_205 <= io_pipe_phv_in_data_205; // @[executor.scala 449:13]
    phv_data_206 <= io_pipe_phv_in_data_206; // @[executor.scala 449:13]
    phv_data_207 <= io_pipe_phv_in_data_207; // @[executor.scala 449:13]
    phv_data_208 <= io_pipe_phv_in_data_208; // @[executor.scala 449:13]
    phv_data_209 <= io_pipe_phv_in_data_209; // @[executor.scala 449:13]
    phv_data_210 <= io_pipe_phv_in_data_210; // @[executor.scala 449:13]
    phv_data_211 <= io_pipe_phv_in_data_211; // @[executor.scala 449:13]
    phv_data_212 <= io_pipe_phv_in_data_212; // @[executor.scala 449:13]
    phv_data_213 <= io_pipe_phv_in_data_213; // @[executor.scala 449:13]
    phv_data_214 <= io_pipe_phv_in_data_214; // @[executor.scala 449:13]
    phv_data_215 <= io_pipe_phv_in_data_215; // @[executor.scala 449:13]
    phv_data_216 <= io_pipe_phv_in_data_216; // @[executor.scala 449:13]
    phv_data_217 <= io_pipe_phv_in_data_217; // @[executor.scala 449:13]
    phv_data_218 <= io_pipe_phv_in_data_218; // @[executor.scala 449:13]
    phv_data_219 <= io_pipe_phv_in_data_219; // @[executor.scala 449:13]
    phv_data_220 <= io_pipe_phv_in_data_220; // @[executor.scala 449:13]
    phv_data_221 <= io_pipe_phv_in_data_221; // @[executor.scala 449:13]
    phv_data_222 <= io_pipe_phv_in_data_222; // @[executor.scala 449:13]
    phv_data_223 <= io_pipe_phv_in_data_223; // @[executor.scala 449:13]
    phv_data_224 <= io_pipe_phv_in_data_224; // @[executor.scala 449:13]
    phv_data_225 <= io_pipe_phv_in_data_225; // @[executor.scala 449:13]
    phv_data_226 <= io_pipe_phv_in_data_226; // @[executor.scala 449:13]
    phv_data_227 <= io_pipe_phv_in_data_227; // @[executor.scala 449:13]
    phv_data_228 <= io_pipe_phv_in_data_228; // @[executor.scala 449:13]
    phv_data_229 <= io_pipe_phv_in_data_229; // @[executor.scala 449:13]
    phv_data_230 <= io_pipe_phv_in_data_230; // @[executor.scala 449:13]
    phv_data_231 <= io_pipe_phv_in_data_231; // @[executor.scala 449:13]
    phv_data_232 <= io_pipe_phv_in_data_232; // @[executor.scala 449:13]
    phv_data_233 <= io_pipe_phv_in_data_233; // @[executor.scala 449:13]
    phv_data_234 <= io_pipe_phv_in_data_234; // @[executor.scala 449:13]
    phv_data_235 <= io_pipe_phv_in_data_235; // @[executor.scala 449:13]
    phv_data_236 <= io_pipe_phv_in_data_236; // @[executor.scala 449:13]
    phv_data_237 <= io_pipe_phv_in_data_237; // @[executor.scala 449:13]
    phv_data_238 <= io_pipe_phv_in_data_238; // @[executor.scala 449:13]
    phv_data_239 <= io_pipe_phv_in_data_239; // @[executor.scala 449:13]
    phv_data_240 <= io_pipe_phv_in_data_240; // @[executor.scala 449:13]
    phv_data_241 <= io_pipe_phv_in_data_241; // @[executor.scala 449:13]
    phv_data_242 <= io_pipe_phv_in_data_242; // @[executor.scala 449:13]
    phv_data_243 <= io_pipe_phv_in_data_243; // @[executor.scala 449:13]
    phv_data_244 <= io_pipe_phv_in_data_244; // @[executor.scala 449:13]
    phv_data_245 <= io_pipe_phv_in_data_245; // @[executor.scala 449:13]
    phv_data_246 <= io_pipe_phv_in_data_246; // @[executor.scala 449:13]
    phv_data_247 <= io_pipe_phv_in_data_247; // @[executor.scala 449:13]
    phv_data_248 <= io_pipe_phv_in_data_248; // @[executor.scala 449:13]
    phv_data_249 <= io_pipe_phv_in_data_249; // @[executor.scala 449:13]
    phv_data_250 <= io_pipe_phv_in_data_250; // @[executor.scala 449:13]
    phv_data_251 <= io_pipe_phv_in_data_251; // @[executor.scala 449:13]
    phv_data_252 <= io_pipe_phv_in_data_252; // @[executor.scala 449:13]
    phv_data_253 <= io_pipe_phv_in_data_253; // @[executor.scala 449:13]
    phv_data_254 <= io_pipe_phv_in_data_254; // @[executor.scala 449:13]
    phv_data_255 <= io_pipe_phv_in_data_255; // @[executor.scala 449:13]
    phv_is_valid_processor <= io_pipe_phv_in_is_valid_processor; // @[executor.scala 449:13]
    vliw_0 <= io_vliw_in_0; // @[executor.scala 453:14]
    vliw_1 <= io_vliw_in_1; // @[executor.scala 453:14]
    vliw_2 <= io_vliw_in_2; // @[executor.scala 453:14]
    vliw_3 <= io_vliw_in_3; // @[executor.scala 453:14]
    field_0 <= io_field_in_0; // @[executor.scala 455:15]
    field_1 <= io_field_in_1; // @[executor.scala 455:15]
    field_2 <= io_field_in_2; // @[executor.scala 455:15]
    field_3 <= io_field_in_3; // @[executor.scala 455:15]
    mask_0 <= io_mask_in_0; // @[executor.scala 457:14]
    mask_1 <= io_mask_in_1; // @[executor.scala 457:14]
    mask_2 <= io_mask_in_2; // @[executor.scala 457:14]
    mask_3 <= io_mask_in_3; // @[executor.scala 457:14]
    dst_offset_0 <= io_dst_offset_in_0; // @[executor.scala 459:20]
    dst_offset_1 <= io_dst_offset_in_1; // @[executor.scala 459:20]
    dst_offset_2 <= io_dst_offset_in_2; // @[executor.scala 459:20]
    dst_offset_3 <= io_dst_offset_in_3; // @[executor.scala 459:20]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  phv_data_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  phv_data_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  phv_data_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  phv_data_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  phv_data_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  phv_data_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  phv_data_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  phv_data_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  phv_data_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  phv_data_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  phv_data_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  phv_data_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  phv_data_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  phv_data_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  phv_data_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  phv_data_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  phv_data_16 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  phv_data_17 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  phv_data_18 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  phv_data_19 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  phv_data_20 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  phv_data_21 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  phv_data_22 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  phv_data_23 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  phv_data_24 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  phv_data_25 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  phv_data_26 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  phv_data_27 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  phv_data_28 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  phv_data_29 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  phv_data_30 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  phv_data_31 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  phv_data_32 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  phv_data_33 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  phv_data_34 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  phv_data_35 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  phv_data_36 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  phv_data_37 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  phv_data_38 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  phv_data_39 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  phv_data_40 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  phv_data_41 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  phv_data_42 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  phv_data_43 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  phv_data_44 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  phv_data_45 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  phv_data_46 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  phv_data_47 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  phv_data_48 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  phv_data_49 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  phv_data_50 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  phv_data_51 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  phv_data_52 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  phv_data_53 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  phv_data_54 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  phv_data_55 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  phv_data_56 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  phv_data_57 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  phv_data_58 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  phv_data_59 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  phv_data_60 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  phv_data_61 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  phv_data_62 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  phv_data_63 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  phv_data_64 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  phv_data_65 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  phv_data_66 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  phv_data_67 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  phv_data_68 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  phv_data_69 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  phv_data_70 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  phv_data_71 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  phv_data_72 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  phv_data_73 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  phv_data_74 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  phv_data_75 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  phv_data_76 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  phv_data_77 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  phv_data_78 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  phv_data_79 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  phv_data_80 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  phv_data_81 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  phv_data_82 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  phv_data_83 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  phv_data_84 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  phv_data_85 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  phv_data_86 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  phv_data_87 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  phv_data_88 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  phv_data_89 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  phv_data_90 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  phv_data_91 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  phv_data_92 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  phv_data_93 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  phv_data_94 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  phv_data_95 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  phv_data_96 = _RAND_96[7:0];
  _RAND_97 = {1{`RANDOM}};
  phv_data_97 = _RAND_97[7:0];
  _RAND_98 = {1{`RANDOM}};
  phv_data_98 = _RAND_98[7:0];
  _RAND_99 = {1{`RANDOM}};
  phv_data_99 = _RAND_99[7:0];
  _RAND_100 = {1{`RANDOM}};
  phv_data_100 = _RAND_100[7:0];
  _RAND_101 = {1{`RANDOM}};
  phv_data_101 = _RAND_101[7:0];
  _RAND_102 = {1{`RANDOM}};
  phv_data_102 = _RAND_102[7:0];
  _RAND_103 = {1{`RANDOM}};
  phv_data_103 = _RAND_103[7:0];
  _RAND_104 = {1{`RANDOM}};
  phv_data_104 = _RAND_104[7:0];
  _RAND_105 = {1{`RANDOM}};
  phv_data_105 = _RAND_105[7:0];
  _RAND_106 = {1{`RANDOM}};
  phv_data_106 = _RAND_106[7:0];
  _RAND_107 = {1{`RANDOM}};
  phv_data_107 = _RAND_107[7:0];
  _RAND_108 = {1{`RANDOM}};
  phv_data_108 = _RAND_108[7:0];
  _RAND_109 = {1{`RANDOM}};
  phv_data_109 = _RAND_109[7:0];
  _RAND_110 = {1{`RANDOM}};
  phv_data_110 = _RAND_110[7:0];
  _RAND_111 = {1{`RANDOM}};
  phv_data_111 = _RAND_111[7:0];
  _RAND_112 = {1{`RANDOM}};
  phv_data_112 = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  phv_data_113 = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  phv_data_114 = _RAND_114[7:0];
  _RAND_115 = {1{`RANDOM}};
  phv_data_115 = _RAND_115[7:0];
  _RAND_116 = {1{`RANDOM}};
  phv_data_116 = _RAND_116[7:0];
  _RAND_117 = {1{`RANDOM}};
  phv_data_117 = _RAND_117[7:0];
  _RAND_118 = {1{`RANDOM}};
  phv_data_118 = _RAND_118[7:0];
  _RAND_119 = {1{`RANDOM}};
  phv_data_119 = _RAND_119[7:0];
  _RAND_120 = {1{`RANDOM}};
  phv_data_120 = _RAND_120[7:0];
  _RAND_121 = {1{`RANDOM}};
  phv_data_121 = _RAND_121[7:0];
  _RAND_122 = {1{`RANDOM}};
  phv_data_122 = _RAND_122[7:0];
  _RAND_123 = {1{`RANDOM}};
  phv_data_123 = _RAND_123[7:0];
  _RAND_124 = {1{`RANDOM}};
  phv_data_124 = _RAND_124[7:0];
  _RAND_125 = {1{`RANDOM}};
  phv_data_125 = _RAND_125[7:0];
  _RAND_126 = {1{`RANDOM}};
  phv_data_126 = _RAND_126[7:0];
  _RAND_127 = {1{`RANDOM}};
  phv_data_127 = _RAND_127[7:0];
  _RAND_128 = {1{`RANDOM}};
  phv_data_128 = _RAND_128[7:0];
  _RAND_129 = {1{`RANDOM}};
  phv_data_129 = _RAND_129[7:0];
  _RAND_130 = {1{`RANDOM}};
  phv_data_130 = _RAND_130[7:0];
  _RAND_131 = {1{`RANDOM}};
  phv_data_131 = _RAND_131[7:0];
  _RAND_132 = {1{`RANDOM}};
  phv_data_132 = _RAND_132[7:0];
  _RAND_133 = {1{`RANDOM}};
  phv_data_133 = _RAND_133[7:0];
  _RAND_134 = {1{`RANDOM}};
  phv_data_134 = _RAND_134[7:0];
  _RAND_135 = {1{`RANDOM}};
  phv_data_135 = _RAND_135[7:0];
  _RAND_136 = {1{`RANDOM}};
  phv_data_136 = _RAND_136[7:0];
  _RAND_137 = {1{`RANDOM}};
  phv_data_137 = _RAND_137[7:0];
  _RAND_138 = {1{`RANDOM}};
  phv_data_138 = _RAND_138[7:0];
  _RAND_139 = {1{`RANDOM}};
  phv_data_139 = _RAND_139[7:0];
  _RAND_140 = {1{`RANDOM}};
  phv_data_140 = _RAND_140[7:0];
  _RAND_141 = {1{`RANDOM}};
  phv_data_141 = _RAND_141[7:0];
  _RAND_142 = {1{`RANDOM}};
  phv_data_142 = _RAND_142[7:0];
  _RAND_143 = {1{`RANDOM}};
  phv_data_143 = _RAND_143[7:0];
  _RAND_144 = {1{`RANDOM}};
  phv_data_144 = _RAND_144[7:0];
  _RAND_145 = {1{`RANDOM}};
  phv_data_145 = _RAND_145[7:0];
  _RAND_146 = {1{`RANDOM}};
  phv_data_146 = _RAND_146[7:0];
  _RAND_147 = {1{`RANDOM}};
  phv_data_147 = _RAND_147[7:0];
  _RAND_148 = {1{`RANDOM}};
  phv_data_148 = _RAND_148[7:0];
  _RAND_149 = {1{`RANDOM}};
  phv_data_149 = _RAND_149[7:0];
  _RAND_150 = {1{`RANDOM}};
  phv_data_150 = _RAND_150[7:0];
  _RAND_151 = {1{`RANDOM}};
  phv_data_151 = _RAND_151[7:0];
  _RAND_152 = {1{`RANDOM}};
  phv_data_152 = _RAND_152[7:0];
  _RAND_153 = {1{`RANDOM}};
  phv_data_153 = _RAND_153[7:0];
  _RAND_154 = {1{`RANDOM}};
  phv_data_154 = _RAND_154[7:0];
  _RAND_155 = {1{`RANDOM}};
  phv_data_155 = _RAND_155[7:0];
  _RAND_156 = {1{`RANDOM}};
  phv_data_156 = _RAND_156[7:0];
  _RAND_157 = {1{`RANDOM}};
  phv_data_157 = _RAND_157[7:0];
  _RAND_158 = {1{`RANDOM}};
  phv_data_158 = _RAND_158[7:0];
  _RAND_159 = {1{`RANDOM}};
  phv_data_159 = _RAND_159[7:0];
  _RAND_160 = {1{`RANDOM}};
  phv_data_160 = _RAND_160[7:0];
  _RAND_161 = {1{`RANDOM}};
  phv_data_161 = _RAND_161[7:0];
  _RAND_162 = {1{`RANDOM}};
  phv_data_162 = _RAND_162[7:0];
  _RAND_163 = {1{`RANDOM}};
  phv_data_163 = _RAND_163[7:0];
  _RAND_164 = {1{`RANDOM}};
  phv_data_164 = _RAND_164[7:0];
  _RAND_165 = {1{`RANDOM}};
  phv_data_165 = _RAND_165[7:0];
  _RAND_166 = {1{`RANDOM}};
  phv_data_166 = _RAND_166[7:0];
  _RAND_167 = {1{`RANDOM}};
  phv_data_167 = _RAND_167[7:0];
  _RAND_168 = {1{`RANDOM}};
  phv_data_168 = _RAND_168[7:0];
  _RAND_169 = {1{`RANDOM}};
  phv_data_169 = _RAND_169[7:0];
  _RAND_170 = {1{`RANDOM}};
  phv_data_170 = _RAND_170[7:0];
  _RAND_171 = {1{`RANDOM}};
  phv_data_171 = _RAND_171[7:0];
  _RAND_172 = {1{`RANDOM}};
  phv_data_172 = _RAND_172[7:0];
  _RAND_173 = {1{`RANDOM}};
  phv_data_173 = _RAND_173[7:0];
  _RAND_174 = {1{`RANDOM}};
  phv_data_174 = _RAND_174[7:0];
  _RAND_175 = {1{`RANDOM}};
  phv_data_175 = _RAND_175[7:0];
  _RAND_176 = {1{`RANDOM}};
  phv_data_176 = _RAND_176[7:0];
  _RAND_177 = {1{`RANDOM}};
  phv_data_177 = _RAND_177[7:0];
  _RAND_178 = {1{`RANDOM}};
  phv_data_178 = _RAND_178[7:0];
  _RAND_179 = {1{`RANDOM}};
  phv_data_179 = _RAND_179[7:0];
  _RAND_180 = {1{`RANDOM}};
  phv_data_180 = _RAND_180[7:0];
  _RAND_181 = {1{`RANDOM}};
  phv_data_181 = _RAND_181[7:0];
  _RAND_182 = {1{`RANDOM}};
  phv_data_182 = _RAND_182[7:0];
  _RAND_183 = {1{`RANDOM}};
  phv_data_183 = _RAND_183[7:0];
  _RAND_184 = {1{`RANDOM}};
  phv_data_184 = _RAND_184[7:0];
  _RAND_185 = {1{`RANDOM}};
  phv_data_185 = _RAND_185[7:0];
  _RAND_186 = {1{`RANDOM}};
  phv_data_186 = _RAND_186[7:0];
  _RAND_187 = {1{`RANDOM}};
  phv_data_187 = _RAND_187[7:0];
  _RAND_188 = {1{`RANDOM}};
  phv_data_188 = _RAND_188[7:0];
  _RAND_189 = {1{`RANDOM}};
  phv_data_189 = _RAND_189[7:0];
  _RAND_190 = {1{`RANDOM}};
  phv_data_190 = _RAND_190[7:0];
  _RAND_191 = {1{`RANDOM}};
  phv_data_191 = _RAND_191[7:0];
  _RAND_192 = {1{`RANDOM}};
  phv_data_192 = _RAND_192[7:0];
  _RAND_193 = {1{`RANDOM}};
  phv_data_193 = _RAND_193[7:0];
  _RAND_194 = {1{`RANDOM}};
  phv_data_194 = _RAND_194[7:0];
  _RAND_195 = {1{`RANDOM}};
  phv_data_195 = _RAND_195[7:0];
  _RAND_196 = {1{`RANDOM}};
  phv_data_196 = _RAND_196[7:0];
  _RAND_197 = {1{`RANDOM}};
  phv_data_197 = _RAND_197[7:0];
  _RAND_198 = {1{`RANDOM}};
  phv_data_198 = _RAND_198[7:0];
  _RAND_199 = {1{`RANDOM}};
  phv_data_199 = _RAND_199[7:0];
  _RAND_200 = {1{`RANDOM}};
  phv_data_200 = _RAND_200[7:0];
  _RAND_201 = {1{`RANDOM}};
  phv_data_201 = _RAND_201[7:0];
  _RAND_202 = {1{`RANDOM}};
  phv_data_202 = _RAND_202[7:0];
  _RAND_203 = {1{`RANDOM}};
  phv_data_203 = _RAND_203[7:0];
  _RAND_204 = {1{`RANDOM}};
  phv_data_204 = _RAND_204[7:0];
  _RAND_205 = {1{`RANDOM}};
  phv_data_205 = _RAND_205[7:0];
  _RAND_206 = {1{`RANDOM}};
  phv_data_206 = _RAND_206[7:0];
  _RAND_207 = {1{`RANDOM}};
  phv_data_207 = _RAND_207[7:0];
  _RAND_208 = {1{`RANDOM}};
  phv_data_208 = _RAND_208[7:0];
  _RAND_209 = {1{`RANDOM}};
  phv_data_209 = _RAND_209[7:0];
  _RAND_210 = {1{`RANDOM}};
  phv_data_210 = _RAND_210[7:0];
  _RAND_211 = {1{`RANDOM}};
  phv_data_211 = _RAND_211[7:0];
  _RAND_212 = {1{`RANDOM}};
  phv_data_212 = _RAND_212[7:0];
  _RAND_213 = {1{`RANDOM}};
  phv_data_213 = _RAND_213[7:0];
  _RAND_214 = {1{`RANDOM}};
  phv_data_214 = _RAND_214[7:0];
  _RAND_215 = {1{`RANDOM}};
  phv_data_215 = _RAND_215[7:0];
  _RAND_216 = {1{`RANDOM}};
  phv_data_216 = _RAND_216[7:0];
  _RAND_217 = {1{`RANDOM}};
  phv_data_217 = _RAND_217[7:0];
  _RAND_218 = {1{`RANDOM}};
  phv_data_218 = _RAND_218[7:0];
  _RAND_219 = {1{`RANDOM}};
  phv_data_219 = _RAND_219[7:0];
  _RAND_220 = {1{`RANDOM}};
  phv_data_220 = _RAND_220[7:0];
  _RAND_221 = {1{`RANDOM}};
  phv_data_221 = _RAND_221[7:0];
  _RAND_222 = {1{`RANDOM}};
  phv_data_222 = _RAND_222[7:0];
  _RAND_223 = {1{`RANDOM}};
  phv_data_223 = _RAND_223[7:0];
  _RAND_224 = {1{`RANDOM}};
  phv_data_224 = _RAND_224[7:0];
  _RAND_225 = {1{`RANDOM}};
  phv_data_225 = _RAND_225[7:0];
  _RAND_226 = {1{`RANDOM}};
  phv_data_226 = _RAND_226[7:0];
  _RAND_227 = {1{`RANDOM}};
  phv_data_227 = _RAND_227[7:0];
  _RAND_228 = {1{`RANDOM}};
  phv_data_228 = _RAND_228[7:0];
  _RAND_229 = {1{`RANDOM}};
  phv_data_229 = _RAND_229[7:0];
  _RAND_230 = {1{`RANDOM}};
  phv_data_230 = _RAND_230[7:0];
  _RAND_231 = {1{`RANDOM}};
  phv_data_231 = _RAND_231[7:0];
  _RAND_232 = {1{`RANDOM}};
  phv_data_232 = _RAND_232[7:0];
  _RAND_233 = {1{`RANDOM}};
  phv_data_233 = _RAND_233[7:0];
  _RAND_234 = {1{`RANDOM}};
  phv_data_234 = _RAND_234[7:0];
  _RAND_235 = {1{`RANDOM}};
  phv_data_235 = _RAND_235[7:0];
  _RAND_236 = {1{`RANDOM}};
  phv_data_236 = _RAND_236[7:0];
  _RAND_237 = {1{`RANDOM}};
  phv_data_237 = _RAND_237[7:0];
  _RAND_238 = {1{`RANDOM}};
  phv_data_238 = _RAND_238[7:0];
  _RAND_239 = {1{`RANDOM}};
  phv_data_239 = _RAND_239[7:0];
  _RAND_240 = {1{`RANDOM}};
  phv_data_240 = _RAND_240[7:0];
  _RAND_241 = {1{`RANDOM}};
  phv_data_241 = _RAND_241[7:0];
  _RAND_242 = {1{`RANDOM}};
  phv_data_242 = _RAND_242[7:0];
  _RAND_243 = {1{`RANDOM}};
  phv_data_243 = _RAND_243[7:0];
  _RAND_244 = {1{`RANDOM}};
  phv_data_244 = _RAND_244[7:0];
  _RAND_245 = {1{`RANDOM}};
  phv_data_245 = _RAND_245[7:0];
  _RAND_246 = {1{`RANDOM}};
  phv_data_246 = _RAND_246[7:0];
  _RAND_247 = {1{`RANDOM}};
  phv_data_247 = _RAND_247[7:0];
  _RAND_248 = {1{`RANDOM}};
  phv_data_248 = _RAND_248[7:0];
  _RAND_249 = {1{`RANDOM}};
  phv_data_249 = _RAND_249[7:0];
  _RAND_250 = {1{`RANDOM}};
  phv_data_250 = _RAND_250[7:0];
  _RAND_251 = {1{`RANDOM}};
  phv_data_251 = _RAND_251[7:0];
  _RAND_252 = {1{`RANDOM}};
  phv_data_252 = _RAND_252[7:0];
  _RAND_253 = {1{`RANDOM}};
  phv_data_253 = _RAND_253[7:0];
  _RAND_254 = {1{`RANDOM}};
  phv_data_254 = _RAND_254[7:0];
  _RAND_255 = {1{`RANDOM}};
  phv_data_255 = _RAND_255[7:0];
  _RAND_256 = {1{`RANDOM}};
  phv_is_valid_processor = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  vliw_0 = _RAND_257[31:0];
  _RAND_258 = {1{`RANDOM}};
  vliw_1 = _RAND_258[31:0];
  _RAND_259 = {1{`RANDOM}};
  vliw_2 = _RAND_259[31:0];
  _RAND_260 = {1{`RANDOM}};
  vliw_3 = _RAND_260[31:0];
  _RAND_261 = {1{`RANDOM}};
  field_0 = _RAND_261[31:0];
  _RAND_262 = {1{`RANDOM}};
  field_1 = _RAND_262[31:0];
  _RAND_263 = {1{`RANDOM}};
  field_2 = _RAND_263[31:0];
  _RAND_264 = {1{`RANDOM}};
  field_3 = _RAND_264[31:0];
  _RAND_265 = {1{`RANDOM}};
  mask_0 = _RAND_265[3:0];
  _RAND_266 = {1{`RANDOM}};
  mask_1 = _RAND_266[3:0];
  _RAND_267 = {1{`RANDOM}};
  mask_2 = _RAND_267[3:0];
  _RAND_268 = {1{`RANDOM}};
  mask_3 = _RAND_268[3:0];
  _RAND_269 = {1{`RANDOM}};
  dst_offset_0 = _RAND_269[5:0];
  _RAND_270 = {1{`RANDOM}};
  dst_offset_1 = _RAND_270[5:0];
  _RAND_271 = {1{`RANDOM}};
  dst_offset_2 = _RAND_271[5:0];
  _RAND_272 = {1{`RANDOM}};
  dst_offset_3 = _RAND_272[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
