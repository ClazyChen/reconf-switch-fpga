module ParserPISA(
  input         clock,
  input  [7:0]  io_pipe_phv_in_data_0,
  input  [7:0]  io_pipe_phv_in_data_1,
  input  [7:0]  io_pipe_phv_in_data_2,
  input  [7:0]  io_pipe_phv_in_data_3,
  input  [7:0]  io_pipe_phv_in_data_4,
  input  [7:0]  io_pipe_phv_in_data_5,
  input  [7:0]  io_pipe_phv_in_data_6,
  input  [7:0]  io_pipe_phv_in_data_7,
  input  [7:0]  io_pipe_phv_in_data_8,
  input  [7:0]  io_pipe_phv_in_data_9,
  input  [7:0]  io_pipe_phv_in_data_10,
  input  [7:0]  io_pipe_phv_in_data_11,
  input  [7:0]  io_pipe_phv_in_data_12,
  input  [7:0]  io_pipe_phv_in_data_13,
  input  [7:0]  io_pipe_phv_in_data_14,
  input  [7:0]  io_pipe_phv_in_data_15,
  input  [7:0]  io_pipe_phv_in_data_16,
  input  [7:0]  io_pipe_phv_in_data_17,
  input  [7:0]  io_pipe_phv_in_data_18,
  input  [7:0]  io_pipe_phv_in_data_19,
  input  [7:0]  io_pipe_phv_in_data_20,
  input  [7:0]  io_pipe_phv_in_data_21,
  input  [7:0]  io_pipe_phv_in_data_22,
  input  [7:0]  io_pipe_phv_in_data_23,
  input  [7:0]  io_pipe_phv_in_data_24,
  input  [7:0]  io_pipe_phv_in_data_25,
  input  [7:0]  io_pipe_phv_in_data_26,
  input  [7:0]  io_pipe_phv_in_data_27,
  input  [7:0]  io_pipe_phv_in_data_28,
  input  [7:0]  io_pipe_phv_in_data_29,
  input  [7:0]  io_pipe_phv_in_data_30,
  input  [7:0]  io_pipe_phv_in_data_31,
  input  [7:0]  io_pipe_phv_in_data_32,
  input  [7:0]  io_pipe_phv_in_data_33,
  input  [7:0]  io_pipe_phv_in_data_34,
  input  [7:0]  io_pipe_phv_in_data_35,
  input  [7:0]  io_pipe_phv_in_data_36,
  input  [7:0]  io_pipe_phv_in_data_37,
  input  [7:0]  io_pipe_phv_in_data_38,
  input  [7:0]  io_pipe_phv_in_data_39,
  input  [7:0]  io_pipe_phv_in_data_40,
  input  [7:0]  io_pipe_phv_in_data_41,
  input  [7:0]  io_pipe_phv_in_data_42,
  input  [7:0]  io_pipe_phv_in_data_43,
  input  [7:0]  io_pipe_phv_in_data_44,
  input  [7:0]  io_pipe_phv_in_data_45,
  input  [7:0]  io_pipe_phv_in_data_46,
  input  [7:0]  io_pipe_phv_in_data_47,
  input  [7:0]  io_pipe_phv_in_data_48,
  input  [7:0]  io_pipe_phv_in_data_49,
  input  [7:0]  io_pipe_phv_in_data_50,
  input  [7:0]  io_pipe_phv_in_data_51,
  input  [7:0]  io_pipe_phv_in_data_52,
  input  [7:0]  io_pipe_phv_in_data_53,
  input  [7:0]  io_pipe_phv_in_data_54,
  input  [7:0]  io_pipe_phv_in_data_55,
  input  [7:0]  io_pipe_phv_in_data_56,
  input  [7:0]  io_pipe_phv_in_data_57,
  input  [7:0]  io_pipe_phv_in_data_58,
  input  [7:0]  io_pipe_phv_in_data_59,
  input  [7:0]  io_pipe_phv_in_data_60,
  input  [7:0]  io_pipe_phv_in_data_61,
  input  [7:0]  io_pipe_phv_in_data_62,
  input  [7:0]  io_pipe_phv_in_data_63,
  input  [7:0]  io_pipe_phv_in_data_64,
  input  [7:0]  io_pipe_phv_in_data_65,
  input  [7:0]  io_pipe_phv_in_data_66,
  input  [7:0]  io_pipe_phv_in_data_67,
  input  [7:0]  io_pipe_phv_in_data_68,
  input  [7:0]  io_pipe_phv_in_data_69,
  input  [7:0]  io_pipe_phv_in_data_70,
  input  [7:0]  io_pipe_phv_in_data_71,
  input  [7:0]  io_pipe_phv_in_data_72,
  input  [7:0]  io_pipe_phv_in_data_73,
  input  [7:0]  io_pipe_phv_in_data_74,
  input  [7:0]  io_pipe_phv_in_data_75,
  input  [7:0]  io_pipe_phv_in_data_76,
  input  [7:0]  io_pipe_phv_in_data_77,
  input  [7:0]  io_pipe_phv_in_data_78,
  input  [7:0]  io_pipe_phv_in_data_79,
  input  [7:0]  io_pipe_phv_in_data_80,
  input  [7:0]  io_pipe_phv_in_data_81,
  input  [7:0]  io_pipe_phv_in_data_82,
  input  [7:0]  io_pipe_phv_in_data_83,
  input  [7:0]  io_pipe_phv_in_data_84,
  input  [7:0]  io_pipe_phv_in_data_85,
  input  [7:0]  io_pipe_phv_in_data_86,
  input  [7:0]  io_pipe_phv_in_data_87,
  input  [7:0]  io_pipe_phv_in_data_88,
  input  [7:0]  io_pipe_phv_in_data_89,
  input  [7:0]  io_pipe_phv_in_data_90,
  input  [7:0]  io_pipe_phv_in_data_91,
  input  [7:0]  io_pipe_phv_in_data_92,
  input  [7:0]  io_pipe_phv_in_data_93,
  input  [7:0]  io_pipe_phv_in_data_94,
  input  [7:0]  io_pipe_phv_in_data_95,
  input  [7:0]  io_pipe_phv_in_data_96,
  input  [7:0]  io_pipe_phv_in_data_97,
  input  [7:0]  io_pipe_phv_in_data_98,
  input  [7:0]  io_pipe_phv_in_data_99,
  input  [7:0]  io_pipe_phv_in_data_100,
  input  [7:0]  io_pipe_phv_in_data_101,
  input  [7:0]  io_pipe_phv_in_data_102,
  input  [7:0]  io_pipe_phv_in_data_103,
  input  [7:0]  io_pipe_phv_in_data_104,
  input  [7:0]  io_pipe_phv_in_data_105,
  input  [7:0]  io_pipe_phv_in_data_106,
  input  [7:0]  io_pipe_phv_in_data_107,
  input  [7:0]  io_pipe_phv_in_data_108,
  input  [7:0]  io_pipe_phv_in_data_109,
  input  [7:0]  io_pipe_phv_in_data_110,
  input  [7:0]  io_pipe_phv_in_data_111,
  input  [7:0]  io_pipe_phv_in_data_112,
  input  [7:0]  io_pipe_phv_in_data_113,
  input  [7:0]  io_pipe_phv_in_data_114,
  input  [7:0]  io_pipe_phv_in_data_115,
  input  [7:0]  io_pipe_phv_in_data_116,
  input  [7:0]  io_pipe_phv_in_data_117,
  input  [7:0]  io_pipe_phv_in_data_118,
  input  [7:0]  io_pipe_phv_in_data_119,
  input  [7:0]  io_pipe_phv_in_data_120,
  input  [7:0]  io_pipe_phv_in_data_121,
  input  [7:0]  io_pipe_phv_in_data_122,
  input  [7:0]  io_pipe_phv_in_data_123,
  input  [7:0]  io_pipe_phv_in_data_124,
  input  [7:0]  io_pipe_phv_in_data_125,
  input  [7:0]  io_pipe_phv_in_data_126,
  input  [7:0]  io_pipe_phv_in_data_127,
  input  [7:0]  io_pipe_phv_in_data_128,
  input  [7:0]  io_pipe_phv_in_data_129,
  input  [7:0]  io_pipe_phv_in_data_130,
  input  [7:0]  io_pipe_phv_in_data_131,
  input  [7:0]  io_pipe_phv_in_data_132,
  input  [7:0]  io_pipe_phv_in_data_133,
  input  [7:0]  io_pipe_phv_in_data_134,
  input  [7:0]  io_pipe_phv_in_data_135,
  input  [7:0]  io_pipe_phv_in_data_136,
  input  [7:0]  io_pipe_phv_in_data_137,
  input  [7:0]  io_pipe_phv_in_data_138,
  input  [7:0]  io_pipe_phv_in_data_139,
  input  [7:0]  io_pipe_phv_in_data_140,
  input  [7:0]  io_pipe_phv_in_data_141,
  input  [7:0]  io_pipe_phv_in_data_142,
  input  [7:0]  io_pipe_phv_in_data_143,
  input  [7:0]  io_pipe_phv_in_data_144,
  input  [7:0]  io_pipe_phv_in_data_145,
  input  [7:0]  io_pipe_phv_in_data_146,
  input  [7:0]  io_pipe_phv_in_data_147,
  input  [7:0]  io_pipe_phv_in_data_148,
  input  [7:0]  io_pipe_phv_in_data_149,
  input  [7:0]  io_pipe_phv_in_data_150,
  input  [7:0]  io_pipe_phv_in_data_151,
  input  [7:0]  io_pipe_phv_in_data_152,
  input  [7:0]  io_pipe_phv_in_data_153,
  input  [7:0]  io_pipe_phv_in_data_154,
  input  [7:0]  io_pipe_phv_in_data_155,
  input  [7:0]  io_pipe_phv_in_data_156,
  input  [7:0]  io_pipe_phv_in_data_157,
  input  [7:0]  io_pipe_phv_in_data_158,
  input  [7:0]  io_pipe_phv_in_data_159,
  input  [7:0]  io_pipe_phv_in_data_160,
  input  [7:0]  io_pipe_phv_in_data_161,
  input  [7:0]  io_pipe_phv_in_data_162,
  input  [7:0]  io_pipe_phv_in_data_163,
  input  [7:0]  io_pipe_phv_in_data_164,
  input  [7:0]  io_pipe_phv_in_data_165,
  input  [7:0]  io_pipe_phv_in_data_166,
  input  [7:0]  io_pipe_phv_in_data_167,
  input  [7:0]  io_pipe_phv_in_data_168,
  input  [7:0]  io_pipe_phv_in_data_169,
  input  [7:0]  io_pipe_phv_in_data_170,
  input  [7:0]  io_pipe_phv_in_data_171,
  input  [7:0]  io_pipe_phv_in_data_172,
  input  [7:0]  io_pipe_phv_in_data_173,
  input  [7:0]  io_pipe_phv_in_data_174,
  input  [7:0]  io_pipe_phv_in_data_175,
  input  [7:0]  io_pipe_phv_in_data_176,
  input  [7:0]  io_pipe_phv_in_data_177,
  input  [7:0]  io_pipe_phv_in_data_178,
  input  [7:0]  io_pipe_phv_in_data_179,
  input  [7:0]  io_pipe_phv_in_data_180,
  input  [7:0]  io_pipe_phv_in_data_181,
  input  [7:0]  io_pipe_phv_in_data_182,
  input  [7:0]  io_pipe_phv_in_data_183,
  input  [7:0]  io_pipe_phv_in_data_184,
  input  [7:0]  io_pipe_phv_in_data_185,
  input  [7:0]  io_pipe_phv_in_data_186,
  input  [7:0]  io_pipe_phv_in_data_187,
  input  [7:0]  io_pipe_phv_in_data_188,
  input  [7:0]  io_pipe_phv_in_data_189,
  input  [7:0]  io_pipe_phv_in_data_190,
  input  [7:0]  io_pipe_phv_in_data_191,
  input  [7:0]  io_pipe_phv_in_data_192,
  input  [7:0]  io_pipe_phv_in_data_193,
  input  [7:0]  io_pipe_phv_in_data_194,
  input  [7:0]  io_pipe_phv_in_data_195,
  input  [7:0]  io_pipe_phv_in_data_196,
  input  [7:0]  io_pipe_phv_in_data_197,
  input  [7:0]  io_pipe_phv_in_data_198,
  input  [7:0]  io_pipe_phv_in_data_199,
  input  [7:0]  io_pipe_phv_in_data_200,
  input  [7:0]  io_pipe_phv_in_data_201,
  input  [7:0]  io_pipe_phv_in_data_202,
  input  [7:0]  io_pipe_phv_in_data_203,
  input  [7:0]  io_pipe_phv_in_data_204,
  input  [7:0]  io_pipe_phv_in_data_205,
  input  [7:0]  io_pipe_phv_in_data_206,
  input  [7:0]  io_pipe_phv_in_data_207,
  input  [7:0]  io_pipe_phv_in_data_208,
  input  [7:0]  io_pipe_phv_in_data_209,
  input  [7:0]  io_pipe_phv_in_data_210,
  input  [7:0]  io_pipe_phv_in_data_211,
  input  [7:0]  io_pipe_phv_in_data_212,
  input  [7:0]  io_pipe_phv_in_data_213,
  input  [7:0]  io_pipe_phv_in_data_214,
  input  [7:0]  io_pipe_phv_in_data_215,
  input  [7:0]  io_pipe_phv_in_data_216,
  input  [7:0]  io_pipe_phv_in_data_217,
  input  [7:0]  io_pipe_phv_in_data_218,
  input  [7:0]  io_pipe_phv_in_data_219,
  input  [7:0]  io_pipe_phv_in_data_220,
  input  [7:0]  io_pipe_phv_in_data_221,
  input  [7:0]  io_pipe_phv_in_data_222,
  input  [7:0]  io_pipe_phv_in_data_223,
  input  [7:0]  io_pipe_phv_in_data_224,
  input  [7:0]  io_pipe_phv_in_data_225,
  input  [7:0]  io_pipe_phv_in_data_226,
  input  [7:0]  io_pipe_phv_in_data_227,
  input  [7:0]  io_pipe_phv_in_data_228,
  input  [7:0]  io_pipe_phv_in_data_229,
  input  [7:0]  io_pipe_phv_in_data_230,
  input  [7:0]  io_pipe_phv_in_data_231,
  input  [7:0]  io_pipe_phv_in_data_232,
  input  [7:0]  io_pipe_phv_in_data_233,
  input  [7:0]  io_pipe_phv_in_data_234,
  input  [7:0]  io_pipe_phv_in_data_235,
  input  [7:0]  io_pipe_phv_in_data_236,
  input  [7:0]  io_pipe_phv_in_data_237,
  input  [7:0]  io_pipe_phv_in_data_238,
  input  [7:0]  io_pipe_phv_in_data_239,
  input  [7:0]  io_pipe_phv_in_data_240,
  input  [7:0]  io_pipe_phv_in_data_241,
  input  [7:0]  io_pipe_phv_in_data_242,
  input  [7:0]  io_pipe_phv_in_data_243,
  input  [7:0]  io_pipe_phv_in_data_244,
  input  [7:0]  io_pipe_phv_in_data_245,
  input  [7:0]  io_pipe_phv_in_data_246,
  input  [7:0]  io_pipe_phv_in_data_247,
  input  [7:0]  io_pipe_phv_in_data_248,
  input  [7:0]  io_pipe_phv_in_data_249,
  input  [7:0]  io_pipe_phv_in_data_250,
  input  [7:0]  io_pipe_phv_in_data_251,
  input  [7:0]  io_pipe_phv_in_data_252,
  input  [7:0]  io_pipe_phv_in_data_253,
  input  [7:0]  io_pipe_phv_in_data_254,
  input  [7:0]  io_pipe_phv_in_data_255,
  input  [7:0]  io_pipe_phv_in_data_256,
  input  [7:0]  io_pipe_phv_in_data_257,
  input  [7:0]  io_pipe_phv_in_data_258,
  input  [7:0]  io_pipe_phv_in_data_259,
  input  [7:0]  io_pipe_phv_in_data_260,
  input  [7:0]  io_pipe_phv_in_data_261,
  input  [7:0]  io_pipe_phv_in_data_262,
  input  [7:0]  io_pipe_phv_in_data_263,
  input  [7:0]  io_pipe_phv_in_data_264,
  input  [7:0]  io_pipe_phv_in_data_265,
  input  [7:0]  io_pipe_phv_in_data_266,
  input  [7:0]  io_pipe_phv_in_data_267,
  input  [7:0]  io_pipe_phv_in_data_268,
  input  [7:0]  io_pipe_phv_in_data_269,
  input  [7:0]  io_pipe_phv_in_data_270,
  input  [7:0]  io_pipe_phv_in_data_271,
  input  [7:0]  io_pipe_phv_in_data_272,
  input  [7:0]  io_pipe_phv_in_data_273,
  input  [7:0]  io_pipe_phv_in_data_274,
  input  [7:0]  io_pipe_phv_in_data_275,
  input  [7:0]  io_pipe_phv_in_data_276,
  input  [7:0]  io_pipe_phv_in_data_277,
  input  [7:0]  io_pipe_phv_in_data_278,
  input  [7:0]  io_pipe_phv_in_data_279,
  input  [7:0]  io_pipe_phv_in_data_280,
  input  [7:0]  io_pipe_phv_in_data_281,
  input  [7:0]  io_pipe_phv_in_data_282,
  input  [7:0]  io_pipe_phv_in_data_283,
  input  [7:0]  io_pipe_phv_in_data_284,
  input  [7:0]  io_pipe_phv_in_data_285,
  input  [7:0]  io_pipe_phv_in_data_286,
  input  [7:0]  io_pipe_phv_in_data_287,
  input  [7:0]  io_pipe_phv_in_data_288,
  input  [7:0]  io_pipe_phv_in_data_289,
  input  [7:0]  io_pipe_phv_in_data_290,
  input  [7:0]  io_pipe_phv_in_data_291,
  input  [7:0]  io_pipe_phv_in_data_292,
  input  [7:0]  io_pipe_phv_in_data_293,
  input  [7:0]  io_pipe_phv_in_data_294,
  input  [7:0]  io_pipe_phv_in_data_295,
  input  [7:0]  io_pipe_phv_in_data_296,
  input  [7:0]  io_pipe_phv_in_data_297,
  input  [7:0]  io_pipe_phv_in_data_298,
  input  [7:0]  io_pipe_phv_in_data_299,
  input  [7:0]  io_pipe_phv_in_data_300,
  input  [7:0]  io_pipe_phv_in_data_301,
  input  [7:0]  io_pipe_phv_in_data_302,
  input  [7:0]  io_pipe_phv_in_data_303,
  input  [7:0]  io_pipe_phv_in_data_304,
  input  [7:0]  io_pipe_phv_in_data_305,
  input  [7:0]  io_pipe_phv_in_data_306,
  input  [7:0]  io_pipe_phv_in_data_307,
  input  [7:0]  io_pipe_phv_in_data_308,
  input  [7:0]  io_pipe_phv_in_data_309,
  input  [7:0]  io_pipe_phv_in_data_310,
  input  [7:0]  io_pipe_phv_in_data_311,
  input  [7:0]  io_pipe_phv_in_data_312,
  input  [7:0]  io_pipe_phv_in_data_313,
  input  [7:0]  io_pipe_phv_in_data_314,
  input  [7:0]  io_pipe_phv_in_data_315,
  input  [7:0]  io_pipe_phv_in_data_316,
  input  [7:0]  io_pipe_phv_in_data_317,
  input  [7:0]  io_pipe_phv_in_data_318,
  input  [7:0]  io_pipe_phv_in_data_319,
  input  [7:0]  io_pipe_phv_in_data_320,
  input  [7:0]  io_pipe_phv_in_data_321,
  input  [7:0]  io_pipe_phv_in_data_322,
  input  [7:0]  io_pipe_phv_in_data_323,
  input  [7:0]  io_pipe_phv_in_data_324,
  input  [7:0]  io_pipe_phv_in_data_325,
  input  [7:0]  io_pipe_phv_in_data_326,
  input  [7:0]  io_pipe_phv_in_data_327,
  input  [7:0]  io_pipe_phv_in_data_328,
  input  [7:0]  io_pipe_phv_in_data_329,
  input  [7:0]  io_pipe_phv_in_data_330,
  input  [7:0]  io_pipe_phv_in_data_331,
  input  [7:0]  io_pipe_phv_in_data_332,
  input  [7:0]  io_pipe_phv_in_data_333,
  input  [7:0]  io_pipe_phv_in_data_334,
  input  [7:0]  io_pipe_phv_in_data_335,
  input  [7:0]  io_pipe_phv_in_data_336,
  input  [7:0]  io_pipe_phv_in_data_337,
  input  [7:0]  io_pipe_phv_in_data_338,
  input  [7:0]  io_pipe_phv_in_data_339,
  input  [7:0]  io_pipe_phv_in_data_340,
  input  [7:0]  io_pipe_phv_in_data_341,
  input  [7:0]  io_pipe_phv_in_data_342,
  input  [7:0]  io_pipe_phv_in_data_343,
  input  [7:0]  io_pipe_phv_in_data_344,
  input  [7:0]  io_pipe_phv_in_data_345,
  input  [7:0]  io_pipe_phv_in_data_346,
  input  [7:0]  io_pipe_phv_in_data_347,
  input  [7:0]  io_pipe_phv_in_data_348,
  input  [7:0]  io_pipe_phv_in_data_349,
  input  [7:0]  io_pipe_phv_in_data_350,
  input  [7:0]  io_pipe_phv_in_data_351,
  input  [7:0]  io_pipe_phv_in_data_352,
  input  [7:0]  io_pipe_phv_in_data_353,
  input  [7:0]  io_pipe_phv_in_data_354,
  input  [7:0]  io_pipe_phv_in_data_355,
  input  [7:0]  io_pipe_phv_in_data_356,
  input  [7:0]  io_pipe_phv_in_data_357,
  input  [7:0]  io_pipe_phv_in_data_358,
  input  [7:0]  io_pipe_phv_in_data_359,
  input  [7:0]  io_pipe_phv_in_data_360,
  input  [7:0]  io_pipe_phv_in_data_361,
  input  [7:0]  io_pipe_phv_in_data_362,
  input  [7:0]  io_pipe_phv_in_data_363,
  input  [7:0]  io_pipe_phv_in_data_364,
  input  [7:0]  io_pipe_phv_in_data_365,
  input  [7:0]  io_pipe_phv_in_data_366,
  input  [7:0]  io_pipe_phv_in_data_367,
  input  [7:0]  io_pipe_phv_in_data_368,
  input  [7:0]  io_pipe_phv_in_data_369,
  input  [7:0]  io_pipe_phv_in_data_370,
  input  [7:0]  io_pipe_phv_in_data_371,
  input  [7:0]  io_pipe_phv_in_data_372,
  input  [7:0]  io_pipe_phv_in_data_373,
  input  [7:0]  io_pipe_phv_in_data_374,
  input  [7:0]  io_pipe_phv_in_data_375,
  input  [7:0]  io_pipe_phv_in_data_376,
  input  [7:0]  io_pipe_phv_in_data_377,
  input  [7:0]  io_pipe_phv_in_data_378,
  input  [7:0]  io_pipe_phv_in_data_379,
  input  [7:0]  io_pipe_phv_in_data_380,
  input  [7:0]  io_pipe_phv_in_data_381,
  input  [7:0]  io_pipe_phv_in_data_382,
  input  [7:0]  io_pipe_phv_in_data_383,
  output [7:0]  io_pipe_phv_out_data_0,
  output [7:0]  io_pipe_phv_out_data_1,
  output [7:0]  io_pipe_phv_out_data_2,
  output [7:0]  io_pipe_phv_out_data_3,
  output [7:0]  io_pipe_phv_out_data_4,
  output [7:0]  io_pipe_phv_out_data_5,
  output [7:0]  io_pipe_phv_out_data_6,
  output [7:0]  io_pipe_phv_out_data_7,
  output [7:0]  io_pipe_phv_out_data_8,
  output [7:0]  io_pipe_phv_out_data_9,
  output [7:0]  io_pipe_phv_out_data_10,
  output [7:0]  io_pipe_phv_out_data_11,
  output [7:0]  io_pipe_phv_out_data_12,
  output [7:0]  io_pipe_phv_out_data_13,
  output [7:0]  io_pipe_phv_out_data_14,
  output [7:0]  io_pipe_phv_out_data_15,
  output [7:0]  io_pipe_phv_out_data_16,
  output [7:0]  io_pipe_phv_out_data_17,
  output [7:0]  io_pipe_phv_out_data_18,
  output [7:0]  io_pipe_phv_out_data_19,
  output [7:0]  io_pipe_phv_out_data_20,
  output [7:0]  io_pipe_phv_out_data_21,
  output [7:0]  io_pipe_phv_out_data_22,
  output [7:0]  io_pipe_phv_out_data_23,
  output [7:0]  io_pipe_phv_out_data_24,
  output [7:0]  io_pipe_phv_out_data_25,
  output [7:0]  io_pipe_phv_out_data_26,
  output [7:0]  io_pipe_phv_out_data_27,
  output [7:0]  io_pipe_phv_out_data_28,
  output [7:0]  io_pipe_phv_out_data_29,
  output [7:0]  io_pipe_phv_out_data_30,
  output [7:0]  io_pipe_phv_out_data_31,
  output [7:0]  io_pipe_phv_out_data_32,
  output [7:0]  io_pipe_phv_out_data_33,
  output [7:0]  io_pipe_phv_out_data_34,
  output [7:0]  io_pipe_phv_out_data_35,
  output [7:0]  io_pipe_phv_out_data_36,
  output [7:0]  io_pipe_phv_out_data_37,
  output [7:0]  io_pipe_phv_out_data_38,
  output [7:0]  io_pipe_phv_out_data_39,
  output [7:0]  io_pipe_phv_out_data_40,
  output [7:0]  io_pipe_phv_out_data_41,
  output [7:0]  io_pipe_phv_out_data_42,
  output [7:0]  io_pipe_phv_out_data_43,
  output [7:0]  io_pipe_phv_out_data_44,
  output [7:0]  io_pipe_phv_out_data_45,
  output [7:0]  io_pipe_phv_out_data_46,
  output [7:0]  io_pipe_phv_out_data_47,
  output [7:0]  io_pipe_phv_out_data_48,
  output [7:0]  io_pipe_phv_out_data_49,
  output [7:0]  io_pipe_phv_out_data_50,
  output [7:0]  io_pipe_phv_out_data_51,
  output [7:0]  io_pipe_phv_out_data_52,
  output [7:0]  io_pipe_phv_out_data_53,
  output [7:0]  io_pipe_phv_out_data_54,
  output [7:0]  io_pipe_phv_out_data_55,
  output [7:0]  io_pipe_phv_out_data_56,
  output [7:0]  io_pipe_phv_out_data_57,
  output [7:0]  io_pipe_phv_out_data_58,
  output [7:0]  io_pipe_phv_out_data_59,
  output [7:0]  io_pipe_phv_out_data_60,
  output [7:0]  io_pipe_phv_out_data_61,
  output [7:0]  io_pipe_phv_out_data_62,
  output [7:0]  io_pipe_phv_out_data_63,
  output [7:0]  io_pipe_phv_out_data_64,
  output [7:0]  io_pipe_phv_out_data_65,
  output [7:0]  io_pipe_phv_out_data_66,
  output [7:0]  io_pipe_phv_out_data_67,
  output [7:0]  io_pipe_phv_out_data_68,
  output [7:0]  io_pipe_phv_out_data_69,
  output [7:0]  io_pipe_phv_out_data_70,
  output [7:0]  io_pipe_phv_out_data_71,
  output [7:0]  io_pipe_phv_out_data_72,
  output [7:0]  io_pipe_phv_out_data_73,
  output [7:0]  io_pipe_phv_out_data_74,
  output [7:0]  io_pipe_phv_out_data_75,
  output [7:0]  io_pipe_phv_out_data_76,
  output [7:0]  io_pipe_phv_out_data_77,
  output [7:0]  io_pipe_phv_out_data_78,
  output [7:0]  io_pipe_phv_out_data_79,
  output [7:0]  io_pipe_phv_out_data_80,
  output [7:0]  io_pipe_phv_out_data_81,
  output [7:0]  io_pipe_phv_out_data_82,
  output [7:0]  io_pipe_phv_out_data_83,
  output [7:0]  io_pipe_phv_out_data_84,
  output [7:0]  io_pipe_phv_out_data_85,
  output [7:0]  io_pipe_phv_out_data_86,
  output [7:0]  io_pipe_phv_out_data_87,
  output [7:0]  io_pipe_phv_out_data_88,
  output [7:0]  io_pipe_phv_out_data_89,
  output [7:0]  io_pipe_phv_out_data_90,
  output [7:0]  io_pipe_phv_out_data_91,
  output [7:0]  io_pipe_phv_out_data_92,
  output [7:0]  io_pipe_phv_out_data_93,
  output [7:0]  io_pipe_phv_out_data_94,
  output [7:0]  io_pipe_phv_out_data_95,
  output [7:0]  io_pipe_phv_out_data_96,
  output [7:0]  io_pipe_phv_out_data_97,
  output [7:0]  io_pipe_phv_out_data_98,
  output [7:0]  io_pipe_phv_out_data_99,
  output [7:0]  io_pipe_phv_out_data_100,
  output [7:0]  io_pipe_phv_out_data_101,
  output [7:0]  io_pipe_phv_out_data_102,
  output [7:0]  io_pipe_phv_out_data_103,
  output [7:0]  io_pipe_phv_out_data_104,
  output [7:0]  io_pipe_phv_out_data_105,
  output [7:0]  io_pipe_phv_out_data_106,
  output [7:0]  io_pipe_phv_out_data_107,
  output [7:0]  io_pipe_phv_out_data_108,
  output [7:0]  io_pipe_phv_out_data_109,
  output [7:0]  io_pipe_phv_out_data_110,
  output [7:0]  io_pipe_phv_out_data_111,
  output [7:0]  io_pipe_phv_out_data_112,
  output [7:0]  io_pipe_phv_out_data_113,
  output [7:0]  io_pipe_phv_out_data_114,
  output [7:0]  io_pipe_phv_out_data_115,
  output [7:0]  io_pipe_phv_out_data_116,
  output [7:0]  io_pipe_phv_out_data_117,
  output [7:0]  io_pipe_phv_out_data_118,
  output [7:0]  io_pipe_phv_out_data_119,
  output [7:0]  io_pipe_phv_out_data_120,
  output [7:0]  io_pipe_phv_out_data_121,
  output [7:0]  io_pipe_phv_out_data_122,
  output [7:0]  io_pipe_phv_out_data_123,
  output [7:0]  io_pipe_phv_out_data_124,
  output [7:0]  io_pipe_phv_out_data_125,
  output [7:0]  io_pipe_phv_out_data_126,
  output [7:0]  io_pipe_phv_out_data_127,
  output [7:0]  io_pipe_phv_out_data_128,
  output [7:0]  io_pipe_phv_out_data_129,
  output [7:0]  io_pipe_phv_out_data_130,
  output [7:0]  io_pipe_phv_out_data_131,
  output [7:0]  io_pipe_phv_out_data_132,
  output [7:0]  io_pipe_phv_out_data_133,
  output [7:0]  io_pipe_phv_out_data_134,
  output [7:0]  io_pipe_phv_out_data_135,
  output [7:0]  io_pipe_phv_out_data_136,
  output [7:0]  io_pipe_phv_out_data_137,
  output [7:0]  io_pipe_phv_out_data_138,
  output [7:0]  io_pipe_phv_out_data_139,
  output [7:0]  io_pipe_phv_out_data_140,
  output [7:0]  io_pipe_phv_out_data_141,
  output [7:0]  io_pipe_phv_out_data_142,
  output [7:0]  io_pipe_phv_out_data_143,
  output [7:0]  io_pipe_phv_out_data_144,
  output [7:0]  io_pipe_phv_out_data_145,
  output [7:0]  io_pipe_phv_out_data_146,
  output [7:0]  io_pipe_phv_out_data_147,
  output [7:0]  io_pipe_phv_out_data_148,
  output [7:0]  io_pipe_phv_out_data_149,
  output [7:0]  io_pipe_phv_out_data_150,
  output [7:0]  io_pipe_phv_out_data_151,
  output [7:0]  io_pipe_phv_out_data_152,
  output [7:0]  io_pipe_phv_out_data_153,
  output [7:0]  io_pipe_phv_out_data_154,
  output [7:0]  io_pipe_phv_out_data_155,
  output [7:0]  io_pipe_phv_out_data_156,
  output [7:0]  io_pipe_phv_out_data_157,
  output [7:0]  io_pipe_phv_out_data_158,
  output [7:0]  io_pipe_phv_out_data_159,
  output [7:0]  io_pipe_phv_out_data_160,
  output [7:0]  io_pipe_phv_out_data_161,
  output [7:0]  io_pipe_phv_out_data_162,
  output [7:0]  io_pipe_phv_out_data_163,
  output [7:0]  io_pipe_phv_out_data_164,
  output [7:0]  io_pipe_phv_out_data_165,
  output [7:0]  io_pipe_phv_out_data_166,
  output [7:0]  io_pipe_phv_out_data_167,
  output [7:0]  io_pipe_phv_out_data_168,
  output [7:0]  io_pipe_phv_out_data_169,
  output [7:0]  io_pipe_phv_out_data_170,
  output [7:0]  io_pipe_phv_out_data_171,
  output [7:0]  io_pipe_phv_out_data_172,
  output [7:0]  io_pipe_phv_out_data_173,
  output [7:0]  io_pipe_phv_out_data_174,
  output [7:0]  io_pipe_phv_out_data_175,
  output [7:0]  io_pipe_phv_out_data_176,
  output [7:0]  io_pipe_phv_out_data_177,
  output [7:0]  io_pipe_phv_out_data_178,
  output [7:0]  io_pipe_phv_out_data_179,
  output [7:0]  io_pipe_phv_out_data_180,
  output [7:0]  io_pipe_phv_out_data_181,
  output [7:0]  io_pipe_phv_out_data_182,
  output [7:0]  io_pipe_phv_out_data_183,
  output [7:0]  io_pipe_phv_out_data_184,
  output [7:0]  io_pipe_phv_out_data_185,
  output [7:0]  io_pipe_phv_out_data_186,
  output [7:0]  io_pipe_phv_out_data_187,
  output [7:0]  io_pipe_phv_out_data_188,
  output [7:0]  io_pipe_phv_out_data_189,
  output [7:0]  io_pipe_phv_out_data_190,
  output [7:0]  io_pipe_phv_out_data_191,
  output [7:0]  io_pipe_phv_out_data_192,
  output [7:0]  io_pipe_phv_out_data_193,
  output [7:0]  io_pipe_phv_out_data_194,
  output [7:0]  io_pipe_phv_out_data_195,
  output [7:0]  io_pipe_phv_out_data_196,
  output [7:0]  io_pipe_phv_out_data_197,
  output [7:0]  io_pipe_phv_out_data_198,
  output [7:0]  io_pipe_phv_out_data_199,
  output [7:0]  io_pipe_phv_out_data_200,
  output [7:0]  io_pipe_phv_out_data_201,
  output [7:0]  io_pipe_phv_out_data_202,
  output [7:0]  io_pipe_phv_out_data_203,
  output [7:0]  io_pipe_phv_out_data_204,
  output [7:0]  io_pipe_phv_out_data_205,
  output [7:0]  io_pipe_phv_out_data_206,
  output [7:0]  io_pipe_phv_out_data_207,
  output [7:0]  io_pipe_phv_out_data_208,
  output [7:0]  io_pipe_phv_out_data_209,
  output [7:0]  io_pipe_phv_out_data_210,
  output [7:0]  io_pipe_phv_out_data_211,
  output [7:0]  io_pipe_phv_out_data_212,
  output [7:0]  io_pipe_phv_out_data_213,
  output [7:0]  io_pipe_phv_out_data_214,
  output [7:0]  io_pipe_phv_out_data_215,
  output [7:0]  io_pipe_phv_out_data_216,
  output [7:0]  io_pipe_phv_out_data_217,
  output [7:0]  io_pipe_phv_out_data_218,
  output [7:0]  io_pipe_phv_out_data_219,
  output [7:0]  io_pipe_phv_out_data_220,
  output [7:0]  io_pipe_phv_out_data_221,
  output [7:0]  io_pipe_phv_out_data_222,
  output [7:0]  io_pipe_phv_out_data_223,
  output [7:0]  io_pipe_phv_out_data_224,
  output [7:0]  io_pipe_phv_out_data_225,
  output [7:0]  io_pipe_phv_out_data_226,
  output [7:0]  io_pipe_phv_out_data_227,
  output [7:0]  io_pipe_phv_out_data_228,
  output [7:0]  io_pipe_phv_out_data_229,
  output [7:0]  io_pipe_phv_out_data_230,
  output [7:0]  io_pipe_phv_out_data_231,
  output [7:0]  io_pipe_phv_out_data_232,
  output [7:0]  io_pipe_phv_out_data_233,
  output [7:0]  io_pipe_phv_out_data_234,
  output [7:0]  io_pipe_phv_out_data_235,
  output [7:0]  io_pipe_phv_out_data_236,
  output [7:0]  io_pipe_phv_out_data_237,
  output [7:0]  io_pipe_phv_out_data_238,
  output [7:0]  io_pipe_phv_out_data_239,
  output [7:0]  io_pipe_phv_out_data_240,
  output [7:0]  io_pipe_phv_out_data_241,
  output [7:0]  io_pipe_phv_out_data_242,
  output [7:0]  io_pipe_phv_out_data_243,
  output [7:0]  io_pipe_phv_out_data_244,
  output [7:0]  io_pipe_phv_out_data_245,
  output [7:0]  io_pipe_phv_out_data_246,
  output [7:0]  io_pipe_phv_out_data_247,
  output [7:0]  io_pipe_phv_out_data_248,
  output [7:0]  io_pipe_phv_out_data_249,
  output [7:0]  io_pipe_phv_out_data_250,
  output [7:0]  io_pipe_phv_out_data_251,
  output [7:0]  io_pipe_phv_out_data_252,
  output [7:0]  io_pipe_phv_out_data_253,
  output [7:0]  io_pipe_phv_out_data_254,
  output [7:0]  io_pipe_phv_out_data_255,
  output [7:0]  io_pipe_phv_out_data_256,
  output [7:0]  io_pipe_phv_out_data_257,
  output [7:0]  io_pipe_phv_out_data_258,
  output [7:0]  io_pipe_phv_out_data_259,
  output [7:0]  io_pipe_phv_out_data_260,
  output [7:0]  io_pipe_phv_out_data_261,
  output [7:0]  io_pipe_phv_out_data_262,
  output [7:0]  io_pipe_phv_out_data_263,
  output [7:0]  io_pipe_phv_out_data_264,
  output [7:0]  io_pipe_phv_out_data_265,
  output [7:0]  io_pipe_phv_out_data_266,
  output [7:0]  io_pipe_phv_out_data_267,
  output [7:0]  io_pipe_phv_out_data_268,
  output [7:0]  io_pipe_phv_out_data_269,
  output [7:0]  io_pipe_phv_out_data_270,
  output [7:0]  io_pipe_phv_out_data_271,
  output [7:0]  io_pipe_phv_out_data_272,
  output [7:0]  io_pipe_phv_out_data_273,
  output [7:0]  io_pipe_phv_out_data_274,
  output [7:0]  io_pipe_phv_out_data_275,
  output [7:0]  io_pipe_phv_out_data_276,
  output [7:0]  io_pipe_phv_out_data_277,
  output [7:0]  io_pipe_phv_out_data_278,
  output [7:0]  io_pipe_phv_out_data_279,
  output [7:0]  io_pipe_phv_out_data_280,
  output [7:0]  io_pipe_phv_out_data_281,
  output [7:0]  io_pipe_phv_out_data_282,
  output [7:0]  io_pipe_phv_out_data_283,
  output [7:0]  io_pipe_phv_out_data_284,
  output [7:0]  io_pipe_phv_out_data_285,
  output [7:0]  io_pipe_phv_out_data_286,
  output [7:0]  io_pipe_phv_out_data_287,
  output [7:0]  io_pipe_phv_out_data_288,
  output [7:0]  io_pipe_phv_out_data_289,
  output [7:0]  io_pipe_phv_out_data_290,
  output [7:0]  io_pipe_phv_out_data_291,
  output [7:0]  io_pipe_phv_out_data_292,
  output [7:0]  io_pipe_phv_out_data_293,
  output [7:0]  io_pipe_phv_out_data_294,
  output [7:0]  io_pipe_phv_out_data_295,
  output [7:0]  io_pipe_phv_out_data_296,
  output [7:0]  io_pipe_phv_out_data_297,
  output [7:0]  io_pipe_phv_out_data_298,
  output [7:0]  io_pipe_phv_out_data_299,
  output [7:0]  io_pipe_phv_out_data_300,
  output [7:0]  io_pipe_phv_out_data_301,
  output [7:0]  io_pipe_phv_out_data_302,
  output [7:0]  io_pipe_phv_out_data_303,
  output [7:0]  io_pipe_phv_out_data_304,
  output [7:0]  io_pipe_phv_out_data_305,
  output [7:0]  io_pipe_phv_out_data_306,
  output [7:0]  io_pipe_phv_out_data_307,
  output [7:0]  io_pipe_phv_out_data_308,
  output [7:0]  io_pipe_phv_out_data_309,
  output [7:0]  io_pipe_phv_out_data_310,
  output [7:0]  io_pipe_phv_out_data_311,
  output [7:0]  io_pipe_phv_out_data_312,
  output [7:0]  io_pipe_phv_out_data_313,
  output [7:0]  io_pipe_phv_out_data_314,
  output [7:0]  io_pipe_phv_out_data_315,
  output [7:0]  io_pipe_phv_out_data_316,
  output [7:0]  io_pipe_phv_out_data_317,
  output [7:0]  io_pipe_phv_out_data_318,
  output [7:0]  io_pipe_phv_out_data_319,
  output [7:0]  io_pipe_phv_out_data_320,
  output [7:0]  io_pipe_phv_out_data_321,
  output [7:0]  io_pipe_phv_out_data_322,
  output [7:0]  io_pipe_phv_out_data_323,
  output [7:0]  io_pipe_phv_out_data_324,
  output [7:0]  io_pipe_phv_out_data_325,
  output [7:0]  io_pipe_phv_out_data_326,
  output [7:0]  io_pipe_phv_out_data_327,
  output [7:0]  io_pipe_phv_out_data_328,
  output [7:0]  io_pipe_phv_out_data_329,
  output [7:0]  io_pipe_phv_out_data_330,
  output [7:0]  io_pipe_phv_out_data_331,
  output [7:0]  io_pipe_phv_out_data_332,
  output [7:0]  io_pipe_phv_out_data_333,
  output [7:0]  io_pipe_phv_out_data_334,
  output [7:0]  io_pipe_phv_out_data_335,
  output [7:0]  io_pipe_phv_out_data_336,
  output [7:0]  io_pipe_phv_out_data_337,
  output [7:0]  io_pipe_phv_out_data_338,
  output [7:0]  io_pipe_phv_out_data_339,
  output [7:0]  io_pipe_phv_out_data_340,
  output [7:0]  io_pipe_phv_out_data_341,
  output [7:0]  io_pipe_phv_out_data_342,
  output [7:0]  io_pipe_phv_out_data_343,
  output [7:0]  io_pipe_phv_out_data_344,
  output [7:0]  io_pipe_phv_out_data_345,
  output [7:0]  io_pipe_phv_out_data_346,
  output [7:0]  io_pipe_phv_out_data_347,
  output [7:0]  io_pipe_phv_out_data_348,
  output [7:0]  io_pipe_phv_out_data_349,
  output [7:0]  io_pipe_phv_out_data_350,
  output [7:0]  io_pipe_phv_out_data_351,
  output [7:0]  io_pipe_phv_out_data_352,
  output [7:0]  io_pipe_phv_out_data_353,
  output [7:0]  io_pipe_phv_out_data_354,
  output [7:0]  io_pipe_phv_out_data_355,
  output [7:0]  io_pipe_phv_out_data_356,
  output [7:0]  io_pipe_phv_out_data_357,
  output [7:0]  io_pipe_phv_out_data_358,
  output [7:0]  io_pipe_phv_out_data_359,
  output [7:0]  io_pipe_phv_out_data_360,
  output [7:0]  io_pipe_phv_out_data_361,
  output [7:0]  io_pipe_phv_out_data_362,
  output [7:0]  io_pipe_phv_out_data_363,
  output [7:0]  io_pipe_phv_out_data_364,
  output [7:0]  io_pipe_phv_out_data_365,
  output [7:0]  io_pipe_phv_out_data_366,
  output [7:0]  io_pipe_phv_out_data_367,
  output [7:0]  io_pipe_phv_out_data_368,
  output [7:0]  io_pipe_phv_out_data_369,
  output [7:0]  io_pipe_phv_out_data_370,
  output [7:0]  io_pipe_phv_out_data_371,
  output [7:0]  io_pipe_phv_out_data_372,
  output [7:0]  io_pipe_phv_out_data_373,
  output [7:0]  io_pipe_phv_out_data_374,
  output [7:0]  io_pipe_phv_out_data_375,
  output [7:0]  io_pipe_phv_out_data_376,
  output [7:0]  io_pipe_phv_out_data_377,
  output [7:0]  io_pipe_phv_out_data_378,
  output [7:0]  io_pipe_phv_out_data_379,
  output [7:0]  io_pipe_phv_out_data_380,
  output [7:0]  io_pipe_phv_out_data_381,
  output [7:0]  io_pipe_phv_out_data_382,
  output [7:0]  io_pipe_phv_out_data_383,
  output [7:0]  io_pipe_phv_out_data_384,
  output [7:0]  io_pipe_phv_out_data_385,
  output [7:0]  io_pipe_phv_out_data_386,
  output [7:0]  io_pipe_phv_out_data_387,
  output [7:0]  io_pipe_phv_out_data_388,
  output [7:0]  io_pipe_phv_out_data_389,
  output [7:0]  io_pipe_phv_out_data_390,
  output [7:0]  io_pipe_phv_out_data_391,
  output [7:0]  io_pipe_phv_out_data_392,
  output [7:0]  io_pipe_phv_out_data_393,
  output [7:0]  io_pipe_phv_out_data_394,
  output [7:0]  io_pipe_phv_out_data_395,
  output [7:0]  io_pipe_phv_out_data_396,
  output [7:0]  io_pipe_phv_out_data_397,
  output [7:0]  io_pipe_phv_out_data_398,
  output [7:0]  io_pipe_phv_out_data_399,
  output [7:0]  io_pipe_phv_out_data_400,
  output [7:0]  io_pipe_phv_out_data_401,
  output [7:0]  io_pipe_phv_out_data_402,
  output [7:0]  io_pipe_phv_out_data_403,
  output [7:0]  io_pipe_phv_out_data_404,
  output [7:0]  io_pipe_phv_out_data_405,
  output [7:0]  io_pipe_phv_out_data_406,
  output [7:0]  io_pipe_phv_out_data_407,
  output [7:0]  io_pipe_phv_out_data_408,
  output [7:0]  io_pipe_phv_out_data_409,
  output [7:0]  io_pipe_phv_out_data_410,
  output [7:0]  io_pipe_phv_out_data_411,
  output [7:0]  io_pipe_phv_out_data_412,
  output [7:0]  io_pipe_phv_out_data_413,
  output [7:0]  io_pipe_phv_out_data_414,
  output [7:0]  io_pipe_phv_out_data_415,
  output [7:0]  io_pipe_phv_out_data_416,
  output [7:0]  io_pipe_phv_out_data_417,
  output [7:0]  io_pipe_phv_out_data_418,
  output [7:0]  io_pipe_phv_out_data_419,
  output [7:0]  io_pipe_phv_out_data_420,
  output [7:0]  io_pipe_phv_out_data_421,
  output [7:0]  io_pipe_phv_out_data_422,
  output [7:0]  io_pipe_phv_out_data_423,
  output [7:0]  io_pipe_phv_out_data_424,
  output [7:0]  io_pipe_phv_out_data_425,
  output [7:0]  io_pipe_phv_out_data_426,
  output [7:0]  io_pipe_phv_out_data_427,
  output [7:0]  io_pipe_phv_out_data_428,
  output [7:0]  io_pipe_phv_out_data_429,
  output [7:0]  io_pipe_phv_out_data_430,
  output [7:0]  io_pipe_phv_out_data_431,
  output [7:0]  io_pipe_phv_out_data_432,
  output [7:0]  io_pipe_phv_out_data_433,
  output [7:0]  io_pipe_phv_out_data_434,
  output [7:0]  io_pipe_phv_out_data_435,
  output [7:0]  io_pipe_phv_out_data_436,
  output [7:0]  io_pipe_phv_out_data_437,
  output [7:0]  io_pipe_phv_out_data_438,
  output [7:0]  io_pipe_phv_out_data_439,
  output [7:0]  io_pipe_phv_out_data_440,
  output [7:0]  io_pipe_phv_out_data_441,
  output [7:0]  io_pipe_phv_out_data_442,
  output [7:0]  io_pipe_phv_out_data_443,
  output [7:0]  io_pipe_phv_out_data_444,
  output [7:0]  io_pipe_phv_out_data_445,
  output [7:0]  io_pipe_phv_out_data_446,
  output [7:0]  io_pipe_phv_out_data_447,
  output [7:0]  io_pipe_phv_out_data_448,
  output [7:0]  io_pipe_phv_out_data_449,
  output [7:0]  io_pipe_phv_out_data_450,
  output [7:0]  io_pipe_phv_out_data_451,
  output [7:0]  io_pipe_phv_out_data_452,
  output [7:0]  io_pipe_phv_out_data_453,
  output [7:0]  io_pipe_phv_out_data_454,
  output [7:0]  io_pipe_phv_out_data_455,
  output [7:0]  io_pipe_phv_out_data_456,
  output [7:0]  io_pipe_phv_out_data_457,
  output [7:0]  io_pipe_phv_out_data_458,
  output [7:0]  io_pipe_phv_out_data_459,
  output [7:0]  io_pipe_phv_out_data_460,
  output [7:0]  io_pipe_phv_out_data_461,
  output [7:0]  io_pipe_phv_out_data_462,
  output [7:0]  io_pipe_phv_out_data_463,
  output [7:0]  io_pipe_phv_out_data_464,
  output [7:0]  io_pipe_phv_out_data_465,
  output [7:0]  io_pipe_phv_out_data_466,
  output [7:0]  io_pipe_phv_out_data_467,
  output [7:0]  io_pipe_phv_out_data_468,
  output [7:0]  io_pipe_phv_out_data_469,
  output [7:0]  io_pipe_phv_out_data_470,
  output [7:0]  io_pipe_phv_out_data_471,
  output [7:0]  io_pipe_phv_out_data_472,
  output [7:0]  io_pipe_phv_out_data_473,
  output [7:0]  io_pipe_phv_out_data_474,
  output [7:0]  io_pipe_phv_out_data_475,
  output [7:0]  io_pipe_phv_out_data_476,
  output [7:0]  io_pipe_phv_out_data_477,
  output [7:0]  io_pipe_phv_out_data_478,
  output [7:0]  io_pipe_phv_out_data_479,
  output [7:0]  io_pipe_phv_out_data_480,
  output [7:0]  io_pipe_phv_out_data_481,
  output [7:0]  io_pipe_phv_out_data_482,
  output [7:0]  io_pipe_phv_out_data_483,
  output [7:0]  io_pipe_phv_out_data_484,
  output [7:0]  io_pipe_phv_out_data_485,
  output [7:0]  io_pipe_phv_out_data_486,
  output [7:0]  io_pipe_phv_out_data_487,
  output [7:0]  io_pipe_phv_out_data_488,
  output [7:0]  io_pipe_phv_out_data_489,
  output [7:0]  io_pipe_phv_out_data_490,
  output [7:0]  io_pipe_phv_out_data_491,
  output [7:0]  io_pipe_phv_out_data_492,
  output [7:0]  io_pipe_phv_out_data_493,
  output [7:0]  io_pipe_phv_out_data_494,
  output [7:0]  io_pipe_phv_out_data_495,
  output [7:0]  io_pipe_phv_out_data_496,
  output [7:0]  io_pipe_phv_out_data_497,
  output [7:0]  io_pipe_phv_out_data_498,
  output [7:0]  io_pipe_phv_out_data_499,
  output [7:0]  io_pipe_phv_out_data_500,
  output [7:0]  io_pipe_phv_out_data_501,
  output [7:0]  io_pipe_phv_out_data_502,
  output [7:0]  io_pipe_phv_out_data_503,
  output [7:0]  io_pipe_phv_out_data_504,
  output [7:0]  io_pipe_phv_out_data_505,
  output [7:0]  io_pipe_phv_out_data_506,
  output [7:0]  io_pipe_phv_out_data_507,
  output [7:0]  io_pipe_phv_out_data_508,
  output [7:0]  io_pipe_phv_out_data_509,
  output [7:0]  io_pipe_phv_out_data_510,
  output [7:0]  io_pipe_phv_out_data_511,
  output [3:0]  io_pipe_phv_out_next_processor_id,
  output        io_pipe_phv_out_next_config_id,
  input         io_mod_en,
  input         io_mod_last_mau_id_mod,
  input  [3:0]  io_mod_last_mau_id,
  input  [2:0]  io_mod_cs,
  input         io_mod_module_mod_state_id_mod,
  input  [7:0]  io_mod_module_mod_state_id,
  input         io_mod_module_mod_sram_w_cs,
  input         io_mod_module_mod_sram_w_en,
  input  [7:0]  io_mod_module_mod_sram_w_addr,
  input  [63:0] io_mod_module_mod_sram_w_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  mau_0_clock; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_0; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_1; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_2; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_3; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_4; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_5; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_6; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_7; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_8; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_9; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_10; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_11; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_12; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_13; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_14; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_15; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_16; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_17; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_18; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_19; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_20; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_21; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_22; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_23; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_24; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_25; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_26; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_27; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_28; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_29; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_30; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_31; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_32; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_33; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_34; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_35; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_36; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_37; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_38; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_39; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_40; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_41; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_42; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_43; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_44; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_45; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_46; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_47; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_48; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_49; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_50; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_51; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_52; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_53; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_54; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_55; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_56; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_57; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_58; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_59; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_60; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_61; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_62; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_63; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_64; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_65; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_66; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_67; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_68; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_69; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_70; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_71; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_72; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_73; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_74; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_75; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_76; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_77; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_78; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_79; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_80; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_81; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_82; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_83; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_84; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_85; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_86; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_87; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_88; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_89; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_90; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_91; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_92; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_93; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_94; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_95; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_96; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_97; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_98; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_99; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_100; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_101; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_102; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_103; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_104; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_105; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_106; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_107; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_108; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_109; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_110; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_111; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_112; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_113; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_114; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_115; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_116; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_117; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_118; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_119; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_120; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_121; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_122; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_123; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_124; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_125; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_126; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_127; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_128; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_129; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_130; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_131; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_132; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_133; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_134; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_135; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_136; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_137; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_138; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_139; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_140; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_141; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_142; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_143; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_144; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_145; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_146; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_147; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_148; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_149; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_150; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_151; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_152; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_153; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_154; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_155; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_156; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_157; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_158; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_159; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_160; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_161; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_162; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_163; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_164; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_165; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_166; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_167; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_168; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_169; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_170; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_171; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_172; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_173; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_174; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_175; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_176; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_177; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_178; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_179; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_180; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_181; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_182; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_183; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_184; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_185; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_186; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_187; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_188; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_189; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_190; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_191; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_192; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_193; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_194; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_195; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_196; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_197; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_198; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_199; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_200; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_201; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_202; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_203; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_204; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_205; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_206; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_207; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_208; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_209; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_210; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_211; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_212; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_213; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_214; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_215; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_216; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_217; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_218; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_219; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_220; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_221; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_222; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_223; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_224; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_225; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_226; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_227; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_228; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_229; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_230; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_231; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_232; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_233; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_234; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_235; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_236; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_237; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_238; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_239; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_240; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_241; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_242; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_243; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_244; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_245; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_246; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_247; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_248; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_249; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_250; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_251; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_252; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_253; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_254; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_255; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_256; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_257; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_258; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_259; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_260; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_261; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_262; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_263; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_264; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_265; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_266; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_267; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_268; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_269; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_270; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_271; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_272; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_273; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_274; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_275; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_276; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_277; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_278; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_279; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_280; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_281; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_282; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_283; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_284; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_285; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_286; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_287; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_288; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_289; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_290; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_291; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_292; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_293; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_294; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_295; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_296; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_297; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_298; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_299; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_300; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_301; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_302; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_303; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_304; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_305; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_306; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_307; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_308; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_309; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_310; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_311; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_312; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_313; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_314; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_315; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_316; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_317; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_318; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_319; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_320; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_321; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_322; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_323; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_324; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_325; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_326; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_327; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_328; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_329; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_330; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_331; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_332; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_333; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_334; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_335; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_336; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_337; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_338; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_339; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_340; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_341; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_342; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_343; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_344; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_345; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_346; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_347; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_348; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_349; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_350; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_351; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_352; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_353; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_354; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_355; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_356; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_357; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_358; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_359; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_360; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_361; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_362; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_363; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_364; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_365; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_366; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_367; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_368; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_369; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_370; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_371; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_372; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_373; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_374; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_375; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_376; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_377; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_378; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_379; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_380; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_381; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_382; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_383; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_384; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_385; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_386; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_387; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_388; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_389; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_390; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_391; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_392; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_393; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_394; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_395; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_396; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_397; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_398; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_399; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_400; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_401; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_402; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_403; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_404; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_405; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_406; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_407; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_408; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_409; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_410; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_411; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_412; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_413; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_414; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_415; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_416; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_417; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_418; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_419; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_420; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_421; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_422; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_423; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_424; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_425; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_426; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_427; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_428; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_429; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_430; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_431; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_432; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_433; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_434; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_435; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_436; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_437; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_438; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_439; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_440; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_441; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_442; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_443; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_444; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_445; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_446; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_447; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_448; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_449; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_450; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_451; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_452; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_453; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_454; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_455; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_456; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_457; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_458; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_459; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_460; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_461; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_462; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_463; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_464; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_465; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_466; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_467; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_468; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_469; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_470; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_471; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_472; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_473; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_474; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_475; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_476; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_477; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_478; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_479; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_480; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_481; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_482; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_483; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_484; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_485; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_486; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_487; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_488; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_489; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_490; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_491; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_492; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_493; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_494; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_495; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_496; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_497; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_498; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_499; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_500; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_501; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_502; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_503; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_504; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_505; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_506; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_507; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_508; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_509; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_510; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_511; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_0; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_1; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_2; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_3; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_4; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_5; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_6; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_7; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_8; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_9; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_10; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_11; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_12; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_13; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_14; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_15; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_parse_current_state; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_parse_current_offset; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_in_parse_transition_field; // @[parser_pisa.scala 31:25]
  wire [3:0] mau_0_io_pipe_phv_in_next_processor_id; // @[parser_pisa.scala 31:25]
  wire  mau_0_io_pipe_phv_in_next_config_id; // @[parser_pisa.scala 31:25]
  wire  mau_0_io_pipe_phv_in_is_valid_processor; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_0; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_1; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_2; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_3; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_4; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_5; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_6; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_7; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_8; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_9; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_10; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_11; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_12; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_13; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_14; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_15; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_16; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_17; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_18; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_19; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_20; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_21; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_22; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_23; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_24; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_25; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_26; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_27; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_28; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_29; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_30; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_31; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_32; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_33; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_34; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_35; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_36; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_37; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_38; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_39; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_40; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_41; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_42; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_43; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_44; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_45; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_46; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_47; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_48; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_49; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_50; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_51; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_52; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_53; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_54; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_55; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_56; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_57; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_58; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_59; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_60; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_61; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_62; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_63; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_64; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_65; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_66; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_67; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_68; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_69; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_70; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_71; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_72; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_73; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_74; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_75; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_76; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_77; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_78; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_79; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_80; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_81; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_82; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_83; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_84; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_85; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_86; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_87; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_88; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_89; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_90; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_91; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_92; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_93; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_94; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_95; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_96; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_97; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_98; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_99; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_100; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_101; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_102; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_103; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_104; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_105; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_106; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_107; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_108; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_109; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_110; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_111; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_112; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_113; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_114; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_115; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_116; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_117; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_118; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_119; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_120; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_121; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_122; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_123; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_124; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_125; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_126; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_127; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_128; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_129; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_130; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_131; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_132; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_133; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_134; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_135; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_136; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_137; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_138; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_139; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_140; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_141; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_142; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_143; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_144; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_145; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_146; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_147; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_148; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_149; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_150; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_151; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_152; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_153; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_154; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_155; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_156; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_157; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_158; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_159; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_160; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_161; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_162; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_163; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_164; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_165; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_166; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_167; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_168; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_169; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_170; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_171; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_172; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_173; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_174; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_175; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_176; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_177; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_178; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_179; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_180; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_181; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_182; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_183; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_184; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_185; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_186; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_187; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_188; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_189; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_190; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_191; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_192; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_193; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_194; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_195; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_196; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_197; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_198; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_199; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_200; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_201; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_202; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_203; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_204; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_205; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_206; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_207; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_208; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_209; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_210; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_211; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_212; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_213; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_214; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_215; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_216; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_217; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_218; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_219; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_220; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_221; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_222; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_223; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_224; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_225; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_226; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_227; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_228; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_229; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_230; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_231; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_232; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_233; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_234; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_235; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_236; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_237; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_238; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_239; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_240; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_241; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_242; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_243; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_244; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_245; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_246; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_247; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_248; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_249; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_250; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_251; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_252; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_253; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_254; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_255; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_256; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_257; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_258; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_259; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_260; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_261; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_262; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_263; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_264; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_265; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_266; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_267; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_268; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_269; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_270; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_271; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_272; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_273; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_274; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_275; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_276; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_277; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_278; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_279; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_280; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_281; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_282; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_283; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_284; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_285; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_286; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_287; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_288; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_289; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_290; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_291; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_292; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_293; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_294; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_295; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_296; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_297; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_298; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_299; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_300; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_301; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_302; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_303; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_304; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_305; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_306; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_307; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_308; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_309; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_310; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_311; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_312; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_313; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_314; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_315; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_316; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_317; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_318; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_319; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_320; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_321; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_322; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_323; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_324; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_325; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_326; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_327; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_328; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_329; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_330; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_331; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_332; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_333; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_334; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_335; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_336; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_337; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_338; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_339; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_340; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_341; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_342; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_343; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_344; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_345; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_346; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_347; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_348; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_349; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_350; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_351; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_352; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_353; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_354; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_355; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_356; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_357; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_358; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_359; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_360; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_361; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_362; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_363; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_364; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_365; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_366; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_367; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_368; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_369; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_370; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_371; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_372; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_373; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_374; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_375; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_376; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_377; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_378; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_379; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_380; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_381; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_382; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_383; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_384; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_385; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_386; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_387; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_388; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_389; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_390; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_391; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_392; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_393; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_394; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_395; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_396; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_397; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_398; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_399; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_400; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_401; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_402; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_403; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_404; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_405; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_406; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_407; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_408; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_409; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_410; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_411; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_412; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_413; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_414; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_415; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_416; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_417; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_418; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_419; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_420; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_421; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_422; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_423; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_424; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_425; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_426; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_427; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_428; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_429; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_430; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_431; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_432; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_433; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_434; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_435; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_436; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_437; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_438; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_439; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_440; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_441; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_442; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_443; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_444; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_445; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_446; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_447; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_448; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_449; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_450; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_451; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_452; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_453; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_454; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_455; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_456; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_457; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_458; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_459; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_460; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_461; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_462; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_463; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_464; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_465; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_466; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_467; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_468; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_469; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_470; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_471; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_472; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_473; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_474; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_475; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_476; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_477; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_478; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_479; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_480; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_481; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_482; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_483; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_484; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_485; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_486; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_487; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_488; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_489; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_490; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_491; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_492; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_493; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_494; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_495; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_496; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_497; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_498; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_499; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_500; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_501; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_502; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_503; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_504; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_505; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_506; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_507; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_508; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_509; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_510; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_511; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_0; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_1; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_2; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_3; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_4; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_5; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_6; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_7; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_8; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_9; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_10; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_11; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_12; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_13; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_14; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_15; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_parse_current_state; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_parse_current_offset; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_out_parse_transition_field; // @[parser_pisa.scala 31:25]
  wire [3:0] mau_0_io_pipe_phv_out_next_processor_id; // @[parser_pisa.scala 31:25]
  wire  mau_0_io_pipe_phv_out_next_config_id; // @[parser_pisa.scala 31:25]
  wire  mau_0_io_pipe_phv_out_is_valid_processor; // @[parser_pisa.scala 31:25]
  wire  mau_0_io_mod_state_id_mod; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_mod_state_id; // @[parser_pisa.scala 31:25]
  wire  mau_0_io_mod_sram_w_cs; // @[parser_pisa.scala 31:25]
  wire  mau_0_io_mod_sram_w_en; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_mod_sram_w_addr; // @[parser_pisa.scala 31:25]
  wire [63:0] mau_0_io_mod_sram_w_data; // @[parser_pisa.scala 31:25]
  wire  mau_1_clock; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_0; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_1; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_2; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_3; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_4; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_5; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_6; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_7; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_8; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_9; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_10; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_11; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_12; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_13; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_14; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_15; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_16; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_17; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_18; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_19; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_20; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_21; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_22; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_23; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_24; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_25; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_26; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_27; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_28; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_29; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_30; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_31; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_32; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_33; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_34; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_35; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_36; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_37; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_38; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_39; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_40; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_41; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_42; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_43; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_44; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_45; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_46; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_47; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_48; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_49; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_50; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_51; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_52; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_53; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_54; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_55; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_56; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_57; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_58; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_59; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_60; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_61; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_62; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_63; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_64; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_65; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_66; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_67; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_68; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_69; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_70; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_71; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_72; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_73; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_74; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_75; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_76; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_77; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_78; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_79; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_80; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_81; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_82; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_83; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_84; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_85; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_86; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_87; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_88; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_89; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_90; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_91; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_92; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_93; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_94; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_95; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_96; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_97; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_98; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_99; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_100; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_101; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_102; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_103; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_104; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_105; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_106; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_107; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_108; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_109; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_110; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_111; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_112; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_113; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_114; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_115; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_116; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_117; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_118; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_119; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_120; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_121; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_122; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_123; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_124; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_125; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_126; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_127; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_128; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_129; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_130; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_131; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_132; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_133; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_134; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_135; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_136; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_137; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_138; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_139; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_140; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_141; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_142; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_143; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_144; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_145; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_146; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_147; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_148; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_149; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_150; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_151; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_152; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_153; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_154; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_155; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_156; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_157; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_158; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_159; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_160; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_161; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_162; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_163; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_164; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_165; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_166; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_167; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_168; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_169; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_170; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_171; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_172; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_173; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_174; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_175; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_176; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_177; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_178; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_179; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_180; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_181; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_182; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_183; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_184; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_185; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_186; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_187; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_188; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_189; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_190; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_191; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_192; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_193; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_194; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_195; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_196; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_197; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_198; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_199; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_200; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_201; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_202; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_203; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_204; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_205; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_206; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_207; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_208; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_209; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_210; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_211; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_212; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_213; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_214; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_215; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_216; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_217; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_218; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_219; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_220; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_221; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_222; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_223; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_224; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_225; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_226; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_227; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_228; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_229; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_230; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_231; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_232; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_233; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_234; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_235; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_236; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_237; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_238; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_239; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_240; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_241; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_242; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_243; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_244; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_245; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_246; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_247; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_248; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_249; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_250; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_251; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_252; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_253; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_254; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_255; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_256; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_257; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_258; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_259; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_260; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_261; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_262; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_263; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_264; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_265; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_266; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_267; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_268; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_269; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_270; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_271; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_272; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_273; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_274; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_275; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_276; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_277; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_278; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_279; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_280; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_281; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_282; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_283; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_284; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_285; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_286; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_287; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_288; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_289; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_290; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_291; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_292; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_293; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_294; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_295; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_296; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_297; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_298; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_299; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_300; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_301; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_302; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_303; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_304; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_305; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_306; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_307; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_308; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_309; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_310; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_311; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_312; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_313; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_314; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_315; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_316; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_317; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_318; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_319; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_320; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_321; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_322; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_323; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_324; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_325; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_326; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_327; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_328; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_329; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_330; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_331; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_332; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_333; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_334; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_335; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_336; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_337; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_338; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_339; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_340; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_341; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_342; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_343; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_344; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_345; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_346; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_347; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_348; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_349; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_350; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_351; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_352; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_353; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_354; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_355; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_356; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_357; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_358; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_359; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_360; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_361; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_362; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_363; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_364; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_365; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_366; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_367; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_368; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_369; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_370; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_371; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_372; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_373; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_374; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_375; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_376; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_377; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_378; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_379; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_380; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_381; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_382; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_383; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_384; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_385; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_386; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_387; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_388; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_389; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_390; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_391; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_392; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_393; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_394; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_395; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_396; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_397; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_398; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_399; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_400; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_401; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_402; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_403; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_404; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_405; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_406; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_407; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_408; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_409; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_410; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_411; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_412; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_413; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_414; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_415; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_416; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_417; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_418; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_419; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_420; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_421; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_422; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_423; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_424; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_425; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_426; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_427; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_428; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_429; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_430; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_431; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_432; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_433; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_434; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_435; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_436; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_437; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_438; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_439; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_440; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_441; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_442; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_443; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_444; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_445; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_446; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_447; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_448; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_449; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_450; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_451; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_452; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_453; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_454; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_455; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_456; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_457; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_458; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_459; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_460; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_461; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_462; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_463; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_464; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_465; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_466; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_467; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_468; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_469; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_470; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_471; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_472; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_473; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_474; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_475; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_476; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_477; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_478; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_479; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_480; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_481; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_482; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_483; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_484; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_485; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_486; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_487; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_488; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_489; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_490; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_491; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_492; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_493; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_494; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_495; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_496; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_497; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_498; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_499; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_500; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_501; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_502; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_503; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_504; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_505; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_506; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_507; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_508; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_509; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_510; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_511; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_0; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_1; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_2; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_3; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_4; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_5; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_6; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_7; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_8; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_9; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_10; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_11; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_12; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_13; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_14; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_15; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_parse_current_state; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_parse_current_offset; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_in_parse_transition_field; // @[parser_pisa.scala 31:25]
  wire [3:0] mau_1_io_pipe_phv_in_next_processor_id; // @[parser_pisa.scala 31:25]
  wire  mau_1_io_pipe_phv_in_next_config_id; // @[parser_pisa.scala 31:25]
  wire  mau_1_io_pipe_phv_in_is_valid_processor; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_0; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_1; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_2; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_3; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_4; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_5; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_6; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_7; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_8; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_9; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_10; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_11; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_12; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_13; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_14; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_15; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_16; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_17; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_18; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_19; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_20; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_21; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_22; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_23; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_24; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_25; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_26; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_27; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_28; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_29; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_30; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_31; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_32; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_33; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_34; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_35; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_36; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_37; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_38; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_39; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_40; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_41; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_42; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_43; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_44; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_45; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_46; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_47; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_48; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_49; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_50; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_51; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_52; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_53; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_54; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_55; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_56; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_57; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_58; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_59; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_60; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_61; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_62; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_63; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_64; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_65; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_66; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_67; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_68; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_69; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_70; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_71; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_72; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_73; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_74; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_75; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_76; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_77; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_78; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_79; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_80; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_81; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_82; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_83; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_84; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_85; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_86; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_87; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_88; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_89; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_90; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_91; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_92; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_93; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_94; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_95; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_96; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_97; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_98; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_99; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_100; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_101; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_102; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_103; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_104; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_105; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_106; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_107; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_108; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_109; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_110; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_111; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_112; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_113; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_114; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_115; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_116; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_117; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_118; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_119; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_120; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_121; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_122; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_123; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_124; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_125; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_126; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_127; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_128; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_129; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_130; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_131; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_132; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_133; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_134; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_135; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_136; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_137; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_138; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_139; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_140; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_141; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_142; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_143; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_144; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_145; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_146; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_147; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_148; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_149; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_150; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_151; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_152; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_153; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_154; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_155; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_156; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_157; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_158; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_159; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_160; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_161; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_162; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_163; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_164; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_165; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_166; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_167; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_168; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_169; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_170; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_171; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_172; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_173; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_174; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_175; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_176; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_177; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_178; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_179; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_180; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_181; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_182; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_183; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_184; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_185; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_186; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_187; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_188; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_189; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_190; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_191; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_192; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_193; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_194; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_195; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_196; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_197; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_198; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_199; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_200; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_201; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_202; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_203; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_204; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_205; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_206; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_207; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_208; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_209; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_210; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_211; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_212; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_213; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_214; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_215; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_216; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_217; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_218; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_219; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_220; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_221; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_222; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_223; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_224; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_225; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_226; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_227; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_228; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_229; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_230; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_231; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_232; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_233; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_234; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_235; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_236; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_237; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_238; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_239; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_240; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_241; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_242; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_243; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_244; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_245; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_246; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_247; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_248; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_249; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_250; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_251; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_252; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_253; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_254; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_255; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_256; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_257; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_258; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_259; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_260; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_261; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_262; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_263; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_264; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_265; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_266; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_267; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_268; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_269; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_270; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_271; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_272; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_273; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_274; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_275; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_276; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_277; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_278; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_279; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_280; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_281; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_282; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_283; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_284; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_285; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_286; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_287; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_288; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_289; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_290; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_291; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_292; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_293; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_294; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_295; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_296; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_297; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_298; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_299; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_300; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_301; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_302; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_303; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_304; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_305; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_306; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_307; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_308; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_309; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_310; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_311; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_312; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_313; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_314; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_315; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_316; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_317; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_318; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_319; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_320; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_321; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_322; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_323; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_324; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_325; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_326; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_327; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_328; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_329; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_330; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_331; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_332; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_333; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_334; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_335; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_336; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_337; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_338; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_339; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_340; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_341; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_342; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_343; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_344; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_345; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_346; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_347; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_348; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_349; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_350; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_351; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_352; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_353; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_354; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_355; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_356; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_357; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_358; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_359; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_360; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_361; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_362; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_363; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_364; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_365; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_366; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_367; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_368; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_369; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_370; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_371; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_372; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_373; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_374; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_375; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_376; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_377; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_378; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_379; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_380; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_381; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_382; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_383; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_384; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_385; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_386; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_387; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_388; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_389; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_390; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_391; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_392; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_393; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_394; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_395; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_396; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_397; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_398; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_399; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_400; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_401; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_402; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_403; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_404; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_405; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_406; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_407; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_408; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_409; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_410; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_411; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_412; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_413; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_414; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_415; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_416; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_417; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_418; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_419; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_420; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_421; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_422; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_423; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_424; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_425; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_426; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_427; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_428; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_429; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_430; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_431; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_432; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_433; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_434; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_435; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_436; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_437; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_438; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_439; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_440; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_441; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_442; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_443; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_444; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_445; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_446; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_447; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_448; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_449; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_450; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_451; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_452; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_453; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_454; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_455; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_456; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_457; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_458; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_459; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_460; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_461; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_462; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_463; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_464; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_465; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_466; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_467; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_468; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_469; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_470; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_471; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_472; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_473; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_474; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_475; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_476; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_477; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_478; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_479; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_480; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_481; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_482; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_483; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_484; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_485; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_486; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_487; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_488; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_489; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_490; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_491; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_492; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_493; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_494; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_495; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_496; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_497; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_498; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_499; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_500; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_501; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_502; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_503; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_504; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_505; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_506; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_507; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_508; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_509; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_510; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_511; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_0; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_1; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_2; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_3; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_4; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_5; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_6; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_7; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_8; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_9; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_10; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_11; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_12; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_13; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_14; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_15; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_parse_current_state; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_parse_current_offset; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_out_parse_transition_field; // @[parser_pisa.scala 31:25]
  wire [3:0] mau_1_io_pipe_phv_out_next_processor_id; // @[parser_pisa.scala 31:25]
  wire  mau_1_io_pipe_phv_out_next_config_id; // @[parser_pisa.scala 31:25]
  wire  mau_1_io_pipe_phv_out_is_valid_processor; // @[parser_pisa.scala 31:25]
  wire  mau_1_io_mod_state_id_mod; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_mod_state_id; // @[parser_pisa.scala 31:25]
  wire  mau_1_io_mod_sram_w_cs; // @[parser_pisa.scala 31:25]
  wire  mau_1_io_mod_sram_w_en; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_mod_sram_w_addr; // @[parser_pisa.scala 31:25]
  wire [63:0] mau_1_io_mod_sram_w_data; // @[parser_pisa.scala 31:25]
  wire  mau_2_clock; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_0; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_1; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_2; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_3; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_4; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_5; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_6; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_7; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_8; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_9; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_10; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_11; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_12; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_13; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_14; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_15; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_16; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_17; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_18; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_19; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_20; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_21; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_22; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_23; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_24; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_25; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_26; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_27; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_28; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_29; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_30; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_31; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_32; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_33; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_34; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_35; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_36; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_37; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_38; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_39; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_40; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_41; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_42; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_43; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_44; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_45; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_46; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_47; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_48; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_49; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_50; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_51; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_52; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_53; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_54; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_55; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_56; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_57; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_58; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_59; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_60; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_61; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_62; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_63; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_64; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_65; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_66; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_67; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_68; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_69; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_70; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_71; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_72; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_73; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_74; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_75; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_76; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_77; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_78; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_79; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_80; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_81; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_82; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_83; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_84; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_85; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_86; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_87; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_88; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_89; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_90; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_91; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_92; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_93; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_94; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_95; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_96; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_97; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_98; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_99; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_100; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_101; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_102; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_103; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_104; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_105; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_106; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_107; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_108; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_109; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_110; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_111; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_112; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_113; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_114; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_115; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_116; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_117; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_118; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_119; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_120; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_121; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_122; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_123; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_124; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_125; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_126; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_127; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_128; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_129; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_130; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_131; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_132; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_133; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_134; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_135; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_136; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_137; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_138; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_139; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_140; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_141; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_142; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_143; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_144; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_145; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_146; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_147; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_148; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_149; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_150; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_151; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_152; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_153; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_154; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_155; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_156; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_157; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_158; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_159; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_160; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_161; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_162; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_163; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_164; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_165; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_166; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_167; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_168; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_169; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_170; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_171; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_172; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_173; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_174; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_175; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_176; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_177; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_178; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_179; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_180; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_181; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_182; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_183; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_184; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_185; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_186; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_187; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_188; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_189; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_190; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_191; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_192; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_193; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_194; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_195; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_196; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_197; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_198; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_199; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_200; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_201; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_202; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_203; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_204; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_205; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_206; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_207; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_208; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_209; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_210; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_211; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_212; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_213; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_214; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_215; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_216; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_217; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_218; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_219; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_220; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_221; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_222; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_223; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_224; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_225; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_226; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_227; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_228; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_229; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_230; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_231; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_232; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_233; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_234; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_235; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_236; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_237; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_238; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_239; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_240; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_241; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_242; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_243; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_244; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_245; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_246; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_247; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_248; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_249; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_250; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_251; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_252; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_253; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_254; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_255; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_256; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_257; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_258; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_259; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_260; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_261; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_262; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_263; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_264; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_265; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_266; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_267; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_268; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_269; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_270; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_271; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_272; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_273; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_274; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_275; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_276; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_277; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_278; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_279; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_280; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_281; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_282; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_283; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_284; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_285; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_286; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_287; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_288; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_289; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_290; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_291; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_292; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_293; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_294; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_295; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_296; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_297; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_298; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_299; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_300; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_301; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_302; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_303; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_304; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_305; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_306; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_307; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_308; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_309; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_310; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_311; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_312; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_313; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_314; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_315; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_316; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_317; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_318; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_319; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_320; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_321; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_322; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_323; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_324; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_325; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_326; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_327; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_328; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_329; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_330; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_331; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_332; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_333; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_334; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_335; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_336; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_337; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_338; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_339; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_340; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_341; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_342; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_343; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_344; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_345; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_346; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_347; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_348; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_349; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_350; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_351; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_352; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_353; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_354; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_355; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_356; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_357; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_358; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_359; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_360; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_361; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_362; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_363; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_364; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_365; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_366; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_367; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_368; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_369; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_370; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_371; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_372; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_373; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_374; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_375; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_376; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_377; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_378; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_379; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_380; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_381; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_382; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_383; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_384; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_385; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_386; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_387; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_388; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_389; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_390; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_391; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_392; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_393; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_394; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_395; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_396; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_397; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_398; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_399; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_400; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_401; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_402; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_403; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_404; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_405; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_406; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_407; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_408; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_409; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_410; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_411; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_412; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_413; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_414; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_415; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_416; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_417; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_418; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_419; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_420; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_421; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_422; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_423; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_424; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_425; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_426; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_427; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_428; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_429; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_430; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_431; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_432; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_433; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_434; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_435; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_436; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_437; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_438; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_439; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_440; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_441; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_442; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_443; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_444; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_445; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_446; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_447; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_448; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_449; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_450; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_451; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_452; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_453; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_454; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_455; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_456; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_457; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_458; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_459; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_460; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_461; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_462; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_463; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_464; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_465; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_466; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_467; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_468; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_469; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_470; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_471; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_472; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_473; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_474; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_475; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_476; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_477; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_478; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_479; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_480; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_481; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_482; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_483; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_484; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_485; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_486; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_487; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_488; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_489; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_490; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_491; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_492; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_493; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_494; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_495; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_496; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_497; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_498; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_499; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_500; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_501; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_502; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_503; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_504; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_505; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_506; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_507; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_508; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_509; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_510; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_511; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_0; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_1; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_2; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_3; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_4; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_5; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_6; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_7; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_8; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_9; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_10; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_11; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_12; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_13; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_14; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_15; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_parse_current_state; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_parse_current_offset; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_in_parse_transition_field; // @[parser_pisa.scala 31:25]
  wire [3:0] mau_2_io_pipe_phv_in_next_processor_id; // @[parser_pisa.scala 31:25]
  wire  mau_2_io_pipe_phv_in_next_config_id; // @[parser_pisa.scala 31:25]
  wire  mau_2_io_pipe_phv_in_is_valid_processor; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_0; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_1; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_2; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_3; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_4; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_5; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_6; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_7; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_8; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_9; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_10; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_11; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_12; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_13; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_14; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_15; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_16; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_17; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_18; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_19; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_20; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_21; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_22; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_23; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_24; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_25; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_26; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_27; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_28; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_29; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_30; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_31; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_32; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_33; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_34; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_35; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_36; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_37; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_38; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_39; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_40; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_41; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_42; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_43; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_44; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_45; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_46; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_47; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_48; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_49; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_50; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_51; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_52; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_53; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_54; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_55; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_56; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_57; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_58; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_59; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_60; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_61; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_62; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_63; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_64; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_65; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_66; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_67; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_68; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_69; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_70; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_71; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_72; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_73; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_74; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_75; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_76; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_77; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_78; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_79; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_80; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_81; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_82; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_83; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_84; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_85; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_86; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_87; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_88; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_89; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_90; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_91; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_92; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_93; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_94; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_95; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_96; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_97; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_98; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_99; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_100; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_101; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_102; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_103; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_104; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_105; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_106; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_107; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_108; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_109; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_110; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_111; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_112; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_113; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_114; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_115; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_116; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_117; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_118; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_119; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_120; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_121; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_122; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_123; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_124; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_125; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_126; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_127; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_128; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_129; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_130; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_131; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_132; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_133; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_134; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_135; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_136; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_137; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_138; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_139; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_140; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_141; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_142; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_143; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_144; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_145; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_146; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_147; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_148; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_149; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_150; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_151; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_152; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_153; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_154; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_155; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_156; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_157; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_158; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_159; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_160; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_161; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_162; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_163; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_164; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_165; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_166; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_167; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_168; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_169; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_170; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_171; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_172; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_173; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_174; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_175; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_176; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_177; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_178; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_179; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_180; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_181; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_182; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_183; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_184; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_185; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_186; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_187; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_188; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_189; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_190; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_191; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_192; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_193; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_194; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_195; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_196; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_197; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_198; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_199; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_200; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_201; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_202; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_203; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_204; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_205; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_206; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_207; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_208; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_209; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_210; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_211; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_212; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_213; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_214; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_215; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_216; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_217; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_218; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_219; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_220; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_221; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_222; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_223; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_224; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_225; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_226; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_227; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_228; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_229; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_230; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_231; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_232; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_233; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_234; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_235; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_236; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_237; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_238; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_239; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_240; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_241; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_242; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_243; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_244; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_245; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_246; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_247; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_248; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_249; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_250; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_251; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_252; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_253; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_254; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_255; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_256; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_257; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_258; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_259; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_260; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_261; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_262; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_263; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_264; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_265; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_266; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_267; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_268; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_269; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_270; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_271; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_272; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_273; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_274; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_275; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_276; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_277; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_278; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_279; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_280; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_281; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_282; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_283; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_284; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_285; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_286; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_287; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_288; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_289; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_290; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_291; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_292; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_293; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_294; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_295; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_296; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_297; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_298; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_299; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_300; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_301; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_302; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_303; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_304; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_305; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_306; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_307; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_308; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_309; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_310; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_311; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_312; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_313; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_314; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_315; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_316; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_317; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_318; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_319; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_320; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_321; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_322; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_323; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_324; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_325; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_326; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_327; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_328; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_329; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_330; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_331; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_332; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_333; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_334; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_335; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_336; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_337; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_338; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_339; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_340; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_341; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_342; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_343; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_344; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_345; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_346; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_347; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_348; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_349; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_350; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_351; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_352; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_353; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_354; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_355; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_356; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_357; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_358; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_359; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_360; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_361; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_362; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_363; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_364; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_365; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_366; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_367; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_368; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_369; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_370; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_371; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_372; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_373; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_374; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_375; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_376; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_377; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_378; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_379; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_380; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_381; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_382; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_383; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_384; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_385; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_386; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_387; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_388; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_389; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_390; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_391; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_392; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_393; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_394; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_395; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_396; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_397; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_398; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_399; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_400; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_401; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_402; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_403; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_404; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_405; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_406; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_407; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_408; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_409; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_410; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_411; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_412; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_413; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_414; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_415; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_416; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_417; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_418; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_419; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_420; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_421; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_422; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_423; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_424; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_425; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_426; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_427; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_428; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_429; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_430; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_431; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_432; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_433; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_434; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_435; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_436; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_437; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_438; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_439; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_440; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_441; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_442; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_443; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_444; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_445; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_446; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_447; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_448; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_449; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_450; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_451; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_452; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_453; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_454; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_455; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_456; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_457; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_458; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_459; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_460; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_461; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_462; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_463; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_464; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_465; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_466; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_467; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_468; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_469; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_470; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_471; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_472; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_473; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_474; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_475; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_476; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_477; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_478; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_479; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_480; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_481; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_482; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_483; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_484; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_485; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_486; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_487; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_488; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_489; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_490; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_491; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_492; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_493; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_494; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_495; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_496; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_497; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_498; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_499; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_500; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_501; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_502; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_503; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_504; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_505; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_506; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_507; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_508; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_509; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_510; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_511; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_0; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_1; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_2; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_3; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_4; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_5; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_6; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_7; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_8; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_9; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_10; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_11; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_12; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_13; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_14; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_15; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_parse_current_state; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_parse_current_offset; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_out_parse_transition_field; // @[parser_pisa.scala 31:25]
  wire [3:0] mau_2_io_pipe_phv_out_next_processor_id; // @[parser_pisa.scala 31:25]
  wire  mau_2_io_pipe_phv_out_next_config_id; // @[parser_pisa.scala 31:25]
  wire  mau_2_io_pipe_phv_out_is_valid_processor; // @[parser_pisa.scala 31:25]
  wire  mau_2_io_mod_state_id_mod; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_mod_state_id; // @[parser_pisa.scala 31:25]
  wire  mau_2_io_mod_sram_w_cs; // @[parser_pisa.scala 31:25]
  wire  mau_2_io_mod_sram_w_en; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_mod_sram_w_addr; // @[parser_pisa.scala 31:25]
  wire [63:0] mau_2_io_mod_sram_w_data; // @[parser_pisa.scala 31:25]
  wire  mau_3_clock; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_0; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_1; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_2; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_3; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_4; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_5; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_6; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_7; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_8; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_9; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_10; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_11; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_12; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_13; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_14; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_15; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_16; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_17; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_18; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_19; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_20; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_21; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_22; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_23; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_24; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_25; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_26; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_27; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_28; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_29; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_30; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_31; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_32; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_33; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_34; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_35; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_36; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_37; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_38; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_39; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_40; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_41; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_42; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_43; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_44; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_45; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_46; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_47; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_48; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_49; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_50; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_51; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_52; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_53; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_54; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_55; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_56; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_57; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_58; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_59; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_60; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_61; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_62; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_63; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_64; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_65; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_66; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_67; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_68; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_69; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_70; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_71; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_72; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_73; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_74; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_75; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_76; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_77; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_78; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_79; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_80; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_81; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_82; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_83; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_84; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_85; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_86; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_87; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_88; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_89; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_90; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_91; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_92; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_93; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_94; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_95; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_96; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_97; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_98; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_99; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_100; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_101; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_102; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_103; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_104; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_105; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_106; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_107; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_108; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_109; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_110; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_111; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_112; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_113; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_114; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_115; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_116; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_117; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_118; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_119; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_120; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_121; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_122; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_123; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_124; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_125; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_126; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_127; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_128; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_129; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_130; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_131; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_132; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_133; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_134; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_135; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_136; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_137; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_138; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_139; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_140; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_141; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_142; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_143; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_144; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_145; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_146; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_147; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_148; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_149; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_150; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_151; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_152; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_153; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_154; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_155; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_156; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_157; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_158; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_159; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_160; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_161; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_162; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_163; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_164; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_165; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_166; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_167; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_168; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_169; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_170; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_171; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_172; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_173; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_174; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_175; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_176; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_177; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_178; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_179; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_180; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_181; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_182; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_183; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_184; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_185; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_186; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_187; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_188; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_189; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_190; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_191; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_192; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_193; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_194; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_195; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_196; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_197; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_198; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_199; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_200; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_201; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_202; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_203; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_204; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_205; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_206; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_207; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_208; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_209; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_210; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_211; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_212; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_213; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_214; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_215; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_216; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_217; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_218; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_219; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_220; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_221; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_222; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_223; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_224; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_225; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_226; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_227; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_228; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_229; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_230; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_231; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_232; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_233; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_234; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_235; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_236; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_237; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_238; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_239; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_240; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_241; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_242; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_243; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_244; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_245; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_246; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_247; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_248; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_249; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_250; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_251; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_252; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_253; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_254; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_255; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_256; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_257; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_258; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_259; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_260; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_261; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_262; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_263; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_264; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_265; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_266; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_267; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_268; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_269; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_270; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_271; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_272; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_273; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_274; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_275; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_276; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_277; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_278; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_279; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_280; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_281; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_282; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_283; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_284; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_285; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_286; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_287; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_288; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_289; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_290; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_291; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_292; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_293; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_294; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_295; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_296; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_297; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_298; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_299; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_300; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_301; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_302; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_303; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_304; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_305; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_306; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_307; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_308; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_309; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_310; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_311; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_312; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_313; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_314; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_315; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_316; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_317; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_318; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_319; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_320; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_321; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_322; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_323; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_324; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_325; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_326; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_327; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_328; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_329; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_330; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_331; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_332; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_333; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_334; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_335; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_336; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_337; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_338; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_339; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_340; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_341; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_342; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_343; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_344; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_345; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_346; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_347; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_348; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_349; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_350; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_351; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_352; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_353; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_354; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_355; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_356; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_357; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_358; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_359; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_360; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_361; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_362; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_363; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_364; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_365; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_366; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_367; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_368; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_369; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_370; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_371; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_372; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_373; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_374; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_375; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_376; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_377; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_378; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_379; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_380; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_381; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_382; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_383; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_384; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_385; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_386; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_387; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_388; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_389; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_390; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_391; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_392; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_393; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_394; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_395; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_396; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_397; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_398; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_399; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_400; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_401; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_402; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_403; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_404; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_405; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_406; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_407; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_408; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_409; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_410; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_411; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_412; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_413; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_414; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_415; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_416; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_417; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_418; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_419; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_420; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_421; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_422; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_423; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_424; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_425; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_426; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_427; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_428; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_429; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_430; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_431; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_432; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_433; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_434; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_435; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_436; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_437; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_438; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_439; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_440; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_441; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_442; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_443; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_444; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_445; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_446; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_447; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_448; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_449; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_450; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_451; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_452; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_453; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_454; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_455; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_456; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_457; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_458; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_459; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_460; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_461; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_462; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_463; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_464; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_465; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_466; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_467; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_468; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_469; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_470; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_471; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_472; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_473; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_474; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_475; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_476; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_477; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_478; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_479; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_480; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_481; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_482; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_483; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_484; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_485; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_486; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_487; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_488; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_489; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_490; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_491; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_492; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_493; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_494; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_495; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_496; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_497; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_498; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_499; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_500; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_501; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_502; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_503; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_504; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_505; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_506; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_507; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_508; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_509; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_510; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_511; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_0; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_1; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_2; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_3; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_4; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_5; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_6; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_7; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_8; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_9; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_10; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_11; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_12; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_13; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_14; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_15; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_parse_current_state; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_parse_current_offset; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_in_parse_transition_field; // @[parser_pisa.scala 31:25]
  wire [3:0] mau_3_io_pipe_phv_in_next_processor_id; // @[parser_pisa.scala 31:25]
  wire  mau_3_io_pipe_phv_in_next_config_id; // @[parser_pisa.scala 31:25]
  wire  mau_3_io_pipe_phv_in_is_valid_processor; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_0; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_1; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_2; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_3; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_4; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_5; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_6; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_7; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_8; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_9; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_10; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_11; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_12; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_13; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_14; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_15; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_16; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_17; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_18; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_19; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_20; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_21; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_22; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_23; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_24; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_25; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_26; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_27; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_28; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_29; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_30; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_31; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_32; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_33; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_34; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_35; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_36; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_37; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_38; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_39; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_40; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_41; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_42; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_43; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_44; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_45; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_46; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_47; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_48; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_49; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_50; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_51; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_52; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_53; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_54; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_55; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_56; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_57; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_58; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_59; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_60; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_61; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_62; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_63; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_64; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_65; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_66; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_67; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_68; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_69; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_70; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_71; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_72; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_73; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_74; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_75; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_76; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_77; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_78; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_79; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_80; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_81; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_82; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_83; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_84; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_85; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_86; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_87; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_88; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_89; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_90; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_91; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_92; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_93; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_94; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_95; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_96; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_97; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_98; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_99; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_100; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_101; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_102; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_103; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_104; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_105; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_106; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_107; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_108; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_109; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_110; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_111; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_112; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_113; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_114; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_115; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_116; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_117; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_118; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_119; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_120; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_121; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_122; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_123; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_124; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_125; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_126; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_127; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_128; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_129; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_130; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_131; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_132; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_133; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_134; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_135; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_136; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_137; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_138; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_139; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_140; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_141; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_142; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_143; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_144; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_145; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_146; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_147; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_148; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_149; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_150; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_151; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_152; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_153; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_154; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_155; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_156; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_157; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_158; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_159; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_160; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_161; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_162; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_163; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_164; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_165; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_166; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_167; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_168; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_169; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_170; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_171; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_172; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_173; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_174; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_175; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_176; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_177; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_178; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_179; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_180; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_181; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_182; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_183; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_184; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_185; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_186; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_187; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_188; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_189; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_190; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_191; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_192; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_193; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_194; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_195; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_196; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_197; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_198; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_199; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_200; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_201; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_202; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_203; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_204; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_205; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_206; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_207; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_208; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_209; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_210; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_211; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_212; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_213; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_214; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_215; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_216; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_217; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_218; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_219; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_220; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_221; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_222; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_223; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_224; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_225; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_226; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_227; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_228; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_229; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_230; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_231; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_232; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_233; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_234; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_235; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_236; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_237; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_238; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_239; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_240; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_241; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_242; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_243; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_244; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_245; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_246; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_247; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_248; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_249; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_250; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_251; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_252; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_253; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_254; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_255; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_256; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_257; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_258; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_259; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_260; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_261; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_262; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_263; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_264; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_265; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_266; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_267; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_268; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_269; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_270; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_271; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_272; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_273; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_274; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_275; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_276; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_277; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_278; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_279; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_280; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_281; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_282; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_283; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_284; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_285; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_286; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_287; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_288; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_289; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_290; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_291; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_292; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_293; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_294; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_295; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_296; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_297; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_298; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_299; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_300; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_301; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_302; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_303; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_304; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_305; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_306; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_307; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_308; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_309; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_310; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_311; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_312; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_313; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_314; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_315; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_316; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_317; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_318; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_319; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_320; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_321; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_322; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_323; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_324; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_325; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_326; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_327; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_328; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_329; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_330; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_331; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_332; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_333; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_334; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_335; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_336; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_337; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_338; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_339; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_340; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_341; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_342; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_343; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_344; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_345; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_346; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_347; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_348; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_349; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_350; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_351; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_352; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_353; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_354; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_355; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_356; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_357; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_358; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_359; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_360; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_361; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_362; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_363; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_364; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_365; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_366; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_367; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_368; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_369; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_370; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_371; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_372; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_373; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_374; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_375; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_376; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_377; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_378; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_379; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_380; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_381; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_382; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_383; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_384; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_385; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_386; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_387; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_388; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_389; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_390; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_391; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_392; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_393; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_394; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_395; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_396; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_397; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_398; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_399; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_400; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_401; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_402; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_403; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_404; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_405; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_406; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_407; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_408; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_409; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_410; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_411; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_412; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_413; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_414; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_415; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_416; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_417; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_418; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_419; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_420; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_421; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_422; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_423; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_424; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_425; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_426; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_427; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_428; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_429; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_430; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_431; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_432; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_433; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_434; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_435; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_436; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_437; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_438; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_439; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_440; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_441; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_442; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_443; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_444; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_445; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_446; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_447; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_448; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_449; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_450; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_451; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_452; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_453; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_454; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_455; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_456; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_457; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_458; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_459; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_460; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_461; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_462; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_463; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_464; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_465; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_466; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_467; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_468; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_469; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_470; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_471; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_472; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_473; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_474; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_475; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_476; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_477; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_478; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_479; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_480; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_481; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_482; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_483; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_484; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_485; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_486; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_487; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_488; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_489; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_490; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_491; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_492; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_493; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_494; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_495; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_496; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_497; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_498; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_499; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_500; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_501; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_502; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_503; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_504; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_505; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_506; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_507; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_508; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_509; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_510; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_511; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_0; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_1; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_2; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_3; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_4; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_5; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_6; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_7; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_8; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_9; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_10; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_11; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_12; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_13; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_14; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_15; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_parse_current_state; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_parse_current_offset; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_out_parse_transition_field; // @[parser_pisa.scala 31:25]
  wire [3:0] mau_3_io_pipe_phv_out_next_processor_id; // @[parser_pisa.scala 31:25]
  wire  mau_3_io_pipe_phv_out_next_config_id; // @[parser_pisa.scala 31:25]
  wire  mau_3_io_pipe_phv_out_is_valid_processor; // @[parser_pisa.scala 31:25]
  wire  mau_3_io_mod_state_id_mod; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_mod_state_id; // @[parser_pisa.scala 31:25]
  wire  mau_3_io_mod_sram_w_cs; // @[parser_pisa.scala 31:25]
  wire  mau_3_io_mod_sram_w_en; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_mod_sram_w_addr; // @[parser_pisa.scala 31:25]
  wire [63:0] mau_3_io_mod_sram_w_data; // @[parser_pisa.scala 31:25]
  wire  mau_4_clock; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_0; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_1; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_2; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_3; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_4; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_5; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_6; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_7; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_8; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_9; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_10; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_11; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_12; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_13; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_14; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_15; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_16; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_17; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_18; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_19; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_20; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_21; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_22; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_23; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_24; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_25; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_26; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_27; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_28; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_29; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_30; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_31; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_32; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_33; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_34; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_35; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_36; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_37; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_38; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_39; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_40; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_41; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_42; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_43; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_44; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_45; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_46; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_47; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_48; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_49; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_50; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_51; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_52; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_53; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_54; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_55; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_56; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_57; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_58; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_59; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_60; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_61; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_62; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_63; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_64; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_65; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_66; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_67; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_68; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_69; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_70; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_71; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_72; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_73; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_74; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_75; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_76; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_77; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_78; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_79; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_80; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_81; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_82; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_83; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_84; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_85; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_86; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_87; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_88; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_89; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_90; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_91; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_92; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_93; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_94; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_95; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_96; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_97; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_98; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_99; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_100; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_101; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_102; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_103; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_104; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_105; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_106; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_107; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_108; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_109; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_110; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_111; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_112; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_113; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_114; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_115; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_116; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_117; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_118; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_119; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_120; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_121; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_122; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_123; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_124; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_125; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_126; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_127; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_128; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_129; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_130; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_131; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_132; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_133; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_134; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_135; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_136; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_137; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_138; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_139; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_140; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_141; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_142; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_143; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_144; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_145; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_146; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_147; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_148; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_149; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_150; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_151; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_152; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_153; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_154; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_155; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_156; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_157; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_158; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_159; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_160; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_161; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_162; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_163; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_164; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_165; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_166; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_167; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_168; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_169; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_170; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_171; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_172; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_173; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_174; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_175; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_176; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_177; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_178; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_179; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_180; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_181; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_182; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_183; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_184; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_185; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_186; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_187; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_188; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_189; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_190; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_191; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_192; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_193; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_194; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_195; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_196; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_197; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_198; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_199; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_200; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_201; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_202; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_203; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_204; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_205; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_206; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_207; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_208; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_209; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_210; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_211; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_212; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_213; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_214; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_215; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_216; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_217; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_218; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_219; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_220; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_221; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_222; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_223; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_224; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_225; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_226; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_227; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_228; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_229; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_230; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_231; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_232; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_233; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_234; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_235; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_236; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_237; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_238; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_239; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_240; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_241; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_242; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_243; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_244; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_245; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_246; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_247; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_248; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_249; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_250; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_251; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_252; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_253; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_254; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_255; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_256; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_257; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_258; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_259; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_260; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_261; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_262; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_263; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_264; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_265; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_266; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_267; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_268; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_269; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_270; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_271; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_272; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_273; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_274; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_275; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_276; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_277; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_278; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_279; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_280; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_281; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_282; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_283; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_284; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_285; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_286; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_287; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_288; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_289; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_290; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_291; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_292; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_293; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_294; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_295; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_296; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_297; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_298; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_299; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_300; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_301; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_302; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_303; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_304; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_305; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_306; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_307; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_308; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_309; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_310; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_311; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_312; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_313; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_314; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_315; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_316; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_317; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_318; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_319; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_320; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_321; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_322; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_323; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_324; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_325; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_326; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_327; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_328; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_329; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_330; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_331; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_332; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_333; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_334; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_335; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_336; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_337; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_338; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_339; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_340; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_341; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_342; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_343; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_344; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_345; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_346; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_347; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_348; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_349; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_350; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_351; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_352; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_353; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_354; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_355; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_356; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_357; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_358; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_359; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_360; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_361; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_362; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_363; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_364; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_365; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_366; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_367; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_368; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_369; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_370; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_371; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_372; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_373; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_374; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_375; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_376; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_377; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_378; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_379; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_380; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_381; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_382; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_383; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_384; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_385; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_386; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_387; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_388; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_389; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_390; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_391; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_392; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_393; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_394; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_395; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_396; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_397; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_398; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_399; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_400; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_401; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_402; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_403; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_404; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_405; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_406; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_407; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_408; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_409; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_410; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_411; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_412; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_413; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_414; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_415; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_416; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_417; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_418; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_419; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_420; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_421; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_422; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_423; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_424; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_425; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_426; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_427; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_428; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_429; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_430; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_431; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_432; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_433; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_434; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_435; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_436; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_437; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_438; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_439; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_440; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_441; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_442; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_443; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_444; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_445; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_446; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_447; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_448; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_449; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_450; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_451; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_452; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_453; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_454; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_455; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_456; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_457; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_458; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_459; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_460; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_461; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_462; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_463; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_464; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_465; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_466; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_467; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_468; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_469; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_470; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_471; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_472; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_473; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_474; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_475; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_476; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_477; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_478; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_479; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_480; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_481; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_482; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_483; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_484; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_485; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_486; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_487; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_488; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_489; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_490; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_491; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_492; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_493; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_494; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_495; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_496; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_497; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_498; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_499; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_500; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_501; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_502; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_503; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_504; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_505; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_506; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_507; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_508; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_509; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_510; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_511; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_in_header_0; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_in_header_1; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_in_header_2; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_in_header_3; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_in_header_4; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_in_header_5; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_in_header_6; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_in_header_7; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_in_header_8; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_in_header_9; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_in_header_10; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_in_header_11; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_in_header_12; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_in_header_13; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_in_header_14; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_in_header_15; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_parse_current_state; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_parse_current_offset; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_in_parse_transition_field; // @[parser_pisa.scala 31:25]
  wire [3:0] mau_4_io_pipe_phv_in_next_processor_id; // @[parser_pisa.scala 31:25]
  wire  mau_4_io_pipe_phv_in_next_config_id; // @[parser_pisa.scala 31:25]
  wire  mau_4_io_pipe_phv_in_is_valid_processor; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_0; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_1; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_2; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_3; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_4; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_5; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_6; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_7; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_8; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_9; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_10; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_11; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_12; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_13; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_14; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_15; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_16; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_17; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_18; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_19; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_20; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_21; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_22; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_23; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_24; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_25; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_26; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_27; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_28; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_29; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_30; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_31; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_32; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_33; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_34; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_35; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_36; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_37; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_38; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_39; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_40; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_41; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_42; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_43; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_44; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_45; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_46; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_47; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_48; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_49; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_50; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_51; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_52; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_53; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_54; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_55; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_56; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_57; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_58; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_59; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_60; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_61; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_62; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_63; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_64; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_65; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_66; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_67; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_68; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_69; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_70; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_71; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_72; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_73; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_74; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_75; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_76; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_77; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_78; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_79; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_80; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_81; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_82; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_83; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_84; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_85; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_86; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_87; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_88; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_89; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_90; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_91; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_92; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_93; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_94; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_95; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_96; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_97; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_98; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_99; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_100; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_101; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_102; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_103; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_104; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_105; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_106; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_107; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_108; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_109; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_110; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_111; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_112; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_113; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_114; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_115; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_116; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_117; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_118; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_119; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_120; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_121; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_122; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_123; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_124; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_125; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_126; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_127; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_128; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_129; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_130; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_131; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_132; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_133; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_134; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_135; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_136; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_137; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_138; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_139; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_140; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_141; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_142; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_143; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_144; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_145; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_146; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_147; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_148; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_149; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_150; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_151; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_152; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_153; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_154; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_155; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_156; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_157; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_158; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_159; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_160; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_161; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_162; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_163; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_164; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_165; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_166; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_167; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_168; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_169; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_170; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_171; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_172; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_173; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_174; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_175; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_176; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_177; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_178; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_179; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_180; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_181; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_182; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_183; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_184; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_185; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_186; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_187; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_188; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_189; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_190; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_191; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_192; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_193; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_194; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_195; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_196; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_197; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_198; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_199; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_200; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_201; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_202; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_203; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_204; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_205; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_206; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_207; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_208; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_209; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_210; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_211; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_212; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_213; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_214; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_215; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_216; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_217; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_218; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_219; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_220; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_221; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_222; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_223; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_224; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_225; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_226; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_227; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_228; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_229; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_230; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_231; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_232; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_233; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_234; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_235; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_236; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_237; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_238; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_239; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_240; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_241; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_242; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_243; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_244; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_245; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_246; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_247; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_248; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_249; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_250; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_251; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_252; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_253; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_254; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_255; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_256; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_257; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_258; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_259; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_260; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_261; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_262; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_263; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_264; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_265; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_266; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_267; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_268; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_269; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_270; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_271; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_272; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_273; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_274; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_275; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_276; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_277; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_278; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_279; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_280; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_281; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_282; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_283; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_284; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_285; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_286; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_287; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_288; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_289; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_290; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_291; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_292; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_293; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_294; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_295; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_296; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_297; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_298; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_299; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_300; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_301; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_302; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_303; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_304; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_305; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_306; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_307; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_308; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_309; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_310; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_311; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_312; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_313; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_314; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_315; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_316; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_317; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_318; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_319; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_320; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_321; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_322; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_323; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_324; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_325; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_326; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_327; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_328; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_329; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_330; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_331; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_332; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_333; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_334; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_335; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_336; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_337; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_338; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_339; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_340; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_341; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_342; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_343; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_344; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_345; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_346; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_347; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_348; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_349; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_350; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_351; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_352; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_353; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_354; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_355; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_356; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_357; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_358; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_359; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_360; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_361; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_362; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_363; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_364; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_365; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_366; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_367; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_368; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_369; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_370; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_371; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_372; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_373; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_374; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_375; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_376; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_377; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_378; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_379; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_380; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_381; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_382; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_383; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_384; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_385; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_386; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_387; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_388; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_389; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_390; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_391; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_392; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_393; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_394; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_395; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_396; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_397; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_398; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_399; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_400; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_401; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_402; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_403; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_404; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_405; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_406; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_407; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_408; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_409; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_410; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_411; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_412; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_413; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_414; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_415; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_416; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_417; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_418; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_419; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_420; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_421; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_422; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_423; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_424; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_425; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_426; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_427; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_428; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_429; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_430; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_431; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_432; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_433; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_434; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_435; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_436; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_437; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_438; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_439; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_440; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_441; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_442; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_443; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_444; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_445; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_446; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_447; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_448; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_449; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_450; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_451; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_452; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_453; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_454; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_455; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_456; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_457; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_458; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_459; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_460; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_461; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_462; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_463; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_464; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_465; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_466; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_467; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_468; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_469; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_470; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_471; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_472; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_473; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_474; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_475; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_476; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_477; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_478; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_479; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_480; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_481; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_482; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_483; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_484; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_485; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_486; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_487; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_488; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_489; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_490; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_491; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_492; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_493; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_494; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_495; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_496; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_497; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_498; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_499; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_500; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_501; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_502; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_503; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_504; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_505; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_506; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_507; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_508; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_509; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_510; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_511; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_out_header_0; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_out_header_1; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_out_header_2; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_out_header_3; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_out_header_4; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_out_header_5; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_out_header_6; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_out_header_7; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_out_header_8; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_out_header_9; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_out_header_10; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_out_header_11; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_out_header_12; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_out_header_13; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_out_header_14; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_out_header_15; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_parse_current_state; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_parse_current_offset; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_out_parse_transition_field; // @[parser_pisa.scala 31:25]
  wire [3:0] mau_4_io_pipe_phv_out_next_processor_id; // @[parser_pisa.scala 31:25]
  wire  mau_4_io_pipe_phv_out_next_config_id; // @[parser_pisa.scala 31:25]
  wire  mau_4_io_pipe_phv_out_is_valid_processor; // @[parser_pisa.scala 31:25]
  wire  mau_4_io_mod_state_id_mod; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_mod_state_id; // @[parser_pisa.scala 31:25]
  wire  mau_4_io_mod_sram_w_cs; // @[parser_pisa.scala 31:25]
  wire  mau_4_io_mod_sram_w_en; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_mod_sram_w_addr; // @[parser_pisa.scala 31:25]
  wire [63:0] mau_4_io_mod_sram_w_data; // @[parser_pisa.scala 31:25]
  wire  mau_5_clock; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_0; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_1; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_2; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_3; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_4; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_5; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_6; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_7; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_8; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_9; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_10; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_11; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_12; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_13; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_14; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_15; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_16; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_17; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_18; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_19; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_20; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_21; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_22; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_23; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_24; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_25; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_26; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_27; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_28; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_29; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_30; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_31; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_32; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_33; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_34; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_35; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_36; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_37; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_38; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_39; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_40; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_41; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_42; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_43; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_44; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_45; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_46; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_47; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_48; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_49; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_50; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_51; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_52; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_53; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_54; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_55; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_56; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_57; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_58; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_59; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_60; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_61; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_62; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_63; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_64; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_65; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_66; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_67; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_68; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_69; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_70; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_71; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_72; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_73; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_74; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_75; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_76; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_77; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_78; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_79; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_80; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_81; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_82; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_83; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_84; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_85; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_86; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_87; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_88; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_89; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_90; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_91; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_92; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_93; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_94; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_95; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_96; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_97; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_98; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_99; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_100; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_101; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_102; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_103; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_104; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_105; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_106; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_107; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_108; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_109; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_110; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_111; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_112; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_113; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_114; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_115; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_116; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_117; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_118; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_119; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_120; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_121; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_122; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_123; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_124; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_125; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_126; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_127; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_128; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_129; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_130; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_131; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_132; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_133; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_134; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_135; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_136; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_137; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_138; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_139; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_140; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_141; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_142; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_143; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_144; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_145; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_146; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_147; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_148; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_149; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_150; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_151; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_152; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_153; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_154; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_155; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_156; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_157; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_158; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_159; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_160; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_161; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_162; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_163; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_164; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_165; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_166; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_167; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_168; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_169; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_170; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_171; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_172; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_173; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_174; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_175; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_176; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_177; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_178; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_179; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_180; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_181; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_182; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_183; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_184; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_185; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_186; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_187; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_188; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_189; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_190; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_191; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_192; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_193; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_194; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_195; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_196; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_197; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_198; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_199; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_200; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_201; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_202; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_203; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_204; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_205; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_206; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_207; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_208; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_209; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_210; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_211; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_212; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_213; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_214; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_215; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_216; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_217; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_218; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_219; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_220; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_221; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_222; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_223; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_224; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_225; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_226; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_227; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_228; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_229; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_230; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_231; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_232; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_233; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_234; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_235; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_236; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_237; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_238; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_239; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_240; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_241; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_242; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_243; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_244; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_245; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_246; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_247; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_248; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_249; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_250; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_251; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_252; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_253; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_254; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_255; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_256; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_257; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_258; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_259; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_260; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_261; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_262; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_263; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_264; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_265; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_266; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_267; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_268; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_269; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_270; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_271; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_272; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_273; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_274; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_275; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_276; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_277; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_278; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_279; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_280; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_281; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_282; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_283; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_284; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_285; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_286; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_287; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_288; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_289; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_290; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_291; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_292; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_293; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_294; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_295; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_296; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_297; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_298; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_299; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_300; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_301; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_302; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_303; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_304; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_305; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_306; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_307; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_308; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_309; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_310; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_311; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_312; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_313; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_314; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_315; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_316; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_317; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_318; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_319; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_320; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_321; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_322; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_323; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_324; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_325; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_326; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_327; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_328; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_329; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_330; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_331; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_332; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_333; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_334; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_335; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_336; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_337; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_338; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_339; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_340; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_341; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_342; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_343; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_344; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_345; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_346; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_347; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_348; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_349; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_350; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_351; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_352; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_353; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_354; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_355; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_356; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_357; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_358; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_359; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_360; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_361; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_362; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_363; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_364; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_365; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_366; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_367; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_368; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_369; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_370; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_371; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_372; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_373; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_374; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_375; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_376; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_377; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_378; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_379; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_380; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_381; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_382; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_383; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_384; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_385; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_386; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_387; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_388; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_389; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_390; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_391; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_392; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_393; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_394; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_395; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_396; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_397; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_398; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_399; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_400; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_401; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_402; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_403; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_404; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_405; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_406; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_407; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_408; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_409; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_410; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_411; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_412; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_413; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_414; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_415; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_416; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_417; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_418; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_419; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_420; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_421; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_422; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_423; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_424; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_425; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_426; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_427; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_428; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_429; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_430; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_431; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_432; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_433; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_434; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_435; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_436; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_437; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_438; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_439; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_440; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_441; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_442; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_443; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_444; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_445; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_446; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_447; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_448; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_449; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_450; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_451; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_452; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_453; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_454; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_455; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_456; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_457; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_458; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_459; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_460; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_461; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_462; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_463; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_464; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_465; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_466; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_467; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_468; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_469; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_470; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_471; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_472; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_473; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_474; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_475; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_476; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_477; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_478; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_479; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_480; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_481; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_482; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_483; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_484; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_485; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_486; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_487; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_488; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_489; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_490; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_491; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_492; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_493; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_494; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_495; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_496; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_497; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_498; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_499; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_500; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_501; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_502; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_503; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_504; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_505; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_506; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_507; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_508; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_509; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_510; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_511; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_in_header_0; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_in_header_1; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_in_header_2; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_in_header_3; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_in_header_4; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_in_header_5; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_in_header_6; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_in_header_7; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_in_header_8; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_in_header_9; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_in_header_10; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_in_header_11; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_in_header_12; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_in_header_13; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_in_header_14; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_in_header_15; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_parse_current_state; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_parse_current_offset; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_in_parse_transition_field; // @[parser_pisa.scala 31:25]
  wire [3:0] mau_5_io_pipe_phv_in_next_processor_id; // @[parser_pisa.scala 31:25]
  wire  mau_5_io_pipe_phv_in_next_config_id; // @[parser_pisa.scala 31:25]
  wire  mau_5_io_pipe_phv_in_is_valid_processor; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_0; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_1; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_2; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_3; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_4; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_5; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_6; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_7; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_8; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_9; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_10; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_11; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_12; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_13; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_14; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_15; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_16; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_17; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_18; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_19; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_20; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_21; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_22; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_23; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_24; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_25; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_26; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_27; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_28; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_29; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_30; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_31; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_32; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_33; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_34; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_35; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_36; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_37; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_38; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_39; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_40; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_41; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_42; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_43; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_44; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_45; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_46; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_47; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_48; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_49; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_50; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_51; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_52; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_53; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_54; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_55; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_56; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_57; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_58; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_59; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_60; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_61; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_62; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_63; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_64; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_65; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_66; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_67; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_68; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_69; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_70; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_71; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_72; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_73; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_74; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_75; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_76; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_77; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_78; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_79; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_80; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_81; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_82; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_83; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_84; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_85; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_86; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_87; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_88; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_89; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_90; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_91; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_92; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_93; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_94; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_95; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_96; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_97; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_98; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_99; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_100; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_101; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_102; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_103; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_104; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_105; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_106; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_107; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_108; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_109; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_110; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_111; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_112; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_113; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_114; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_115; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_116; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_117; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_118; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_119; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_120; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_121; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_122; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_123; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_124; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_125; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_126; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_127; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_128; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_129; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_130; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_131; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_132; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_133; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_134; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_135; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_136; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_137; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_138; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_139; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_140; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_141; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_142; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_143; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_144; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_145; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_146; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_147; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_148; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_149; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_150; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_151; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_152; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_153; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_154; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_155; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_156; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_157; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_158; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_159; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_160; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_161; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_162; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_163; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_164; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_165; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_166; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_167; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_168; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_169; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_170; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_171; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_172; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_173; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_174; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_175; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_176; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_177; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_178; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_179; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_180; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_181; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_182; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_183; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_184; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_185; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_186; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_187; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_188; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_189; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_190; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_191; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_192; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_193; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_194; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_195; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_196; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_197; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_198; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_199; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_200; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_201; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_202; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_203; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_204; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_205; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_206; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_207; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_208; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_209; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_210; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_211; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_212; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_213; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_214; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_215; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_216; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_217; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_218; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_219; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_220; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_221; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_222; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_223; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_224; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_225; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_226; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_227; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_228; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_229; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_230; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_231; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_232; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_233; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_234; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_235; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_236; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_237; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_238; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_239; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_240; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_241; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_242; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_243; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_244; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_245; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_246; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_247; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_248; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_249; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_250; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_251; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_252; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_253; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_254; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_255; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_256; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_257; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_258; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_259; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_260; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_261; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_262; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_263; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_264; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_265; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_266; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_267; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_268; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_269; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_270; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_271; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_272; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_273; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_274; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_275; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_276; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_277; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_278; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_279; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_280; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_281; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_282; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_283; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_284; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_285; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_286; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_287; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_288; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_289; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_290; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_291; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_292; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_293; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_294; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_295; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_296; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_297; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_298; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_299; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_300; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_301; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_302; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_303; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_304; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_305; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_306; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_307; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_308; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_309; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_310; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_311; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_312; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_313; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_314; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_315; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_316; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_317; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_318; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_319; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_320; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_321; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_322; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_323; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_324; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_325; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_326; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_327; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_328; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_329; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_330; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_331; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_332; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_333; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_334; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_335; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_336; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_337; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_338; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_339; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_340; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_341; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_342; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_343; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_344; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_345; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_346; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_347; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_348; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_349; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_350; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_351; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_352; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_353; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_354; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_355; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_356; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_357; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_358; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_359; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_360; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_361; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_362; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_363; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_364; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_365; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_366; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_367; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_368; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_369; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_370; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_371; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_372; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_373; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_374; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_375; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_376; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_377; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_378; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_379; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_380; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_381; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_382; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_383; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_384; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_385; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_386; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_387; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_388; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_389; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_390; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_391; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_392; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_393; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_394; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_395; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_396; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_397; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_398; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_399; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_400; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_401; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_402; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_403; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_404; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_405; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_406; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_407; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_408; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_409; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_410; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_411; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_412; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_413; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_414; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_415; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_416; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_417; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_418; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_419; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_420; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_421; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_422; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_423; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_424; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_425; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_426; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_427; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_428; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_429; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_430; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_431; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_432; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_433; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_434; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_435; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_436; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_437; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_438; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_439; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_440; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_441; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_442; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_443; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_444; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_445; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_446; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_447; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_448; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_449; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_450; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_451; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_452; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_453; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_454; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_455; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_456; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_457; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_458; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_459; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_460; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_461; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_462; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_463; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_464; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_465; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_466; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_467; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_468; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_469; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_470; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_471; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_472; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_473; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_474; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_475; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_476; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_477; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_478; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_479; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_480; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_481; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_482; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_483; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_484; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_485; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_486; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_487; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_488; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_489; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_490; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_491; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_492; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_493; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_494; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_495; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_496; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_497; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_498; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_499; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_500; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_501; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_502; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_503; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_504; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_505; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_506; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_507; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_508; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_509; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_510; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_511; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_out_header_0; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_out_header_1; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_out_header_2; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_out_header_3; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_out_header_4; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_out_header_5; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_out_header_6; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_out_header_7; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_out_header_8; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_out_header_9; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_out_header_10; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_out_header_11; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_out_header_12; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_out_header_13; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_out_header_14; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_out_header_15; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_parse_current_state; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_parse_current_offset; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_out_parse_transition_field; // @[parser_pisa.scala 31:25]
  wire [3:0] mau_5_io_pipe_phv_out_next_processor_id; // @[parser_pisa.scala 31:25]
  wire  mau_5_io_pipe_phv_out_next_config_id; // @[parser_pisa.scala 31:25]
  wire  mau_5_io_pipe_phv_out_is_valid_processor; // @[parser_pisa.scala 31:25]
  wire  mau_5_io_mod_state_id_mod; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_mod_state_id; // @[parser_pisa.scala 31:25]
  wire  mau_5_io_mod_sram_w_cs; // @[parser_pisa.scala 31:25]
  wire  mau_5_io_mod_sram_w_en; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_mod_sram_w_addr; // @[parser_pisa.scala 31:25]
  wire [63:0] mau_5_io_mod_sram_w_data; // @[parser_pisa.scala 31:25]
  wire  mau_6_clock; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_0; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_1; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_2; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_3; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_4; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_5; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_6; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_7; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_8; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_9; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_10; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_11; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_12; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_13; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_14; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_15; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_16; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_17; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_18; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_19; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_20; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_21; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_22; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_23; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_24; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_25; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_26; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_27; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_28; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_29; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_30; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_31; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_32; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_33; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_34; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_35; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_36; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_37; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_38; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_39; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_40; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_41; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_42; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_43; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_44; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_45; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_46; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_47; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_48; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_49; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_50; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_51; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_52; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_53; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_54; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_55; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_56; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_57; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_58; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_59; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_60; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_61; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_62; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_63; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_64; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_65; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_66; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_67; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_68; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_69; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_70; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_71; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_72; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_73; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_74; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_75; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_76; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_77; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_78; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_79; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_80; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_81; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_82; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_83; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_84; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_85; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_86; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_87; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_88; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_89; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_90; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_91; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_92; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_93; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_94; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_95; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_96; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_97; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_98; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_99; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_100; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_101; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_102; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_103; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_104; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_105; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_106; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_107; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_108; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_109; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_110; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_111; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_112; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_113; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_114; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_115; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_116; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_117; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_118; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_119; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_120; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_121; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_122; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_123; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_124; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_125; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_126; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_127; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_128; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_129; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_130; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_131; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_132; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_133; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_134; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_135; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_136; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_137; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_138; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_139; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_140; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_141; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_142; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_143; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_144; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_145; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_146; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_147; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_148; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_149; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_150; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_151; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_152; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_153; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_154; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_155; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_156; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_157; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_158; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_159; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_160; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_161; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_162; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_163; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_164; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_165; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_166; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_167; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_168; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_169; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_170; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_171; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_172; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_173; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_174; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_175; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_176; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_177; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_178; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_179; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_180; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_181; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_182; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_183; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_184; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_185; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_186; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_187; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_188; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_189; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_190; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_191; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_192; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_193; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_194; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_195; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_196; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_197; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_198; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_199; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_200; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_201; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_202; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_203; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_204; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_205; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_206; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_207; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_208; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_209; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_210; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_211; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_212; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_213; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_214; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_215; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_216; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_217; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_218; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_219; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_220; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_221; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_222; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_223; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_224; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_225; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_226; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_227; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_228; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_229; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_230; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_231; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_232; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_233; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_234; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_235; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_236; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_237; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_238; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_239; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_240; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_241; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_242; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_243; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_244; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_245; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_246; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_247; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_248; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_249; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_250; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_251; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_252; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_253; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_254; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_255; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_256; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_257; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_258; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_259; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_260; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_261; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_262; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_263; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_264; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_265; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_266; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_267; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_268; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_269; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_270; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_271; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_272; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_273; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_274; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_275; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_276; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_277; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_278; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_279; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_280; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_281; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_282; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_283; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_284; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_285; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_286; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_287; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_288; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_289; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_290; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_291; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_292; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_293; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_294; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_295; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_296; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_297; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_298; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_299; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_300; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_301; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_302; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_303; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_304; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_305; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_306; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_307; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_308; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_309; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_310; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_311; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_312; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_313; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_314; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_315; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_316; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_317; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_318; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_319; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_320; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_321; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_322; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_323; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_324; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_325; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_326; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_327; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_328; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_329; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_330; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_331; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_332; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_333; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_334; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_335; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_336; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_337; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_338; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_339; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_340; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_341; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_342; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_343; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_344; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_345; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_346; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_347; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_348; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_349; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_350; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_351; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_352; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_353; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_354; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_355; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_356; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_357; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_358; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_359; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_360; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_361; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_362; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_363; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_364; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_365; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_366; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_367; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_368; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_369; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_370; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_371; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_372; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_373; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_374; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_375; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_376; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_377; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_378; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_379; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_380; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_381; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_382; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_383; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_384; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_385; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_386; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_387; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_388; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_389; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_390; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_391; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_392; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_393; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_394; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_395; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_396; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_397; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_398; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_399; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_400; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_401; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_402; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_403; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_404; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_405; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_406; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_407; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_408; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_409; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_410; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_411; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_412; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_413; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_414; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_415; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_416; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_417; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_418; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_419; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_420; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_421; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_422; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_423; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_424; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_425; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_426; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_427; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_428; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_429; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_430; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_431; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_432; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_433; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_434; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_435; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_436; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_437; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_438; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_439; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_440; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_441; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_442; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_443; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_444; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_445; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_446; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_447; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_448; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_449; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_450; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_451; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_452; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_453; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_454; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_455; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_456; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_457; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_458; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_459; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_460; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_461; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_462; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_463; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_464; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_465; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_466; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_467; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_468; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_469; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_470; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_471; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_472; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_473; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_474; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_475; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_476; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_477; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_478; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_479; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_480; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_481; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_482; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_483; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_484; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_485; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_486; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_487; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_488; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_489; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_490; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_491; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_492; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_493; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_494; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_495; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_496; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_497; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_498; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_499; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_500; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_501; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_502; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_503; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_504; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_505; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_506; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_507; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_508; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_509; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_510; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_511; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_in_header_0; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_in_header_1; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_in_header_2; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_in_header_3; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_in_header_4; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_in_header_5; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_in_header_6; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_in_header_7; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_in_header_8; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_in_header_9; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_in_header_10; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_in_header_11; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_in_header_12; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_in_header_13; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_in_header_14; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_in_header_15; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_parse_current_state; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_parse_current_offset; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_in_parse_transition_field; // @[parser_pisa.scala 31:25]
  wire [3:0] mau_6_io_pipe_phv_in_next_processor_id; // @[parser_pisa.scala 31:25]
  wire  mau_6_io_pipe_phv_in_next_config_id; // @[parser_pisa.scala 31:25]
  wire  mau_6_io_pipe_phv_in_is_valid_processor; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_0; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_1; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_2; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_3; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_4; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_5; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_6; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_7; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_8; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_9; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_10; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_11; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_12; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_13; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_14; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_15; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_16; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_17; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_18; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_19; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_20; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_21; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_22; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_23; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_24; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_25; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_26; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_27; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_28; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_29; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_30; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_31; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_32; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_33; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_34; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_35; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_36; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_37; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_38; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_39; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_40; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_41; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_42; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_43; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_44; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_45; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_46; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_47; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_48; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_49; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_50; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_51; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_52; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_53; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_54; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_55; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_56; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_57; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_58; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_59; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_60; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_61; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_62; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_63; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_64; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_65; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_66; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_67; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_68; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_69; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_70; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_71; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_72; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_73; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_74; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_75; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_76; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_77; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_78; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_79; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_80; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_81; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_82; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_83; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_84; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_85; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_86; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_87; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_88; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_89; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_90; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_91; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_92; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_93; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_94; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_95; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_96; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_97; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_98; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_99; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_100; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_101; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_102; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_103; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_104; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_105; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_106; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_107; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_108; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_109; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_110; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_111; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_112; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_113; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_114; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_115; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_116; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_117; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_118; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_119; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_120; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_121; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_122; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_123; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_124; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_125; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_126; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_127; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_128; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_129; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_130; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_131; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_132; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_133; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_134; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_135; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_136; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_137; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_138; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_139; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_140; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_141; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_142; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_143; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_144; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_145; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_146; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_147; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_148; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_149; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_150; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_151; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_152; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_153; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_154; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_155; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_156; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_157; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_158; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_159; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_160; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_161; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_162; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_163; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_164; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_165; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_166; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_167; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_168; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_169; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_170; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_171; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_172; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_173; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_174; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_175; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_176; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_177; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_178; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_179; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_180; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_181; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_182; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_183; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_184; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_185; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_186; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_187; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_188; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_189; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_190; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_191; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_192; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_193; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_194; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_195; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_196; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_197; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_198; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_199; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_200; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_201; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_202; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_203; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_204; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_205; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_206; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_207; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_208; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_209; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_210; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_211; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_212; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_213; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_214; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_215; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_216; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_217; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_218; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_219; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_220; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_221; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_222; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_223; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_224; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_225; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_226; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_227; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_228; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_229; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_230; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_231; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_232; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_233; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_234; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_235; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_236; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_237; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_238; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_239; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_240; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_241; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_242; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_243; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_244; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_245; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_246; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_247; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_248; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_249; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_250; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_251; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_252; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_253; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_254; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_255; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_256; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_257; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_258; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_259; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_260; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_261; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_262; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_263; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_264; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_265; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_266; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_267; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_268; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_269; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_270; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_271; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_272; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_273; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_274; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_275; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_276; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_277; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_278; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_279; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_280; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_281; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_282; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_283; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_284; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_285; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_286; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_287; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_288; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_289; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_290; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_291; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_292; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_293; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_294; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_295; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_296; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_297; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_298; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_299; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_300; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_301; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_302; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_303; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_304; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_305; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_306; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_307; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_308; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_309; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_310; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_311; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_312; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_313; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_314; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_315; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_316; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_317; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_318; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_319; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_320; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_321; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_322; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_323; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_324; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_325; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_326; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_327; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_328; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_329; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_330; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_331; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_332; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_333; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_334; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_335; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_336; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_337; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_338; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_339; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_340; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_341; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_342; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_343; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_344; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_345; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_346; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_347; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_348; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_349; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_350; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_351; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_352; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_353; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_354; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_355; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_356; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_357; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_358; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_359; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_360; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_361; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_362; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_363; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_364; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_365; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_366; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_367; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_368; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_369; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_370; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_371; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_372; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_373; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_374; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_375; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_376; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_377; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_378; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_379; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_380; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_381; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_382; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_383; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_384; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_385; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_386; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_387; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_388; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_389; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_390; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_391; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_392; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_393; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_394; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_395; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_396; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_397; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_398; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_399; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_400; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_401; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_402; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_403; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_404; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_405; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_406; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_407; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_408; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_409; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_410; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_411; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_412; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_413; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_414; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_415; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_416; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_417; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_418; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_419; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_420; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_421; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_422; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_423; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_424; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_425; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_426; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_427; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_428; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_429; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_430; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_431; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_432; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_433; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_434; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_435; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_436; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_437; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_438; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_439; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_440; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_441; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_442; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_443; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_444; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_445; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_446; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_447; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_448; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_449; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_450; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_451; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_452; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_453; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_454; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_455; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_456; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_457; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_458; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_459; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_460; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_461; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_462; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_463; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_464; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_465; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_466; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_467; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_468; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_469; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_470; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_471; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_472; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_473; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_474; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_475; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_476; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_477; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_478; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_479; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_480; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_481; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_482; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_483; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_484; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_485; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_486; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_487; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_488; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_489; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_490; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_491; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_492; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_493; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_494; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_495; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_496; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_497; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_498; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_499; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_500; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_501; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_502; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_503; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_504; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_505; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_506; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_507; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_508; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_509; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_510; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_511; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_out_header_0; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_out_header_1; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_out_header_2; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_out_header_3; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_out_header_4; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_out_header_5; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_out_header_6; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_out_header_7; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_out_header_8; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_out_header_9; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_out_header_10; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_out_header_11; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_out_header_12; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_out_header_13; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_out_header_14; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_out_header_15; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_parse_current_state; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_parse_current_offset; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_out_parse_transition_field; // @[parser_pisa.scala 31:25]
  wire [3:0] mau_6_io_pipe_phv_out_next_processor_id; // @[parser_pisa.scala 31:25]
  wire  mau_6_io_pipe_phv_out_next_config_id; // @[parser_pisa.scala 31:25]
  wire  mau_6_io_pipe_phv_out_is_valid_processor; // @[parser_pisa.scala 31:25]
  wire  mau_6_io_mod_state_id_mod; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_mod_state_id; // @[parser_pisa.scala 31:25]
  wire  mau_6_io_mod_sram_w_cs; // @[parser_pisa.scala 31:25]
  wire  mau_6_io_mod_sram_w_en; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_mod_sram_w_addr; // @[parser_pisa.scala 31:25]
  wire [63:0] mau_6_io_mod_sram_w_data; // @[parser_pisa.scala 31:25]
  wire  mau_7_clock; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_0; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_1; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_2; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_3; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_4; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_5; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_6; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_7; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_8; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_9; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_10; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_11; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_12; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_13; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_14; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_15; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_16; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_17; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_18; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_19; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_20; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_21; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_22; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_23; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_24; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_25; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_26; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_27; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_28; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_29; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_30; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_31; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_32; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_33; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_34; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_35; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_36; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_37; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_38; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_39; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_40; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_41; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_42; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_43; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_44; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_45; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_46; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_47; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_48; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_49; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_50; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_51; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_52; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_53; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_54; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_55; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_56; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_57; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_58; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_59; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_60; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_61; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_62; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_63; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_64; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_65; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_66; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_67; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_68; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_69; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_70; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_71; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_72; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_73; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_74; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_75; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_76; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_77; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_78; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_79; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_80; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_81; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_82; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_83; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_84; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_85; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_86; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_87; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_88; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_89; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_90; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_91; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_92; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_93; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_94; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_95; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_96; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_97; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_98; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_99; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_100; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_101; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_102; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_103; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_104; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_105; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_106; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_107; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_108; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_109; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_110; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_111; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_112; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_113; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_114; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_115; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_116; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_117; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_118; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_119; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_120; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_121; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_122; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_123; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_124; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_125; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_126; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_127; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_128; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_129; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_130; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_131; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_132; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_133; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_134; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_135; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_136; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_137; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_138; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_139; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_140; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_141; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_142; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_143; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_144; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_145; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_146; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_147; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_148; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_149; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_150; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_151; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_152; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_153; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_154; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_155; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_156; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_157; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_158; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_159; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_160; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_161; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_162; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_163; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_164; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_165; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_166; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_167; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_168; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_169; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_170; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_171; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_172; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_173; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_174; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_175; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_176; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_177; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_178; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_179; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_180; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_181; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_182; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_183; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_184; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_185; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_186; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_187; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_188; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_189; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_190; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_191; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_192; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_193; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_194; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_195; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_196; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_197; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_198; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_199; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_200; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_201; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_202; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_203; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_204; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_205; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_206; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_207; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_208; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_209; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_210; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_211; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_212; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_213; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_214; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_215; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_216; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_217; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_218; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_219; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_220; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_221; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_222; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_223; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_224; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_225; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_226; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_227; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_228; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_229; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_230; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_231; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_232; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_233; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_234; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_235; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_236; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_237; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_238; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_239; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_240; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_241; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_242; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_243; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_244; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_245; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_246; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_247; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_248; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_249; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_250; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_251; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_252; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_253; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_254; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_255; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_256; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_257; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_258; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_259; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_260; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_261; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_262; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_263; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_264; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_265; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_266; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_267; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_268; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_269; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_270; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_271; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_272; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_273; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_274; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_275; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_276; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_277; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_278; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_279; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_280; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_281; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_282; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_283; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_284; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_285; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_286; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_287; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_288; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_289; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_290; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_291; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_292; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_293; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_294; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_295; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_296; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_297; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_298; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_299; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_300; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_301; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_302; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_303; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_304; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_305; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_306; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_307; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_308; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_309; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_310; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_311; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_312; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_313; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_314; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_315; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_316; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_317; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_318; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_319; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_320; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_321; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_322; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_323; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_324; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_325; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_326; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_327; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_328; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_329; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_330; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_331; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_332; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_333; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_334; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_335; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_336; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_337; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_338; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_339; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_340; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_341; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_342; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_343; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_344; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_345; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_346; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_347; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_348; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_349; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_350; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_351; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_352; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_353; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_354; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_355; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_356; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_357; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_358; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_359; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_360; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_361; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_362; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_363; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_364; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_365; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_366; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_367; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_368; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_369; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_370; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_371; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_372; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_373; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_374; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_375; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_376; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_377; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_378; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_379; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_380; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_381; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_382; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_383; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_384; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_385; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_386; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_387; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_388; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_389; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_390; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_391; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_392; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_393; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_394; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_395; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_396; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_397; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_398; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_399; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_400; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_401; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_402; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_403; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_404; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_405; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_406; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_407; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_408; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_409; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_410; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_411; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_412; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_413; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_414; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_415; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_416; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_417; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_418; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_419; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_420; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_421; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_422; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_423; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_424; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_425; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_426; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_427; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_428; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_429; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_430; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_431; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_432; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_433; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_434; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_435; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_436; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_437; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_438; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_439; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_440; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_441; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_442; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_443; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_444; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_445; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_446; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_447; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_448; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_449; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_450; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_451; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_452; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_453; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_454; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_455; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_456; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_457; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_458; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_459; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_460; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_461; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_462; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_463; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_464; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_465; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_466; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_467; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_468; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_469; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_470; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_471; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_472; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_473; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_474; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_475; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_476; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_477; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_478; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_479; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_480; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_481; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_482; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_483; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_484; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_485; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_486; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_487; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_488; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_489; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_490; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_491; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_492; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_493; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_494; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_495; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_496; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_497; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_498; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_499; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_500; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_501; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_502; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_503; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_504; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_505; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_506; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_507; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_508; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_509; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_510; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_511; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_in_header_0; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_in_header_1; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_in_header_2; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_in_header_3; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_in_header_4; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_in_header_5; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_in_header_6; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_in_header_7; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_in_header_8; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_in_header_9; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_in_header_10; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_in_header_11; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_in_header_12; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_in_header_13; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_in_header_14; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_in_header_15; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_parse_current_state; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_parse_current_offset; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_in_parse_transition_field; // @[parser_pisa.scala 31:25]
  wire [3:0] mau_7_io_pipe_phv_in_next_processor_id; // @[parser_pisa.scala 31:25]
  wire  mau_7_io_pipe_phv_in_next_config_id; // @[parser_pisa.scala 31:25]
  wire  mau_7_io_pipe_phv_in_is_valid_processor; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_0; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_1; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_2; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_3; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_4; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_5; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_6; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_7; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_8; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_9; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_10; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_11; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_12; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_13; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_14; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_15; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_16; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_17; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_18; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_19; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_20; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_21; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_22; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_23; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_24; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_25; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_26; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_27; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_28; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_29; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_30; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_31; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_32; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_33; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_34; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_35; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_36; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_37; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_38; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_39; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_40; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_41; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_42; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_43; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_44; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_45; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_46; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_47; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_48; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_49; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_50; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_51; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_52; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_53; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_54; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_55; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_56; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_57; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_58; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_59; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_60; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_61; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_62; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_63; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_64; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_65; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_66; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_67; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_68; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_69; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_70; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_71; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_72; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_73; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_74; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_75; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_76; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_77; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_78; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_79; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_80; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_81; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_82; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_83; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_84; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_85; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_86; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_87; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_88; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_89; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_90; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_91; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_92; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_93; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_94; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_95; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_96; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_97; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_98; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_99; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_100; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_101; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_102; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_103; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_104; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_105; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_106; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_107; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_108; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_109; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_110; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_111; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_112; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_113; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_114; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_115; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_116; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_117; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_118; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_119; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_120; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_121; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_122; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_123; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_124; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_125; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_126; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_127; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_128; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_129; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_130; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_131; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_132; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_133; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_134; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_135; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_136; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_137; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_138; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_139; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_140; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_141; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_142; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_143; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_144; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_145; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_146; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_147; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_148; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_149; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_150; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_151; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_152; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_153; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_154; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_155; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_156; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_157; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_158; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_159; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_160; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_161; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_162; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_163; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_164; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_165; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_166; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_167; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_168; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_169; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_170; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_171; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_172; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_173; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_174; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_175; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_176; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_177; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_178; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_179; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_180; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_181; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_182; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_183; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_184; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_185; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_186; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_187; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_188; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_189; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_190; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_191; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_192; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_193; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_194; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_195; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_196; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_197; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_198; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_199; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_200; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_201; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_202; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_203; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_204; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_205; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_206; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_207; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_208; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_209; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_210; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_211; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_212; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_213; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_214; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_215; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_216; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_217; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_218; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_219; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_220; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_221; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_222; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_223; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_224; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_225; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_226; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_227; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_228; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_229; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_230; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_231; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_232; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_233; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_234; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_235; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_236; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_237; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_238; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_239; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_240; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_241; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_242; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_243; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_244; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_245; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_246; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_247; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_248; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_249; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_250; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_251; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_252; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_253; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_254; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_255; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_256; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_257; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_258; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_259; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_260; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_261; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_262; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_263; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_264; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_265; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_266; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_267; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_268; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_269; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_270; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_271; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_272; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_273; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_274; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_275; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_276; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_277; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_278; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_279; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_280; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_281; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_282; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_283; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_284; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_285; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_286; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_287; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_288; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_289; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_290; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_291; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_292; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_293; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_294; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_295; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_296; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_297; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_298; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_299; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_300; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_301; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_302; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_303; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_304; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_305; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_306; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_307; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_308; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_309; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_310; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_311; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_312; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_313; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_314; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_315; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_316; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_317; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_318; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_319; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_320; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_321; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_322; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_323; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_324; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_325; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_326; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_327; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_328; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_329; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_330; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_331; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_332; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_333; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_334; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_335; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_336; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_337; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_338; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_339; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_340; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_341; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_342; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_343; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_344; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_345; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_346; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_347; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_348; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_349; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_350; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_351; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_352; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_353; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_354; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_355; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_356; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_357; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_358; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_359; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_360; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_361; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_362; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_363; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_364; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_365; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_366; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_367; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_368; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_369; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_370; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_371; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_372; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_373; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_374; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_375; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_376; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_377; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_378; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_379; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_380; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_381; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_382; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_383; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_384; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_385; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_386; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_387; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_388; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_389; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_390; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_391; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_392; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_393; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_394; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_395; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_396; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_397; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_398; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_399; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_400; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_401; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_402; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_403; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_404; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_405; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_406; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_407; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_408; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_409; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_410; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_411; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_412; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_413; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_414; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_415; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_416; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_417; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_418; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_419; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_420; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_421; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_422; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_423; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_424; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_425; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_426; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_427; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_428; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_429; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_430; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_431; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_432; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_433; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_434; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_435; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_436; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_437; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_438; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_439; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_440; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_441; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_442; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_443; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_444; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_445; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_446; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_447; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_448; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_449; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_450; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_451; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_452; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_453; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_454; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_455; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_456; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_457; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_458; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_459; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_460; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_461; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_462; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_463; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_464; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_465; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_466; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_467; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_468; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_469; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_470; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_471; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_472; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_473; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_474; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_475; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_476; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_477; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_478; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_479; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_480; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_481; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_482; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_483; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_484; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_485; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_486; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_487; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_488; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_489; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_490; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_491; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_492; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_493; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_494; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_495; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_496; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_497; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_498; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_499; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_500; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_501; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_502; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_503; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_504; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_505; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_506; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_507; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_508; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_509; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_510; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_511; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_out_header_0; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_out_header_1; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_out_header_2; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_out_header_3; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_out_header_4; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_out_header_5; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_out_header_6; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_out_header_7; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_out_header_8; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_out_header_9; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_out_header_10; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_out_header_11; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_out_header_12; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_out_header_13; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_out_header_14; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_out_header_15; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_parse_current_state; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_parse_current_offset; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_out_parse_transition_field; // @[parser_pisa.scala 31:25]
  wire [3:0] mau_7_io_pipe_phv_out_next_processor_id; // @[parser_pisa.scala 31:25]
  wire  mau_7_io_pipe_phv_out_next_config_id; // @[parser_pisa.scala 31:25]
  wire  mau_7_io_pipe_phv_out_is_valid_processor; // @[parser_pisa.scala 31:25]
  wire  mau_7_io_mod_state_id_mod; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_mod_state_id; // @[parser_pisa.scala 31:25]
  wire  mau_7_io_mod_sram_w_cs; // @[parser_pisa.scala 31:25]
  wire  mau_7_io_mod_sram_w_en; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_mod_sram_w_addr; // @[parser_pisa.scala 31:25]
  wire [63:0] mau_7_io_mod_sram_w_data; // @[parser_pisa.scala 31:25]
  reg [3:0] last_mau_id; // @[parser_pisa.scala 24:26]
  wire  _GEN_1 = 4'h1 == last_mau_id & mau_1_io_pipe_phv_out_next_config_id; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [3:0] _GEN_2 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_next_processor_id : 4'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_22 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_0 : io_pipe_phv_in_data_0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_23 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_1 : io_pipe_phv_in_data_1; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_24 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_2 : io_pipe_phv_in_data_2; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_25 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_3 : io_pipe_phv_in_data_3; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_26 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_4 : io_pipe_phv_in_data_4; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_27 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_5 : io_pipe_phv_in_data_5; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_28 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_6 : io_pipe_phv_in_data_6; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_29 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_7 : io_pipe_phv_in_data_7; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_30 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_8 : io_pipe_phv_in_data_8; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_31 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_9 : io_pipe_phv_in_data_9; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_32 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_10 : io_pipe_phv_in_data_10; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_33 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_11 : io_pipe_phv_in_data_11; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_34 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_12 : io_pipe_phv_in_data_12; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_35 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_13 : io_pipe_phv_in_data_13; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_36 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_14 : io_pipe_phv_in_data_14; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_37 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_15 : io_pipe_phv_in_data_15; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_38 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_16 : io_pipe_phv_in_data_16; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_39 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_17 : io_pipe_phv_in_data_17; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_40 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_18 : io_pipe_phv_in_data_18; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_41 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_19 : io_pipe_phv_in_data_19; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_42 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_20 : io_pipe_phv_in_data_20; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_43 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_21 : io_pipe_phv_in_data_21; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_44 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_22 : io_pipe_phv_in_data_22; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_45 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_23 : io_pipe_phv_in_data_23; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_46 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_24 : io_pipe_phv_in_data_24; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_47 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_25 : io_pipe_phv_in_data_25; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_48 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_26 : io_pipe_phv_in_data_26; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_49 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_27 : io_pipe_phv_in_data_27; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_50 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_28 : io_pipe_phv_in_data_28; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_51 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_29 : io_pipe_phv_in_data_29; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_52 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_30 : io_pipe_phv_in_data_30; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_53 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_31 : io_pipe_phv_in_data_31; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_54 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_32 : io_pipe_phv_in_data_32; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_55 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_33 : io_pipe_phv_in_data_33; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_56 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_34 : io_pipe_phv_in_data_34; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_57 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_35 : io_pipe_phv_in_data_35; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_58 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_36 : io_pipe_phv_in_data_36; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_59 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_37 : io_pipe_phv_in_data_37; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_60 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_38 : io_pipe_phv_in_data_38; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_61 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_39 : io_pipe_phv_in_data_39; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_62 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_40 : io_pipe_phv_in_data_40; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_63 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_41 : io_pipe_phv_in_data_41; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_64 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_42 : io_pipe_phv_in_data_42; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_65 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_43 : io_pipe_phv_in_data_43; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_66 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_44 : io_pipe_phv_in_data_44; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_67 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_45 : io_pipe_phv_in_data_45; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_68 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_46 : io_pipe_phv_in_data_46; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_69 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_47 : io_pipe_phv_in_data_47; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_70 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_48 : io_pipe_phv_in_data_48; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_71 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_49 : io_pipe_phv_in_data_49; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_72 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_50 : io_pipe_phv_in_data_50; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_73 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_51 : io_pipe_phv_in_data_51; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_74 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_52 : io_pipe_phv_in_data_52; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_75 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_53 : io_pipe_phv_in_data_53; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_76 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_54 : io_pipe_phv_in_data_54; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_77 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_55 : io_pipe_phv_in_data_55; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_78 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_56 : io_pipe_phv_in_data_56; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_79 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_57 : io_pipe_phv_in_data_57; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_80 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_58 : io_pipe_phv_in_data_58; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_81 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_59 : io_pipe_phv_in_data_59; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_82 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_60 : io_pipe_phv_in_data_60; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_83 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_61 : io_pipe_phv_in_data_61; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_84 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_62 : io_pipe_phv_in_data_62; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_85 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_63 : io_pipe_phv_in_data_63; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_86 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_64 : io_pipe_phv_in_data_64; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_87 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_65 : io_pipe_phv_in_data_65; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_88 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_66 : io_pipe_phv_in_data_66; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_89 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_67 : io_pipe_phv_in_data_67; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_90 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_68 : io_pipe_phv_in_data_68; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_91 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_69 : io_pipe_phv_in_data_69; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_92 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_70 : io_pipe_phv_in_data_70; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_93 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_71 : io_pipe_phv_in_data_71; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_94 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_72 : io_pipe_phv_in_data_72; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_95 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_73 : io_pipe_phv_in_data_73; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_96 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_74 : io_pipe_phv_in_data_74; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_97 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_75 : io_pipe_phv_in_data_75; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_98 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_76 : io_pipe_phv_in_data_76; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_99 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_77 : io_pipe_phv_in_data_77; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_100 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_78 : io_pipe_phv_in_data_78; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_101 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_79 : io_pipe_phv_in_data_79; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_102 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_80 : io_pipe_phv_in_data_80; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_103 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_81 : io_pipe_phv_in_data_81; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_104 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_82 : io_pipe_phv_in_data_82; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_105 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_83 : io_pipe_phv_in_data_83; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_106 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_84 : io_pipe_phv_in_data_84; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_107 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_85 : io_pipe_phv_in_data_85; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_108 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_86 : io_pipe_phv_in_data_86; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_109 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_87 : io_pipe_phv_in_data_87; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_110 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_88 : io_pipe_phv_in_data_88; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_111 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_89 : io_pipe_phv_in_data_89; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_112 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_90 : io_pipe_phv_in_data_90; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_113 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_91 : io_pipe_phv_in_data_91; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_114 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_92 : io_pipe_phv_in_data_92; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_115 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_93 : io_pipe_phv_in_data_93; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_116 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_94 : io_pipe_phv_in_data_94; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_117 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_95 : io_pipe_phv_in_data_95; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_118 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_96 : io_pipe_phv_in_data_96; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_119 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_97 : io_pipe_phv_in_data_97; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_120 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_98 : io_pipe_phv_in_data_98; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_121 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_99 : io_pipe_phv_in_data_99; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_122 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_100 : io_pipe_phv_in_data_100; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_123 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_101 : io_pipe_phv_in_data_101; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_124 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_102 : io_pipe_phv_in_data_102; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_125 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_103 : io_pipe_phv_in_data_103; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_126 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_104 : io_pipe_phv_in_data_104; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_127 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_105 : io_pipe_phv_in_data_105; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_128 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_106 : io_pipe_phv_in_data_106; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_129 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_107 : io_pipe_phv_in_data_107; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_130 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_108 : io_pipe_phv_in_data_108; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_131 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_109 : io_pipe_phv_in_data_109; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_132 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_110 : io_pipe_phv_in_data_110; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_133 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_111 : io_pipe_phv_in_data_111; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_134 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_112 : io_pipe_phv_in_data_112; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_135 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_113 : io_pipe_phv_in_data_113; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_136 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_114 : io_pipe_phv_in_data_114; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_137 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_115 : io_pipe_phv_in_data_115; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_138 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_116 : io_pipe_phv_in_data_116; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_139 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_117 : io_pipe_phv_in_data_117; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_140 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_118 : io_pipe_phv_in_data_118; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_141 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_119 : io_pipe_phv_in_data_119; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_142 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_120 : io_pipe_phv_in_data_120; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_143 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_121 : io_pipe_phv_in_data_121; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_144 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_122 : io_pipe_phv_in_data_122; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_145 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_123 : io_pipe_phv_in_data_123; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_146 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_124 : io_pipe_phv_in_data_124; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_147 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_125 : io_pipe_phv_in_data_125; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_148 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_126 : io_pipe_phv_in_data_126; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_149 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_127 : io_pipe_phv_in_data_127; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_150 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_128 : io_pipe_phv_in_data_128; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_151 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_129 : io_pipe_phv_in_data_129; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_152 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_130 : io_pipe_phv_in_data_130; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_153 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_131 : io_pipe_phv_in_data_131; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_154 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_132 : io_pipe_phv_in_data_132; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_155 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_133 : io_pipe_phv_in_data_133; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_156 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_134 : io_pipe_phv_in_data_134; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_157 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_135 : io_pipe_phv_in_data_135; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_158 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_136 : io_pipe_phv_in_data_136; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_159 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_137 : io_pipe_phv_in_data_137; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_160 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_138 : io_pipe_phv_in_data_138; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_161 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_139 : io_pipe_phv_in_data_139; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_162 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_140 : io_pipe_phv_in_data_140; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_163 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_141 : io_pipe_phv_in_data_141; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_164 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_142 : io_pipe_phv_in_data_142; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_165 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_143 : io_pipe_phv_in_data_143; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_166 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_144 : io_pipe_phv_in_data_144; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_167 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_145 : io_pipe_phv_in_data_145; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_168 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_146 : io_pipe_phv_in_data_146; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_169 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_147 : io_pipe_phv_in_data_147; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_170 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_148 : io_pipe_phv_in_data_148; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_171 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_149 : io_pipe_phv_in_data_149; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_172 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_150 : io_pipe_phv_in_data_150; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_173 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_151 : io_pipe_phv_in_data_151; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_174 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_152 : io_pipe_phv_in_data_152; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_175 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_153 : io_pipe_phv_in_data_153; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_176 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_154 : io_pipe_phv_in_data_154; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_177 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_155 : io_pipe_phv_in_data_155; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_178 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_156 : io_pipe_phv_in_data_156; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_179 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_157 : io_pipe_phv_in_data_157; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_180 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_158 : io_pipe_phv_in_data_158; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_181 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_159 : io_pipe_phv_in_data_159; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_182 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_160 : io_pipe_phv_in_data_160; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_183 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_161 : io_pipe_phv_in_data_161; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_184 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_162 : io_pipe_phv_in_data_162; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_185 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_163 : io_pipe_phv_in_data_163; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_186 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_164 : io_pipe_phv_in_data_164; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_187 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_165 : io_pipe_phv_in_data_165; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_188 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_166 : io_pipe_phv_in_data_166; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_189 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_167 : io_pipe_phv_in_data_167; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_190 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_168 : io_pipe_phv_in_data_168; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_191 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_169 : io_pipe_phv_in_data_169; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_192 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_170 : io_pipe_phv_in_data_170; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_193 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_171 : io_pipe_phv_in_data_171; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_194 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_172 : io_pipe_phv_in_data_172; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_195 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_173 : io_pipe_phv_in_data_173; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_196 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_174 : io_pipe_phv_in_data_174; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_197 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_175 : io_pipe_phv_in_data_175; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_198 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_176 : io_pipe_phv_in_data_176; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_199 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_177 : io_pipe_phv_in_data_177; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_200 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_178 : io_pipe_phv_in_data_178; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_201 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_179 : io_pipe_phv_in_data_179; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_202 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_180 : io_pipe_phv_in_data_180; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_203 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_181 : io_pipe_phv_in_data_181; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_204 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_182 : io_pipe_phv_in_data_182; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_205 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_183 : io_pipe_phv_in_data_183; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_206 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_184 : io_pipe_phv_in_data_184; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_207 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_185 : io_pipe_phv_in_data_185; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_208 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_186 : io_pipe_phv_in_data_186; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_209 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_187 : io_pipe_phv_in_data_187; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_210 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_188 : io_pipe_phv_in_data_188; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_211 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_189 : io_pipe_phv_in_data_189; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_212 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_190 : io_pipe_phv_in_data_190; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_213 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_191 : io_pipe_phv_in_data_191; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_214 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_192 : io_pipe_phv_in_data_192; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_215 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_193 : io_pipe_phv_in_data_193; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_216 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_194 : io_pipe_phv_in_data_194; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_217 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_195 : io_pipe_phv_in_data_195; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_218 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_196 : io_pipe_phv_in_data_196; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_219 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_197 : io_pipe_phv_in_data_197; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_220 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_198 : io_pipe_phv_in_data_198; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_221 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_199 : io_pipe_phv_in_data_199; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_222 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_200 : io_pipe_phv_in_data_200; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_223 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_201 : io_pipe_phv_in_data_201; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_224 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_202 : io_pipe_phv_in_data_202; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_225 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_203 : io_pipe_phv_in_data_203; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_226 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_204 : io_pipe_phv_in_data_204; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_227 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_205 : io_pipe_phv_in_data_205; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_228 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_206 : io_pipe_phv_in_data_206; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_229 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_207 : io_pipe_phv_in_data_207; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_230 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_208 : io_pipe_phv_in_data_208; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_231 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_209 : io_pipe_phv_in_data_209; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_232 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_210 : io_pipe_phv_in_data_210; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_233 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_211 : io_pipe_phv_in_data_211; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_234 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_212 : io_pipe_phv_in_data_212; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_235 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_213 : io_pipe_phv_in_data_213; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_236 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_214 : io_pipe_phv_in_data_214; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_237 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_215 : io_pipe_phv_in_data_215; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_238 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_216 : io_pipe_phv_in_data_216; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_239 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_217 : io_pipe_phv_in_data_217; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_240 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_218 : io_pipe_phv_in_data_218; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_241 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_219 : io_pipe_phv_in_data_219; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_242 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_220 : io_pipe_phv_in_data_220; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_243 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_221 : io_pipe_phv_in_data_221; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_244 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_222 : io_pipe_phv_in_data_222; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_245 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_223 : io_pipe_phv_in_data_223; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_246 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_224 : io_pipe_phv_in_data_224; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_247 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_225 : io_pipe_phv_in_data_225; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_248 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_226 : io_pipe_phv_in_data_226; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_249 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_227 : io_pipe_phv_in_data_227; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_250 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_228 : io_pipe_phv_in_data_228; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_251 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_229 : io_pipe_phv_in_data_229; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_252 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_230 : io_pipe_phv_in_data_230; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_253 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_231 : io_pipe_phv_in_data_231; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_254 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_232 : io_pipe_phv_in_data_232; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_255 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_233 : io_pipe_phv_in_data_233; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_256 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_234 : io_pipe_phv_in_data_234; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_257 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_235 : io_pipe_phv_in_data_235; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_258 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_236 : io_pipe_phv_in_data_236; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_259 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_237 : io_pipe_phv_in_data_237; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_260 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_238 : io_pipe_phv_in_data_238; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_261 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_239 : io_pipe_phv_in_data_239; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_262 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_240 : io_pipe_phv_in_data_240; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_263 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_241 : io_pipe_phv_in_data_241; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_264 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_242 : io_pipe_phv_in_data_242; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_265 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_243 : io_pipe_phv_in_data_243; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_266 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_244 : io_pipe_phv_in_data_244; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_267 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_245 : io_pipe_phv_in_data_245; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_268 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_246 : io_pipe_phv_in_data_246; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_269 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_247 : io_pipe_phv_in_data_247; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_270 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_248 : io_pipe_phv_in_data_248; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_271 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_249 : io_pipe_phv_in_data_249; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_272 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_250 : io_pipe_phv_in_data_250; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_273 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_251 : io_pipe_phv_in_data_251; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_274 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_252 : io_pipe_phv_in_data_252; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_275 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_253 : io_pipe_phv_in_data_253; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_276 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_254 : io_pipe_phv_in_data_254; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_277 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_255 : io_pipe_phv_in_data_255; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_278 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_256 : io_pipe_phv_in_data_256; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_279 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_257 : io_pipe_phv_in_data_257; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_280 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_258 : io_pipe_phv_in_data_258; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_281 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_259 : io_pipe_phv_in_data_259; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_282 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_260 : io_pipe_phv_in_data_260; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_283 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_261 : io_pipe_phv_in_data_261; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_284 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_262 : io_pipe_phv_in_data_262; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_285 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_263 : io_pipe_phv_in_data_263; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_286 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_264 : io_pipe_phv_in_data_264; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_287 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_265 : io_pipe_phv_in_data_265; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_288 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_266 : io_pipe_phv_in_data_266; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_289 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_267 : io_pipe_phv_in_data_267; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_290 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_268 : io_pipe_phv_in_data_268; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_291 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_269 : io_pipe_phv_in_data_269; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_292 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_270 : io_pipe_phv_in_data_270; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_293 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_271 : io_pipe_phv_in_data_271; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_294 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_272 : io_pipe_phv_in_data_272; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_295 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_273 : io_pipe_phv_in_data_273; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_296 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_274 : io_pipe_phv_in_data_274; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_297 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_275 : io_pipe_phv_in_data_275; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_298 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_276 : io_pipe_phv_in_data_276; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_299 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_277 : io_pipe_phv_in_data_277; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_300 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_278 : io_pipe_phv_in_data_278; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_301 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_279 : io_pipe_phv_in_data_279; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_302 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_280 : io_pipe_phv_in_data_280; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_303 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_281 : io_pipe_phv_in_data_281; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_304 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_282 : io_pipe_phv_in_data_282; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_305 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_283 : io_pipe_phv_in_data_283; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_306 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_284 : io_pipe_phv_in_data_284; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_307 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_285 : io_pipe_phv_in_data_285; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_308 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_286 : io_pipe_phv_in_data_286; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_309 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_287 : io_pipe_phv_in_data_287; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_310 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_288 : io_pipe_phv_in_data_288; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_311 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_289 : io_pipe_phv_in_data_289; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_312 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_290 : io_pipe_phv_in_data_290; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_313 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_291 : io_pipe_phv_in_data_291; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_314 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_292 : io_pipe_phv_in_data_292; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_315 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_293 : io_pipe_phv_in_data_293; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_316 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_294 : io_pipe_phv_in_data_294; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_317 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_295 : io_pipe_phv_in_data_295; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_318 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_296 : io_pipe_phv_in_data_296; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_319 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_297 : io_pipe_phv_in_data_297; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_320 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_298 : io_pipe_phv_in_data_298; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_321 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_299 : io_pipe_phv_in_data_299; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_322 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_300 : io_pipe_phv_in_data_300; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_323 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_301 : io_pipe_phv_in_data_301; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_324 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_302 : io_pipe_phv_in_data_302; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_325 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_303 : io_pipe_phv_in_data_303; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_326 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_304 : io_pipe_phv_in_data_304; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_327 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_305 : io_pipe_phv_in_data_305; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_328 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_306 : io_pipe_phv_in_data_306; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_329 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_307 : io_pipe_phv_in_data_307; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_330 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_308 : io_pipe_phv_in_data_308; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_331 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_309 : io_pipe_phv_in_data_309; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_332 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_310 : io_pipe_phv_in_data_310; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_333 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_311 : io_pipe_phv_in_data_311; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_334 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_312 : io_pipe_phv_in_data_312; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_335 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_313 : io_pipe_phv_in_data_313; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_336 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_314 : io_pipe_phv_in_data_314; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_337 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_315 : io_pipe_phv_in_data_315; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_338 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_316 : io_pipe_phv_in_data_316; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_339 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_317 : io_pipe_phv_in_data_317; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_340 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_318 : io_pipe_phv_in_data_318; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_341 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_319 : io_pipe_phv_in_data_319; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_342 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_320 : io_pipe_phv_in_data_320; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_343 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_321 : io_pipe_phv_in_data_321; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_344 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_322 : io_pipe_phv_in_data_322; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_345 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_323 : io_pipe_phv_in_data_323; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_346 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_324 : io_pipe_phv_in_data_324; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_347 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_325 : io_pipe_phv_in_data_325; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_348 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_326 : io_pipe_phv_in_data_326; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_349 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_327 : io_pipe_phv_in_data_327; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_350 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_328 : io_pipe_phv_in_data_328; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_351 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_329 : io_pipe_phv_in_data_329; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_352 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_330 : io_pipe_phv_in_data_330; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_353 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_331 : io_pipe_phv_in_data_331; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_354 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_332 : io_pipe_phv_in_data_332; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_355 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_333 : io_pipe_phv_in_data_333; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_356 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_334 : io_pipe_phv_in_data_334; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_357 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_335 : io_pipe_phv_in_data_335; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_358 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_336 : io_pipe_phv_in_data_336; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_359 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_337 : io_pipe_phv_in_data_337; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_360 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_338 : io_pipe_phv_in_data_338; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_361 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_339 : io_pipe_phv_in_data_339; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_362 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_340 : io_pipe_phv_in_data_340; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_363 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_341 : io_pipe_phv_in_data_341; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_364 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_342 : io_pipe_phv_in_data_342; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_365 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_343 : io_pipe_phv_in_data_343; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_366 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_344 : io_pipe_phv_in_data_344; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_367 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_345 : io_pipe_phv_in_data_345; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_368 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_346 : io_pipe_phv_in_data_346; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_369 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_347 : io_pipe_phv_in_data_347; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_370 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_348 : io_pipe_phv_in_data_348; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_371 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_349 : io_pipe_phv_in_data_349; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_372 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_350 : io_pipe_phv_in_data_350; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_373 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_351 : io_pipe_phv_in_data_351; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_374 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_352 : io_pipe_phv_in_data_352; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_375 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_353 : io_pipe_phv_in_data_353; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_376 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_354 : io_pipe_phv_in_data_354; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_377 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_355 : io_pipe_phv_in_data_355; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_378 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_356 : io_pipe_phv_in_data_356; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_379 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_357 : io_pipe_phv_in_data_357; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_380 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_358 : io_pipe_phv_in_data_358; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_381 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_359 : io_pipe_phv_in_data_359; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_382 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_360 : io_pipe_phv_in_data_360; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_383 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_361 : io_pipe_phv_in_data_361; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_384 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_362 : io_pipe_phv_in_data_362; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_385 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_363 : io_pipe_phv_in_data_363; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_386 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_364 : io_pipe_phv_in_data_364; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_387 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_365 : io_pipe_phv_in_data_365; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_388 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_366 : io_pipe_phv_in_data_366; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_389 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_367 : io_pipe_phv_in_data_367; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_390 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_368 : io_pipe_phv_in_data_368; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_391 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_369 : io_pipe_phv_in_data_369; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_392 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_370 : io_pipe_phv_in_data_370; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_393 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_371 : io_pipe_phv_in_data_371; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_394 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_372 : io_pipe_phv_in_data_372; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_395 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_373 : io_pipe_phv_in_data_373; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_396 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_374 : io_pipe_phv_in_data_374; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_397 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_375 : io_pipe_phv_in_data_375; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_398 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_376 : io_pipe_phv_in_data_376; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_399 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_377 : io_pipe_phv_in_data_377; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_400 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_378 : io_pipe_phv_in_data_378; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_401 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_379 : io_pipe_phv_in_data_379; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_402 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_380 : io_pipe_phv_in_data_380; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_403 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_381 : io_pipe_phv_in_data_381; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_404 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_382 : io_pipe_phv_in_data_382; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_405 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_383 : io_pipe_phv_in_data_383; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_406 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_384 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_407 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_385 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_408 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_386 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_409 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_387 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_410 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_388 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_411 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_389 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_412 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_390 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_413 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_391 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_414 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_392 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_415 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_393 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_416 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_394 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_417 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_395 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_418 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_396 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_419 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_397 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_420 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_398 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_421 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_399 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_422 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_400 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_423 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_401 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_424 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_402 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_425 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_403 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_426 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_404 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_427 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_405 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_428 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_406 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_429 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_407 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_430 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_408 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_431 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_409 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_432 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_410 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_433 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_411 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_434 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_412 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_435 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_413 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_436 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_414 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_437 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_415 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_438 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_416 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_439 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_417 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_440 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_418 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_441 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_419 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_442 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_420 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_443 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_421 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_444 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_422 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_445 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_423 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_446 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_424 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_447 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_425 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_448 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_426 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_449 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_427 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_450 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_428 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_451 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_429 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_452 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_430 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_453 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_431 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_454 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_432 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_455 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_433 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_456 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_434 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_457 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_435 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_458 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_436 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_459 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_437 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_460 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_438 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_461 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_439 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_462 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_440 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_463 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_441 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_464 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_442 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_465 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_443 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_466 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_444 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_467 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_445 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_468 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_446 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_469 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_447 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_470 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_448 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_471 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_449 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_472 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_450 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_473 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_451 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_474 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_452 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_475 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_453 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_476 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_454 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_477 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_455 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_478 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_456 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_479 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_457 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_480 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_458 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_481 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_459 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_482 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_460 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_483 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_461 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_484 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_462 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_485 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_463 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_486 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_464 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_487 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_465 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_488 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_466 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_489 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_467 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_490 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_468 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_491 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_469 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_492 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_470 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_493 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_471 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_494 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_472 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_495 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_473 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_496 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_474 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_497 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_475 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_498 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_476 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_499 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_477 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_500 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_478 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_501 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_479 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_502 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_480 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_503 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_481 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_504 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_482 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_505 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_483 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_506 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_484 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_507 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_485 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_508 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_486 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_509 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_487 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_510 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_488 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_511 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_489 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_512 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_490 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_513 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_491 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_514 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_492 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_515 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_493 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_516 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_494 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_517 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_495 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_518 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_496 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_519 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_497 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_520 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_498 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_521 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_499 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_522 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_500 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_523 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_501 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_524 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_502 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_525 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_503 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_526 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_504 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_527 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_505 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_528 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_506 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_529 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_507 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_530 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_508 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_531 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_509 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_532 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_510 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_533 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_511 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire  _GEN_535 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_next_config_id : _GEN_1; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [3:0] _GEN_536 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_next_processor_id : _GEN_2; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_556 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_0 : _GEN_22; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_557 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_1 : _GEN_23; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_558 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_2 : _GEN_24; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_559 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_3 : _GEN_25; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_560 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_4 : _GEN_26; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_561 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_5 : _GEN_27; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_562 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_6 : _GEN_28; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_563 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_7 : _GEN_29; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_564 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_8 : _GEN_30; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_565 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_9 : _GEN_31; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_566 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_10 : _GEN_32; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_567 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_11 : _GEN_33; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_568 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_12 : _GEN_34; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_569 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_13 : _GEN_35; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_570 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_14 : _GEN_36; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_571 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_15 : _GEN_37; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_572 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_16 : _GEN_38; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_573 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_17 : _GEN_39; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_574 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_18 : _GEN_40; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_575 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_19 : _GEN_41; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_576 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_20 : _GEN_42; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_577 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_21 : _GEN_43; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_578 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_22 : _GEN_44; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_579 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_23 : _GEN_45; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_580 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_24 : _GEN_46; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_581 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_25 : _GEN_47; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_582 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_26 : _GEN_48; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_583 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_27 : _GEN_49; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_584 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_28 : _GEN_50; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_585 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_29 : _GEN_51; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_586 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_30 : _GEN_52; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_587 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_31 : _GEN_53; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_588 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_32 : _GEN_54; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_589 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_33 : _GEN_55; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_590 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_34 : _GEN_56; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_591 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_35 : _GEN_57; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_592 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_36 : _GEN_58; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_593 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_37 : _GEN_59; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_594 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_38 : _GEN_60; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_595 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_39 : _GEN_61; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_596 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_40 : _GEN_62; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_597 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_41 : _GEN_63; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_598 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_42 : _GEN_64; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_599 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_43 : _GEN_65; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_600 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_44 : _GEN_66; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_601 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_45 : _GEN_67; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_602 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_46 : _GEN_68; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_603 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_47 : _GEN_69; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_604 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_48 : _GEN_70; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_605 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_49 : _GEN_71; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_606 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_50 : _GEN_72; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_607 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_51 : _GEN_73; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_608 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_52 : _GEN_74; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_609 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_53 : _GEN_75; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_610 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_54 : _GEN_76; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_611 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_55 : _GEN_77; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_612 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_56 : _GEN_78; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_613 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_57 : _GEN_79; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_614 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_58 : _GEN_80; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_615 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_59 : _GEN_81; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_616 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_60 : _GEN_82; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_617 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_61 : _GEN_83; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_618 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_62 : _GEN_84; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_619 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_63 : _GEN_85; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_620 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_64 : _GEN_86; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_621 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_65 : _GEN_87; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_622 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_66 : _GEN_88; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_623 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_67 : _GEN_89; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_624 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_68 : _GEN_90; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_625 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_69 : _GEN_91; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_626 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_70 : _GEN_92; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_627 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_71 : _GEN_93; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_628 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_72 : _GEN_94; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_629 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_73 : _GEN_95; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_630 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_74 : _GEN_96; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_631 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_75 : _GEN_97; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_632 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_76 : _GEN_98; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_633 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_77 : _GEN_99; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_634 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_78 : _GEN_100; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_635 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_79 : _GEN_101; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_636 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_80 : _GEN_102; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_637 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_81 : _GEN_103; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_638 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_82 : _GEN_104; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_639 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_83 : _GEN_105; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_640 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_84 : _GEN_106; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_641 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_85 : _GEN_107; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_642 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_86 : _GEN_108; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_643 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_87 : _GEN_109; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_644 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_88 : _GEN_110; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_645 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_89 : _GEN_111; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_646 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_90 : _GEN_112; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_647 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_91 : _GEN_113; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_648 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_92 : _GEN_114; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_649 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_93 : _GEN_115; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_650 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_94 : _GEN_116; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_651 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_95 : _GEN_117; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_652 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_96 : _GEN_118; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_653 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_97 : _GEN_119; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_654 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_98 : _GEN_120; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_655 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_99 : _GEN_121; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_656 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_100 : _GEN_122; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_657 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_101 : _GEN_123; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_658 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_102 : _GEN_124; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_659 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_103 : _GEN_125; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_660 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_104 : _GEN_126; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_661 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_105 : _GEN_127; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_662 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_106 : _GEN_128; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_663 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_107 : _GEN_129; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_664 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_108 : _GEN_130; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_665 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_109 : _GEN_131; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_666 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_110 : _GEN_132; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_667 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_111 : _GEN_133; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_668 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_112 : _GEN_134; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_669 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_113 : _GEN_135; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_670 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_114 : _GEN_136; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_671 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_115 : _GEN_137; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_672 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_116 : _GEN_138; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_673 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_117 : _GEN_139; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_674 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_118 : _GEN_140; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_675 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_119 : _GEN_141; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_676 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_120 : _GEN_142; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_677 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_121 : _GEN_143; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_678 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_122 : _GEN_144; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_679 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_123 : _GEN_145; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_680 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_124 : _GEN_146; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_681 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_125 : _GEN_147; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_682 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_126 : _GEN_148; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_683 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_127 : _GEN_149; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_684 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_128 : _GEN_150; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_685 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_129 : _GEN_151; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_686 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_130 : _GEN_152; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_687 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_131 : _GEN_153; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_688 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_132 : _GEN_154; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_689 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_133 : _GEN_155; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_690 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_134 : _GEN_156; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_691 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_135 : _GEN_157; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_692 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_136 : _GEN_158; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_693 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_137 : _GEN_159; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_694 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_138 : _GEN_160; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_695 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_139 : _GEN_161; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_696 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_140 : _GEN_162; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_697 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_141 : _GEN_163; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_698 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_142 : _GEN_164; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_699 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_143 : _GEN_165; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_700 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_144 : _GEN_166; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_701 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_145 : _GEN_167; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_702 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_146 : _GEN_168; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_703 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_147 : _GEN_169; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_704 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_148 : _GEN_170; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_705 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_149 : _GEN_171; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_706 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_150 : _GEN_172; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_707 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_151 : _GEN_173; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_708 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_152 : _GEN_174; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_709 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_153 : _GEN_175; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_710 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_154 : _GEN_176; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_711 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_155 : _GEN_177; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_712 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_156 : _GEN_178; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_713 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_157 : _GEN_179; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_714 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_158 : _GEN_180; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_715 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_159 : _GEN_181; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_716 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_160 : _GEN_182; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_717 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_161 : _GEN_183; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_718 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_162 : _GEN_184; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_719 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_163 : _GEN_185; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_720 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_164 : _GEN_186; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_721 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_165 : _GEN_187; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_722 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_166 : _GEN_188; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_723 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_167 : _GEN_189; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_724 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_168 : _GEN_190; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_725 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_169 : _GEN_191; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_726 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_170 : _GEN_192; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_727 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_171 : _GEN_193; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_728 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_172 : _GEN_194; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_729 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_173 : _GEN_195; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_730 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_174 : _GEN_196; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_731 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_175 : _GEN_197; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_732 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_176 : _GEN_198; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_733 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_177 : _GEN_199; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_734 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_178 : _GEN_200; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_735 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_179 : _GEN_201; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_736 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_180 : _GEN_202; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_737 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_181 : _GEN_203; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_738 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_182 : _GEN_204; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_739 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_183 : _GEN_205; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_740 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_184 : _GEN_206; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_741 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_185 : _GEN_207; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_742 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_186 : _GEN_208; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_743 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_187 : _GEN_209; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_744 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_188 : _GEN_210; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_745 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_189 : _GEN_211; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_746 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_190 : _GEN_212; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_747 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_191 : _GEN_213; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_748 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_192 : _GEN_214; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_749 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_193 : _GEN_215; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_750 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_194 : _GEN_216; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_751 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_195 : _GEN_217; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_752 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_196 : _GEN_218; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_753 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_197 : _GEN_219; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_754 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_198 : _GEN_220; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_755 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_199 : _GEN_221; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_756 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_200 : _GEN_222; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_757 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_201 : _GEN_223; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_758 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_202 : _GEN_224; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_759 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_203 : _GEN_225; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_760 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_204 : _GEN_226; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_761 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_205 : _GEN_227; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_762 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_206 : _GEN_228; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_763 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_207 : _GEN_229; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_764 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_208 : _GEN_230; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_765 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_209 : _GEN_231; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_766 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_210 : _GEN_232; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_767 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_211 : _GEN_233; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_768 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_212 : _GEN_234; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_769 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_213 : _GEN_235; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_770 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_214 : _GEN_236; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_771 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_215 : _GEN_237; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_772 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_216 : _GEN_238; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_773 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_217 : _GEN_239; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_774 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_218 : _GEN_240; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_775 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_219 : _GEN_241; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_776 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_220 : _GEN_242; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_777 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_221 : _GEN_243; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_778 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_222 : _GEN_244; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_779 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_223 : _GEN_245; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_780 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_224 : _GEN_246; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_781 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_225 : _GEN_247; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_782 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_226 : _GEN_248; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_783 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_227 : _GEN_249; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_784 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_228 : _GEN_250; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_785 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_229 : _GEN_251; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_786 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_230 : _GEN_252; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_787 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_231 : _GEN_253; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_788 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_232 : _GEN_254; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_789 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_233 : _GEN_255; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_790 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_234 : _GEN_256; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_791 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_235 : _GEN_257; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_792 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_236 : _GEN_258; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_793 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_237 : _GEN_259; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_794 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_238 : _GEN_260; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_795 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_239 : _GEN_261; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_796 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_240 : _GEN_262; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_797 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_241 : _GEN_263; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_798 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_242 : _GEN_264; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_799 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_243 : _GEN_265; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_800 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_244 : _GEN_266; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_801 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_245 : _GEN_267; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_802 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_246 : _GEN_268; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_803 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_247 : _GEN_269; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_804 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_248 : _GEN_270; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_805 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_249 : _GEN_271; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_806 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_250 : _GEN_272; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_807 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_251 : _GEN_273; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_808 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_252 : _GEN_274; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_809 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_253 : _GEN_275; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_810 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_254 : _GEN_276; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_811 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_255 : _GEN_277; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_812 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_256 : _GEN_278; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_813 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_257 : _GEN_279; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_814 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_258 : _GEN_280; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_815 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_259 : _GEN_281; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_816 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_260 : _GEN_282; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_817 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_261 : _GEN_283; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_818 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_262 : _GEN_284; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_819 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_263 : _GEN_285; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_820 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_264 : _GEN_286; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_821 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_265 : _GEN_287; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_822 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_266 : _GEN_288; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_823 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_267 : _GEN_289; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_824 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_268 : _GEN_290; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_825 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_269 : _GEN_291; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_826 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_270 : _GEN_292; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_827 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_271 : _GEN_293; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_828 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_272 : _GEN_294; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_829 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_273 : _GEN_295; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_830 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_274 : _GEN_296; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_831 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_275 : _GEN_297; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_832 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_276 : _GEN_298; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_833 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_277 : _GEN_299; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_834 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_278 : _GEN_300; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_835 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_279 : _GEN_301; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_836 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_280 : _GEN_302; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_837 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_281 : _GEN_303; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_838 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_282 : _GEN_304; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_839 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_283 : _GEN_305; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_840 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_284 : _GEN_306; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_841 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_285 : _GEN_307; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_842 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_286 : _GEN_308; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_843 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_287 : _GEN_309; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_844 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_288 : _GEN_310; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_845 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_289 : _GEN_311; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_846 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_290 : _GEN_312; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_847 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_291 : _GEN_313; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_848 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_292 : _GEN_314; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_849 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_293 : _GEN_315; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_850 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_294 : _GEN_316; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_851 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_295 : _GEN_317; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_852 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_296 : _GEN_318; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_853 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_297 : _GEN_319; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_854 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_298 : _GEN_320; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_855 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_299 : _GEN_321; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_856 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_300 : _GEN_322; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_857 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_301 : _GEN_323; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_858 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_302 : _GEN_324; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_859 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_303 : _GEN_325; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_860 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_304 : _GEN_326; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_861 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_305 : _GEN_327; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_862 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_306 : _GEN_328; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_863 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_307 : _GEN_329; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_864 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_308 : _GEN_330; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_865 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_309 : _GEN_331; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_866 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_310 : _GEN_332; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_867 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_311 : _GEN_333; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_868 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_312 : _GEN_334; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_869 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_313 : _GEN_335; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_870 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_314 : _GEN_336; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_871 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_315 : _GEN_337; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_872 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_316 : _GEN_338; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_873 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_317 : _GEN_339; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_874 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_318 : _GEN_340; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_875 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_319 : _GEN_341; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_876 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_320 : _GEN_342; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_877 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_321 : _GEN_343; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_878 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_322 : _GEN_344; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_879 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_323 : _GEN_345; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_880 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_324 : _GEN_346; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_881 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_325 : _GEN_347; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_882 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_326 : _GEN_348; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_883 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_327 : _GEN_349; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_884 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_328 : _GEN_350; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_885 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_329 : _GEN_351; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_886 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_330 : _GEN_352; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_887 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_331 : _GEN_353; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_888 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_332 : _GEN_354; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_889 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_333 : _GEN_355; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_890 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_334 : _GEN_356; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_891 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_335 : _GEN_357; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_892 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_336 : _GEN_358; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_893 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_337 : _GEN_359; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_894 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_338 : _GEN_360; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_895 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_339 : _GEN_361; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_896 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_340 : _GEN_362; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_897 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_341 : _GEN_363; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_898 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_342 : _GEN_364; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_899 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_343 : _GEN_365; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_900 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_344 : _GEN_366; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_901 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_345 : _GEN_367; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_902 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_346 : _GEN_368; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_903 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_347 : _GEN_369; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_904 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_348 : _GEN_370; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_905 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_349 : _GEN_371; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_906 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_350 : _GEN_372; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_907 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_351 : _GEN_373; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_908 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_352 : _GEN_374; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_909 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_353 : _GEN_375; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_910 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_354 : _GEN_376; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_911 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_355 : _GEN_377; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_912 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_356 : _GEN_378; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_913 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_357 : _GEN_379; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_914 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_358 : _GEN_380; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_915 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_359 : _GEN_381; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_916 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_360 : _GEN_382; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_917 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_361 : _GEN_383; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_918 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_362 : _GEN_384; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_919 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_363 : _GEN_385; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_920 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_364 : _GEN_386; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_921 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_365 : _GEN_387; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_922 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_366 : _GEN_388; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_923 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_367 : _GEN_389; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_924 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_368 : _GEN_390; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_925 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_369 : _GEN_391; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_926 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_370 : _GEN_392; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_927 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_371 : _GEN_393; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_928 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_372 : _GEN_394; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_929 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_373 : _GEN_395; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_930 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_374 : _GEN_396; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_931 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_375 : _GEN_397; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_932 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_376 : _GEN_398; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_933 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_377 : _GEN_399; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_934 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_378 : _GEN_400; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_935 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_379 : _GEN_401; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_936 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_380 : _GEN_402; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_937 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_381 : _GEN_403; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_938 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_382 : _GEN_404; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_939 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_383 : _GEN_405; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_940 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_384 : _GEN_406; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_941 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_385 : _GEN_407; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_942 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_386 : _GEN_408; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_943 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_387 : _GEN_409; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_944 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_388 : _GEN_410; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_945 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_389 : _GEN_411; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_946 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_390 : _GEN_412; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_947 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_391 : _GEN_413; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_948 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_392 : _GEN_414; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_949 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_393 : _GEN_415; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_950 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_394 : _GEN_416; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_951 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_395 : _GEN_417; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_952 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_396 : _GEN_418; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_953 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_397 : _GEN_419; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_954 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_398 : _GEN_420; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_955 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_399 : _GEN_421; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_956 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_400 : _GEN_422; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_957 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_401 : _GEN_423; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_958 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_402 : _GEN_424; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_959 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_403 : _GEN_425; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_960 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_404 : _GEN_426; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_961 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_405 : _GEN_427; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_962 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_406 : _GEN_428; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_963 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_407 : _GEN_429; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_964 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_408 : _GEN_430; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_965 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_409 : _GEN_431; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_966 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_410 : _GEN_432; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_967 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_411 : _GEN_433; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_968 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_412 : _GEN_434; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_969 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_413 : _GEN_435; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_970 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_414 : _GEN_436; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_971 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_415 : _GEN_437; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_972 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_416 : _GEN_438; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_973 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_417 : _GEN_439; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_974 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_418 : _GEN_440; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_975 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_419 : _GEN_441; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_976 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_420 : _GEN_442; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_977 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_421 : _GEN_443; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_978 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_422 : _GEN_444; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_979 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_423 : _GEN_445; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_980 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_424 : _GEN_446; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_981 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_425 : _GEN_447; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_982 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_426 : _GEN_448; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_983 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_427 : _GEN_449; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_984 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_428 : _GEN_450; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_985 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_429 : _GEN_451; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_986 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_430 : _GEN_452; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_987 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_431 : _GEN_453; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_988 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_432 : _GEN_454; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_989 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_433 : _GEN_455; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_990 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_434 : _GEN_456; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_991 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_435 : _GEN_457; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_992 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_436 : _GEN_458; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_993 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_437 : _GEN_459; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_994 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_438 : _GEN_460; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_995 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_439 : _GEN_461; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_996 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_440 : _GEN_462; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_997 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_441 : _GEN_463; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_998 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_442 : _GEN_464; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_999 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_443 : _GEN_465; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1000 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_444 : _GEN_466; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1001 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_445 : _GEN_467; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1002 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_446 : _GEN_468; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1003 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_447 : _GEN_469; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1004 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_448 : _GEN_470; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1005 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_449 : _GEN_471; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1006 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_450 : _GEN_472; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1007 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_451 : _GEN_473; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1008 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_452 : _GEN_474; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1009 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_453 : _GEN_475; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1010 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_454 : _GEN_476; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1011 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_455 : _GEN_477; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1012 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_456 : _GEN_478; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1013 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_457 : _GEN_479; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1014 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_458 : _GEN_480; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1015 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_459 : _GEN_481; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1016 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_460 : _GEN_482; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1017 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_461 : _GEN_483; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1018 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_462 : _GEN_484; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1019 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_463 : _GEN_485; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1020 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_464 : _GEN_486; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1021 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_465 : _GEN_487; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1022 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_466 : _GEN_488; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1023 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_467 : _GEN_489; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1024 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_468 : _GEN_490; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1025 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_469 : _GEN_491; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1026 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_470 : _GEN_492; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1027 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_471 : _GEN_493; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1028 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_472 : _GEN_494; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1029 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_473 : _GEN_495; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1030 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_474 : _GEN_496; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1031 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_475 : _GEN_497; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1032 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_476 : _GEN_498; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1033 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_477 : _GEN_499; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1034 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_478 : _GEN_500; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1035 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_479 : _GEN_501; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1036 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_480 : _GEN_502; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1037 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_481 : _GEN_503; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1038 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_482 : _GEN_504; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1039 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_483 : _GEN_505; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1040 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_484 : _GEN_506; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1041 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_485 : _GEN_507; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1042 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_486 : _GEN_508; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1043 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_487 : _GEN_509; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1044 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_488 : _GEN_510; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1045 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_489 : _GEN_511; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1046 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_490 : _GEN_512; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1047 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_491 : _GEN_513; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1048 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_492 : _GEN_514; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1049 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_493 : _GEN_515; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1050 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_494 : _GEN_516; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1051 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_495 : _GEN_517; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1052 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_496 : _GEN_518; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1053 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_497 : _GEN_519; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1054 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_498 : _GEN_520; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1055 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_499 : _GEN_521; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1056 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_500 : _GEN_522; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1057 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_501 : _GEN_523; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1058 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_502 : _GEN_524; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1059 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_503 : _GEN_525; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1060 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_504 : _GEN_526; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1061 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_505 : _GEN_527; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1062 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_506 : _GEN_528; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1063 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_507 : _GEN_529; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1064 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_508 : _GEN_530; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1065 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_509 : _GEN_531; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1066 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_510 : _GEN_532; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1067 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_511 : _GEN_533; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire  _GEN_1069 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_next_config_id : _GEN_535; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [3:0] _GEN_1070 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_next_processor_id : _GEN_536; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1090 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_0 : _GEN_556; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1091 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_1 : _GEN_557; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1092 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_2 : _GEN_558; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1093 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_3 : _GEN_559; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1094 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_4 : _GEN_560; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1095 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_5 : _GEN_561; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1096 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_6 : _GEN_562; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1097 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_7 : _GEN_563; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1098 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_8 : _GEN_564; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1099 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_9 : _GEN_565; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1100 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_10 : _GEN_566; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1101 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_11 : _GEN_567; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1102 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_12 : _GEN_568; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1103 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_13 : _GEN_569; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1104 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_14 : _GEN_570; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1105 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_15 : _GEN_571; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1106 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_16 : _GEN_572; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1107 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_17 : _GEN_573; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1108 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_18 : _GEN_574; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1109 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_19 : _GEN_575; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1110 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_20 : _GEN_576; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1111 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_21 : _GEN_577; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1112 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_22 : _GEN_578; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1113 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_23 : _GEN_579; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1114 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_24 : _GEN_580; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1115 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_25 : _GEN_581; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1116 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_26 : _GEN_582; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1117 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_27 : _GEN_583; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1118 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_28 : _GEN_584; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1119 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_29 : _GEN_585; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1120 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_30 : _GEN_586; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1121 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_31 : _GEN_587; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1122 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_32 : _GEN_588; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1123 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_33 : _GEN_589; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1124 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_34 : _GEN_590; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1125 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_35 : _GEN_591; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1126 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_36 : _GEN_592; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1127 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_37 : _GEN_593; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1128 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_38 : _GEN_594; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1129 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_39 : _GEN_595; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1130 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_40 : _GEN_596; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1131 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_41 : _GEN_597; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1132 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_42 : _GEN_598; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1133 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_43 : _GEN_599; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1134 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_44 : _GEN_600; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1135 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_45 : _GEN_601; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1136 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_46 : _GEN_602; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1137 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_47 : _GEN_603; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1138 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_48 : _GEN_604; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1139 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_49 : _GEN_605; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1140 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_50 : _GEN_606; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1141 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_51 : _GEN_607; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1142 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_52 : _GEN_608; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1143 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_53 : _GEN_609; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1144 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_54 : _GEN_610; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1145 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_55 : _GEN_611; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1146 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_56 : _GEN_612; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1147 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_57 : _GEN_613; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1148 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_58 : _GEN_614; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1149 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_59 : _GEN_615; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1150 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_60 : _GEN_616; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1151 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_61 : _GEN_617; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1152 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_62 : _GEN_618; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1153 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_63 : _GEN_619; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1154 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_64 : _GEN_620; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1155 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_65 : _GEN_621; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1156 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_66 : _GEN_622; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1157 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_67 : _GEN_623; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1158 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_68 : _GEN_624; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1159 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_69 : _GEN_625; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1160 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_70 : _GEN_626; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1161 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_71 : _GEN_627; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1162 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_72 : _GEN_628; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1163 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_73 : _GEN_629; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1164 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_74 : _GEN_630; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1165 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_75 : _GEN_631; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1166 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_76 : _GEN_632; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1167 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_77 : _GEN_633; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1168 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_78 : _GEN_634; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1169 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_79 : _GEN_635; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1170 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_80 : _GEN_636; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1171 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_81 : _GEN_637; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1172 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_82 : _GEN_638; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1173 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_83 : _GEN_639; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1174 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_84 : _GEN_640; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1175 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_85 : _GEN_641; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1176 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_86 : _GEN_642; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1177 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_87 : _GEN_643; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1178 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_88 : _GEN_644; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1179 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_89 : _GEN_645; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1180 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_90 : _GEN_646; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1181 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_91 : _GEN_647; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1182 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_92 : _GEN_648; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1183 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_93 : _GEN_649; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1184 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_94 : _GEN_650; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1185 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_95 : _GEN_651; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1186 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_96 : _GEN_652; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1187 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_97 : _GEN_653; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1188 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_98 : _GEN_654; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1189 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_99 : _GEN_655; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1190 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_100 : _GEN_656; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1191 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_101 : _GEN_657; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1192 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_102 : _GEN_658; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1193 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_103 : _GEN_659; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1194 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_104 : _GEN_660; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1195 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_105 : _GEN_661; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1196 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_106 : _GEN_662; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1197 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_107 : _GEN_663; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1198 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_108 : _GEN_664; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1199 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_109 : _GEN_665; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1200 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_110 : _GEN_666; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1201 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_111 : _GEN_667; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1202 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_112 : _GEN_668; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1203 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_113 : _GEN_669; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1204 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_114 : _GEN_670; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1205 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_115 : _GEN_671; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1206 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_116 : _GEN_672; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1207 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_117 : _GEN_673; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1208 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_118 : _GEN_674; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1209 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_119 : _GEN_675; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1210 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_120 : _GEN_676; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1211 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_121 : _GEN_677; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1212 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_122 : _GEN_678; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1213 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_123 : _GEN_679; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1214 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_124 : _GEN_680; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1215 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_125 : _GEN_681; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1216 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_126 : _GEN_682; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1217 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_127 : _GEN_683; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1218 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_128 : _GEN_684; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1219 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_129 : _GEN_685; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1220 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_130 : _GEN_686; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1221 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_131 : _GEN_687; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1222 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_132 : _GEN_688; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1223 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_133 : _GEN_689; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1224 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_134 : _GEN_690; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1225 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_135 : _GEN_691; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1226 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_136 : _GEN_692; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1227 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_137 : _GEN_693; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1228 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_138 : _GEN_694; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1229 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_139 : _GEN_695; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1230 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_140 : _GEN_696; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1231 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_141 : _GEN_697; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1232 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_142 : _GEN_698; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1233 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_143 : _GEN_699; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1234 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_144 : _GEN_700; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1235 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_145 : _GEN_701; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1236 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_146 : _GEN_702; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1237 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_147 : _GEN_703; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1238 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_148 : _GEN_704; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1239 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_149 : _GEN_705; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1240 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_150 : _GEN_706; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1241 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_151 : _GEN_707; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1242 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_152 : _GEN_708; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1243 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_153 : _GEN_709; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1244 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_154 : _GEN_710; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1245 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_155 : _GEN_711; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1246 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_156 : _GEN_712; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1247 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_157 : _GEN_713; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1248 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_158 : _GEN_714; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1249 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_159 : _GEN_715; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1250 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_160 : _GEN_716; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1251 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_161 : _GEN_717; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1252 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_162 : _GEN_718; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1253 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_163 : _GEN_719; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1254 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_164 : _GEN_720; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1255 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_165 : _GEN_721; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1256 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_166 : _GEN_722; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1257 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_167 : _GEN_723; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1258 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_168 : _GEN_724; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1259 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_169 : _GEN_725; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1260 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_170 : _GEN_726; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1261 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_171 : _GEN_727; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1262 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_172 : _GEN_728; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1263 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_173 : _GEN_729; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1264 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_174 : _GEN_730; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1265 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_175 : _GEN_731; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1266 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_176 : _GEN_732; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1267 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_177 : _GEN_733; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1268 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_178 : _GEN_734; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1269 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_179 : _GEN_735; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1270 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_180 : _GEN_736; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1271 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_181 : _GEN_737; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1272 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_182 : _GEN_738; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1273 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_183 : _GEN_739; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1274 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_184 : _GEN_740; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1275 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_185 : _GEN_741; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1276 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_186 : _GEN_742; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1277 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_187 : _GEN_743; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1278 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_188 : _GEN_744; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1279 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_189 : _GEN_745; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1280 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_190 : _GEN_746; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1281 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_191 : _GEN_747; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1282 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_192 : _GEN_748; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1283 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_193 : _GEN_749; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1284 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_194 : _GEN_750; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1285 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_195 : _GEN_751; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1286 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_196 : _GEN_752; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1287 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_197 : _GEN_753; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1288 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_198 : _GEN_754; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1289 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_199 : _GEN_755; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1290 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_200 : _GEN_756; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1291 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_201 : _GEN_757; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1292 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_202 : _GEN_758; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1293 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_203 : _GEN_759; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1294 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_204 : _GEN_760; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1295 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_205 : _GEN_761; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1296 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_206 : _GEN_762; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1297 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_207 : _GEN_763; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1298 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_208 : _GEN_764; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1299 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_209 : _GEN_765; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1300 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_210 : _GEN_766; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1301 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_211 : _GEN_767; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1302 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_212 : _GEN_768; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1303 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_213 : _GEN_769; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1304 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_214 : _GEN_770; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1305 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_215 : _GEN_771; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1306 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_216 : _GEN_772; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1307 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_217 : _GEN_773; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1308 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_218 : _GEN_774; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1309 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_219 : _GEN_775; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1310 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_220 : _GEN_776; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1311 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_221 : _GEN_777; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1312 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_222 : _GEN_778; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1313 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_223 : _GEN_779; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1314 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_224 : _GEN_780; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1315 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_225 : _GEN_781; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1316 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_226 : _GEN_782; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1317 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_227 : _GEN_783; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1318 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_228 : _GEN_784; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1319 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_229 : _GEN_785; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1320 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_230 : _GEN_786; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1321 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_231 : _GEN_787; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1322 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_232 : _GEN_788; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1323 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_233 : _GEN_789; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1324 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_234 : _GEN_790; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1325 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_235 : _GEN_791; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1326 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_236 : _GEN_792; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1327 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_237 : _GEN_793; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1328 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_238 : _GEN_794; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1329 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_239 : _GEN_795; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1330 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_240 : _GEN_796; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1331 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_241 : _GEN_797; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1332 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_242 : _GEN_798; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1333 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_243 : _GEN_799; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1334 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_244 : _GEN_800; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1335 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_245 : _GEN_801; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1336 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_246 : _GEN_802; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1337 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_247 : _GEN_803; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1338 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_248 : _GEN_804; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1339 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_249 : _GEN_805; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1340 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_250 : _GEN_806; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1341 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_251 : _GEN_807; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1342 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_252 : _GEN_808; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1343 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_253 : _GEN_809; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1344 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_254 : _GEN_810; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1345 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_255 : _GEN_811; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1346 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_256 : _GEN_812; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1347 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_257 : _GEN_813; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1348 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_258 : _GEN_814; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1349 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_259 : _GEN_815; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1350 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_260 : _GEN_816; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1351 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_261 : _GEN_817; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1352 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_262 : _GEN_818; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1353 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_263 : _GEN_819; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1354 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_264 : _GEN_820; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1355 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_265 : _GEN_821; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1356 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_266 : _GEN_822; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1357 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_267 : _GEN_823; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1358 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_268 : _GEN_824; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1359 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_269 : _GEN_825; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1360 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_270 : _GEN_826; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1361 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_271 : _GEN_827; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1362 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_272 : _GEN_828; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1363 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_273 : _GEN_829; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1364 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_274 : _GEN_830; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1365 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_275 : _GEN_831; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1366 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_276 : _GEN_832; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1367 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_277 : _GEN_833; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1368 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_278 : _GEN_834; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1369 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_279 : _GEN_835; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1370 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_280 : _GEN_836; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1371 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_281 : _GEN_837; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1372 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_282 : _GEN_838; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1373 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_283 : _GEN_839; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1374 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_284 : _GEN_840; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1375 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_285 : _GEN_841; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1376 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_286 : _GEN_842; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1377 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_287 : _GEN_843; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1378 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_288 : _GEN_844; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1379 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_289 : _GEN_845; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1380 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_290 : _GEN_846; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1381 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_291 : _GEN_847; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1382 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_292 : _GEN_848; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1383 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_293 : _GEN_849; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1384 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_294 : _GEN_850; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1385 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_295 : _GEN_851; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1386 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_296 : _GEN_852; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1387 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_297 : _GEN_853; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1388 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_298 : _GEN_854; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1389 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_299 : _GEN_855; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1390 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_300 : _GEN_856; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1391 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_301 : _GEN_857; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1392 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_302 : _GEN_858; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1393 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_303 : _GEN_859; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1394 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_304 : _GEN_860; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1395 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_305 : _GEN_861; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1396 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_306 : _GEN_862; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1397 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_307 : _GEN_863; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1398 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_308 : _GEN_864; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1399 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_309 : _GEN_865; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1400 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_310 : _GEN_866; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1401 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_311 : _GEN_867; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1402 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_312 : _GEN_868; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1403 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_313 : _GEN_869; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1404 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_314 : _GEN_870; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1405 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_315 : _GEN_871; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1406 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_316 : _GEN_872; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1407 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_317 : _GEN_873; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1408 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_318 : _GEN_874; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1409 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_319 : _GEN_875; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1410 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_320 : _GEN_876; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1411 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_321 : _GEN_877; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1412 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_322 : _GEN_878; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1413 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_323 : _GEN_879; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1414 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_324 : _GEN_880; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1415 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_325 : _GEN_881; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1416 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_326 : _GEN_882; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1417 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_327 : _GEN_883; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1418 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_328 : _GEN_884; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1419 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_329 : _GEN_885; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1420 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_330 : _GEN_886; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1421 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_331 : _GEN_887; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1422 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_332 : _GEN_888; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1423 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_333 : _GEN_889; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1424 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_334 : _GEN_890; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1425 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_335 : _GEN_891; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1426 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_336 : _GEN_892; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1427 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_337 : _GEN_893; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1428 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_338 : _GEN_894; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1429 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_339 : _GEN_895; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1430 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_340 : _GEN_896; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1431 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_341 : _GEN_897; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1432 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_342 : _GEN_898; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1433 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_343 : _GEN_899; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1434 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_344 : _GEN_900; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1435 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_345 : _GEN_901; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1436 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_346 : _GEN_902; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1437 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_347 : _GEN_903; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1438 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_348 : _GEN_904; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1439 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_349 : _GEN_905; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1440 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_350 : _GEN_906; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1441 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_351 : _GEN_907; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1442 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_352 : _GEN_908; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1443 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_353 : _GEN_909; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1444 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_354 : _GEN_910; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1445 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_355 : _GEN_911; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1446 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_356 : _GEN_912; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1447 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_357 : _GEN_913; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1448 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_358 : _GEN_914; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1449 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_359 : _GEN_915; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1450 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_360 : _GEN_916; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1451 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_361 : _GEN_917; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1452 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_362 : _GEN_918; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1453 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_363 : _GEN_919; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1454 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_364 : _GEN_920; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1455 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_365 : _GEN_921; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1456 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_366 : _GEN_922; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1457 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_367 : _GEN_923; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1458 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_368 : _GEN_924; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1459 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_369 : _GEN_925; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1460 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_370 : _GEN_926; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1461 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_371 : _GEN_927; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1462 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_372 : _GEN_928; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1463 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_373 : _GEN_929; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1464 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_374 : _GEN_930; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1465 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_375 : _GEN_931; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1466 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_376 : _GEN_932; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1467 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_377 : _GEN_933; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1468 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_378 : _GEN_934; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1469 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_379 : _GEN_935; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1470 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_380 : _GEN_936; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1471 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_381 : _GEN_937; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1472 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_382 : _GEN_938; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1473 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_383 : _GEN_939; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1474 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_384 : _GEN_940; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1475 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_385 : _GEN_941; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1476 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_386 : _GEN_942; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1477 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_387 : _GEN_943; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1478 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_388 : _GEN_944; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1479 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_389 : _GEN_945; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1480 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_390 : _GEN_946; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1481 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_391 : _GEN_947; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1482 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_392 : _GEN_948; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1483 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_393 : _GEN_949; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1484 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_394 : _GEN_950; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1485 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_395 : _GEN_951; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1486 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_396 : _GEN_952; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1487 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_397 : _GEN_953; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1488 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_398 : _GEN_954; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1489 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_399 : _GEN_955; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1490 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_400 : _GEN_956; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1491 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_401 : _GEN_957; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1492 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_402 : _GEN_958; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1493 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_403 : _GEN_959; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1494 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_404 : _GEN_960; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1495 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_405 : _GEN_961; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1496 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_406 : _GEN_962; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1497 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_407 : _GEN_963; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1498 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_408 : _GEN_964; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1499 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_409 : _GEN_965; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1500 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_410 : _GEN_966; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1501 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_411 : _GEN_967; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1502 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_412 : _GEN_968; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1503 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_413 : _GEN_969; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1504 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_414 : _GEN_970; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1505 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_415 : _GEN_971; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1506 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_416 : _GEN_972; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1507 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_417 : _GEN_973; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1508 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_418 : _GEN_974; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1509 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_419 : _GEN_975; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1510 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_420 : _GEN_976; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1511 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_421 : _GEN_977; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1512 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_422 : _GEN_978; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1513 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_423 : _GEN_979; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1514 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_424 : _GEN_980; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1515 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_425 : _GEN_981; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1516 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_426 : _GEN_982; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1517 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_427 : _GEN_983; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1518 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_428 : _GEN_984; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1519 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_429 : _GEN_985; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1520 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_430 : _GEN_986; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1521 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_431 : _GEN_987; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1522 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_432 : _GEN_988; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1523 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_433 : _GEN_989; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1524 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_434 : _GEN_990; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1525 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_435 : _GEN_991; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1526 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_436 : _GEN_992; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1527 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_437 : _GEN_993; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1528 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_438 : _GEN_994; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1529 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_439 : _GEN_995; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1530 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_440 : _GEN_996; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1531 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_441 : _GEN_997; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1532 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_442 : _GEN_998; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1533 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_443 : _GEN_999; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1534 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_444 : _GEN_1000; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1535 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_445 : _GEN_1001; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1536 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_446 : _GEN_1002; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1537 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_447 : _GEN_1003; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1538 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_448 : _GEN_1004; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1539 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_449 : _GEN_1005; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1540 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_450 : _GEN_1006; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1541 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_451 : _GEN_1007; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1542 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_452 : _GEN_1008; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1543 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_453 : _GEN_1009; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1544 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_454 : _GEN_1010; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1545 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_455 : _GEN_1011; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1546 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_456 : _GEN_1012; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1547 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_457 : _GEN_1013; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1548 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_458 : _GEN_1014; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1549 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_459 : _GEN_1015; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1550 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_460 : _GEN_1016; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1551 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_461 : _GEN_1017; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1552 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_462 : _GEN_1018; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1553 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_463 : _GEN_1019; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1554 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_464 : _GEN_1020; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1555 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_465 : _GEN_1021; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1556 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_466 : _GEN_1022; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1557 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_467 : _GEN_1023; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1558 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_468 : _GEN_1024; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1559 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_469 : _GEN_1025; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1560 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_470 : _GEN_1026; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1561 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_471 : _GEN_1027; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1562 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_472 : _GEN_1028; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1563 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_473 : _GEN_1029; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1564 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_474 : _GEN_1030; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1565 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_475 : _GEN_1031; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1566 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_476 : _GEN_1032; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1567 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_477 : _GEN_1033; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1568 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_478 : _GEN_1034; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1569 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_479 : _GEN_1035; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1570 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_480 : _GEN_1036; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1571 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_481 : _GEN_1037; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1572 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_482 : _GEN_1038; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1573 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_483 : _GEN_1039; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1574 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_484 : _GEN_1040; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1575 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_485 : _GEN_1041; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1576 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_486 : _GEN_1042; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1577 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_487 : _GEN_1043; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1578 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_488 : _GEN_1044; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1579 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_489 : _GEN_1045; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1580 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_490 : _GEN_1046; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1581 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_491 : _GEN_1047; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1582 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_492 : _GEN_1048; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1583 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_493 : _GEN_1049; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1584 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_494 : _GEN_1050; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1585 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_495 : _GEN_1051; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1586 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_496 : _GEN_1052; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1587 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_497 : _GEN_1053; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1588 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_498 : _GEN_1054; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1589 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_499 : _GEN_1055; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1590 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_500 : _GEN_1056; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1591 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_501 : _GEN_1057; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1592 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_502 : _GEN_1058; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1593 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_503 : _GEN_1059; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1594 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_504 : _GEN_1060; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1595 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_505 : _GEN_1061; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1596 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_506 : _GEN_1062; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1597 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_507 : _GEN_1063; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1598 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_508 : _GEN_1064; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1599 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_509 : _GEN_1065; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1600 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_510 : _GEN_1066; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1601 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_511 : _GEN_1067; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire  _GEN_1603 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_next_config_id : _GEN_1069; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [3:0] _GEN_1604 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_next_processor_id : _GEN_1070; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1624 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_0 : _GEN_1090; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1625 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_1 : _GEN_1091; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1626 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_2 : _GEN_1092; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1627 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_3 : _GEN_1093; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1628 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_4 : _GEN_1094; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1629 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_5 : _GEN_1095; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1630 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_6 : _GEN_1096; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1631 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_7 : _GEN_1097; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1632 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_8 : _GEN_1098; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1633 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_9 : _GEN_1099; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1634 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_10 : _GEN_1100; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1635 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_11 : _GEN_1101; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1636 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_12 : _GEN_1102; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1637 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_13 : _GEN_1103; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1638 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_14 : _GEN_1104; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1639 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_15 : _GEN_1105; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1640 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_16 : _GEN_1106; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1641 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_17 : _GEN_1107; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1642 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_18 : _GEN_1108; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1643 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_19 : _GEN_1109; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1644 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_20 : _GEN_1110; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1645 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_21 : _GEN_1111; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1646 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_22 : _GEN_1112; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1647 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_23 : _GEN_1113; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1648 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_24 : _GEN_1114; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1649 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_25 : _GEN_1115; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1650 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_26 : _GEN_1116; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1651 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_27 : _GEN_1117; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1652 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_28 : _GEN_1118; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1653 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_29 : _GEN_1119; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1654 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_30 : _GEN_1120; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1655 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_31 : _GEN_1121; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1656 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_32 : _GEN_1122; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1657 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_33 : _GEN_1123; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1658 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_34 : _GEN_1124; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1659 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_35 : _GEN_1125; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1660 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_36 : _GEN_1126; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1661 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_37 : _GEN_1127; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1662 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_38 : _GEN_1128; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1663 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_39 : _GEN_1129; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1664 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_40 : _GEN_1130; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1665 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_41 : _GEN_1131; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1666 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_42 : _GEN_1132; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1667 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_43 : _GEN_1133; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1668 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_44 : _GEN_1134; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1669 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_45 : _GEN_1135; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1670 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_46 : _GEN_1136; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1671 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_47 : _GEN_1137; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1672 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_48 : _GEN_1138; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1673 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_49 : _GEN_1139; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1674 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_50 : _GEN_1140; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1675 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_51 : _GEN_1141; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1676 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_52 : _GEN_1142; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1677 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_53 : _GEN_1143; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1678 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_54 : _GEN_1144; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1679 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_55 : _GEN_1145; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1680 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_56 : _GEN_1146; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1681 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_57 : _GEN_1147; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1682 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_58 : _GEN_1148; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1683 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_59 : _GEN_1149; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1684 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_60 : _GEN_1150; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1685 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_61 : _GEN_1151; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1686 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_62 : _GEN_1152; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1687 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_63 : _GEN_1153; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1688 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_64 : _GEN_1154; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1689 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_65 : _GEN_1155; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1690 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_66 : _GEN_1156; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1691 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_67 : _GEN_1157; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1692 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_68 : _GEN_1158; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1693 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_69 : _GEN_1159; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1694 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_70 : _GEN_1160; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1695 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_71 : _GEN_1161; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1696 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_72 : _GEN_1162; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1697 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_73 : _GEN_1163; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1698 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_74 : _GEN_1164; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1699 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_75 : _GEN_1165; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1700 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_76 : _GEN_1166; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1701 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_77 : _GEN_1167; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1702 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_78 : _GEN_1168; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1703 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_79 : _GEN_1169; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1704 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_80 : _GEN_1170; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1705 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_81 : _GEN_1171; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1706 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_82 : _GEN_1172; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1707 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_83 : _GEN_1173; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1708 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_84 : _GEN_1174; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1709 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_85 : _GEN_1175; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1710 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_86 : _GEN_1176; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1711 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_87 : _GEN_1177; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1712 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_88 : _GEN_1178; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1713 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_89 : _GEN_1179; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1714 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_90 : _GEN_1180; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1715 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_91 : _GEN_1181; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1716 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_92 : _GEN_1182; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1717 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_93 : _GEN_1183; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1718 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_94 : _GEN_1184; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1719 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_95 : _GEN_1185; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1720 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_96 : _GEN_1186; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1721 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_97 : _GEN_1187; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1722 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_98 : _GEN_1188; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1723 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_99 : _GEN_1189; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1724 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_100 : _GEN_1190; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1725 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_101 : _GEN_1191; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1726 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_102 : _GEN_1192; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1727 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_103 : _GEN_1193; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1728 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_104 : _GEN_1194; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1729 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_105 : _GEN_1195; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1730 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_106 : _GEN_1196; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1731 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_107 : _GEN_1197; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1732 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_108 : _GEN_1198; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1733 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_109 : _GEN_1199; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1734 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_110 : _GEN_1200; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1735 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_111 : _GEN_1201; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1736 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_112 : _GEN_1202; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1737 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_113 : _GEN_1203; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1738 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_114 : _GEN_1204; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1739 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_115 : _GEN_1205; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1740 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_116 : _GEN_1206; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1741 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_117 : _GEN_1207; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1742 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_118 : _GEN_1208; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1743 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_119 : _GEN_1209; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1744 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_120 : _GEN_1210; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1745 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_121 : _GEN_1211; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1746 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_122 : _GEN_1212; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1747 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_123 : _GEN_1213; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1748 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_124 : _GEN_1214; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1749 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_125 : _GEN_1215; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1750 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_126 : _GEN_1216; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1751 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_127 : _GEN_1217; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1752 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_128 : _GEN_1218; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1753 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_129 : _GEN_1219; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1754 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_130 : _GEN_1220; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1755 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_131 : _GEN_1221; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1756 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_132 : _GEN_1222; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1757 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_133 : _GEN_1223; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1758 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_134 : _GEN_1224; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1759 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_135 : _GEN_1225; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1760 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_136 : _GEN_1226; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1761 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_137 : _GEN_1227; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1762 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_138 : _GEN_1228; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1763 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_139 : _GEN_1229; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1764 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_140 : _GEN_1230; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1765 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_141 : _GEN_1231; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1766 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_142 : _GEN_1232; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1767 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_143 : _GEN_1233; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1768 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_144 : _GEN_1234; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1769 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_145 : _GEN_1235; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1770 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_146 : _GEN_1236; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1771 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_147 : _GEN_1237; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1772 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_148 : _GEN_1238; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1773 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_149 : _GEN_1239; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1774 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_150 : _GEN_1240; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1775 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_151 : _GEN_1241; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1776 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_152 : _GEN_1242; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1777 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_153 : _GEN_1243; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1778 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_154 : _GEN_1244; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1779 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_155 : _GEN_1245; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1780 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_156 : _GEN_1246; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1781 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_157 : _GEN_1247; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1782 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_158 : _GEN_1248; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1783 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_159 : _GEN_1249; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1784 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_160 : _GEN_1250; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1785 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_161 : _GEN_1251; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1786 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_162 : _GEN_1252; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1787 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_163 : _GEN_1253; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1788 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_164 : _GEN_1254; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1789 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_165 : _GEN_1255; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1790 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_166 : _GEN_1256; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1791 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_167 : _GEN_1257; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1792 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_168 : _GEN_1258; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1793 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_169 : _GEN_1259; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1794 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_170 : _GEN_1260; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1795 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_171 : _GEN_1261; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1796 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_172 : _GEN_1262; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1797 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_173 : _GEN_1263; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1798 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_174 : _GEN_1264; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1799 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_175 : _GEN_1265; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1800 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_176 : _GEN_1266; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1801 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_177 : _GEN_1267; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1802 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_178 : _GEN_1268; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1803 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_179 : _GEN_1269; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1804 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_180 : _GEN_1270; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1805 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_181 : _GEN_1271; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1806 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_182 : _GEN_1272; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1807 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_183 : _GEN_1273; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1808 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_184 : _GEN_1274; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1809 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_185 : _GEN_1275; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1810 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_186 : _GEN_1276; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1811 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_187 : _GEN_1277; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1812 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_188 : _GEN_1278; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1813 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_189 : _GEN_1279; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1814 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_190 : _GEN_1280; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1815 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_191 : _GEN_1281; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1816 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_192 : _GEN_1282; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1817 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_193 : _GEN_1283; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1818 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_194 : _GEN_1284; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1819 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_195 : _GEN_1285; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1820 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_196 : _GEN_1286; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1821 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_197 : _GEN_1287; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1822 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_198 : _GEN_1288; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1823 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_199 : _GEN_1289; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1824 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_200 : _GEN_1290; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1825 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_201 : _GEN_1291; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1826 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_202 : _GEN_1292; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1827 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_203 : _GEN_1293; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1828 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_204 : _GEN_1294; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1829 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_205 : _GEN_1295; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1830 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_206 : _GEN_1296; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1831 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_207 : _GEN_1297; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1832 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_208 : _GEN_1298; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1833 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_209 : _GEN_1299; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1834 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_210 : _GEN_1300; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1835 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_211 : _GEN_1301; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1836 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_212 : _GEN_1302; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1837 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_213 : _GEN_1303; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1838 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_214 : _GEN_1304; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1839 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_215 : _GEN_1305; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1840 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_216 : _GEN_1306; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1841 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_217 : _GEN_1307; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1842 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_218 : _GEN_1308; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1843 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_219 : _GEN_1309; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1844 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_220 : _GEN_1310; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1845 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_221 : _GEN_1311; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1846 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_222 : _GEN_1312; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1847 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_223 : _GEN_1313; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1848 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_224 : _GEN_1314; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1849 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_225 : _GEN_1315; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1850 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_226 : _GEN_1316; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1851 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_227 : _GEN_1317; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1852 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_228 : _GEN_1318; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1853 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_229 : _GEN_1319; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1854 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_230 : _GEN_1320; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1855 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_231 : _GEN_1321; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1856 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_232 : _GEN_1322; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1857 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_233 : _GEN_1323; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1858 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_234 : _GEN_1324; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1859 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_235 : _GEN_1325; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1860 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_236 : _GEN_1326; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1861 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_237 : _GEN_1327; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1862 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_238 : _GEN_1328; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1863 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_239 : _GEN_1329; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1864 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_240 : _GEN_1330; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1865 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_241 : _GEN_1331; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1866 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_242 : _GEN_1332; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1867 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_243 : _GEN_1333; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1868 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_244 : _GEN_1334; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1869 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_245 : _GEN_1335; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1870 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_246 : _GEN_1336; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1871 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_247 : _GEN_1337; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1872 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_248 : _GEN_1338; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1873 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_249 : _GEN_1339; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1874 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_250 : _GEN_1340; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1875 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_251 : _GEN_1341; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1876 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_252 : _GEN_1342; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1877 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_253 : _GEN_1343; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1878 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_254 : _GEN_1344; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1879 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_255 : _GEN_1345; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1880 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_256 : _GEN_1346; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1881 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_257 : _GEN_1347; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1882 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_258 : _GEN_1348; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1883 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_259 : _GEN_1349; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1884 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_260 : _GEN_1350; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1885 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_261 : _GEN_1351; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1886 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_262 : _GEN_1352; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1887 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_263 : _GEN_1353; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1888 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_264 : _GEN_1354; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1889 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_265 : _GEN_1355; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1890 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_266 : _GEN_1356; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1891 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_267 : _GEN_1357; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1892 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_268 : _GEN_1358; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1893 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_269 : _GEN_1359; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1894 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_270 : _GEN_1360; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1895 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_271 : _GEN_1361; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1896 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_272 : _GEN_1362; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1897 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_273 : _GEN_1363; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1898 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_274 : _GEN_1364; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1899 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_275 : _GEN_1365; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1900 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_276 : _GEN_1366; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1901 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_277 : _GEN_1367; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1902 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_278 : _GEN_1368; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1903 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_279 : _GEN_1369; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1904 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_280 : _GEN_1370; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1905 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_281 : _GEN_1371; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1906 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_282 : _GEN_1372; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1907 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_283 : _GEN_1373; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1908 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_284 : _GEN_1374; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1909 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_285 : _GEN_1375; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1910 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_286 : _GEN_1376; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1911 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_287 : _GEN_1377; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1912 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_288 : _GEN_1378; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1913 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_289 : _GEN_1379; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1914 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_290 : _GEN_1380; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1915 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_291 : _GEN_1381; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1916 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_292 : _GEN_1382; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1917 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_293 : _GEN_1383; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1918 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_294 : _GEN_1384; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1919 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_295 : _GEN_1385; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1920 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_296 : _GEN_1386; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1921 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_297 : _GEN_1387; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1922 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_298 : _GEN_1388; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1923 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_299 : _GEN_1389; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1924 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_300 : _GEN_1390; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1925 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_301 : _GEN_1391; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1926 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_302 : _GEN_1392; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1927 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_303 : _GEN_1393; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1928 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_304 : _GEN_1394; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1929 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_305 : _GEN_1395; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1930 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_306 : _GEN_1396; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1931 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_307 : _GEN_1397; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1932 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_308 : _GEN_1398; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1933 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_309 : _GEN_1399; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1934 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_310 : _GEN_1400; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1935 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_311 : _GEN_1401; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1936 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_312 : _GEN_1402; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1937 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_313 : _GEN_1403; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1938 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_314 : _GEN_1404; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1939 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_315 : _GEN_1405; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1940 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_316 : _GEN_1406; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1941 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_317 : _GEN_1407; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1942 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_318 : _GEN_1408; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1943 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_319 : _GEN_1409; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1944 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_320 : _GEN_1410; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1945 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_321 : _GEN_1411; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1946 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_322 : _GEN_1412; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1947 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_323 : _GEN_1413; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1948 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_324 : _GEN_1414; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1949 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_325 : _GEN_1415; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1950 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_326 : _GEN_1416; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1951 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_327 : _GEN_1417; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1952 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_328 : _GEN_1418; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1953 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_329 : _GEN_1419; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1954 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_330 : _GEN_1420; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1955 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_331 : _GEN_1421; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1956 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_332 : _GEN_1422; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1957 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_333 : _GEN_1423; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1958 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_334 : _GEN_1424; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1959 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_335 : _GEN_1425; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1960 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_336 : _GEN_1426; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1961 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_337 : _GEN_1427; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1962 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_338 : _GEN_1428; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1963 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_339 : _GEN_1429; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1964 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_340 : _GEN_1430; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1965 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_341 : _GEN_1431; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1966 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_342 : _GEN_1432; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1967 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_343 : _GEN_1433; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1968 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_344 : _GEN_1434; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1969 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_345 : _GEN_1435; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1970 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_346 : _GEN_1436; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1971 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_347 : _GEN_1437; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1972 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_348 : _GEN_1438; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1973 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_349 : _GEN_1439; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1974 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_350 : _GEN_1440; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1975 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_351 : _GEN_1441; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1976 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_352 : _GEN_1442; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1977 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_353 : _GEN_1443; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1978 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_354 : _GEN_1444; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1979 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_355 : _GEN_1445; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1980 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_356 : _GEN_1446; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1981 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_357 : _GEN_1447; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1982 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_358 : _GEN_1448; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1983 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_359 : _GEN_1449; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1984 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_360 : _GEN_1450; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1985 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_361 : _GEN_1451; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1986 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_362 : _GEN_1452; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1987 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_363 : _GEN_1453; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1988 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_364 : _GEN_1454; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1989 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_365 : _GEN_1455; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1990 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_366 : _GEN_1456; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1991 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_367 : _GEN_1457; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1992 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_368 : _GEN_1458; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1993 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_369 : _GEN_1459; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1994 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_370 : _GEN_1460; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1995 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_371 : _GEN_1461; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1996 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_372 : _GEN_1462; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1997 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_373 : _GEN_1463; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1998 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_374 : _GEN_1464; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1999 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_375 : _GEN_1465; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2000 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_376 : _GEN_1466; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2001 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_377 : _GEN_1467; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2002 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_378 : _GEN_1468; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2003 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_379 : _GEN_1469; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2004 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_380 : _GEN_1470; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2005 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_381 : _GEN_1471; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2006 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_382 : _GEN_1472; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2007 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_383 : _GEN_1473; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2008 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_384 : _GEN_1474; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2009 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_385 : _GEN_1475; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2010 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_386 : _GEN_1476; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2011 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_387 : _GEN_1477; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2012 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_388 : _GEN_1478; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2013 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_389 : _GEN_1479; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2014 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_390 : _GEN_1480; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2015 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_391 : _GEN_1481; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2016 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_392 : _GEN_1482; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2017 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_393 : _GEN_1483; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2018 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_394 : _GEN_1484; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2019 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_395 : _GEN_1485; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2020 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_396 : _GEN_1486; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2021 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_397 : _GEN_1487; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2022 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_398 : _GEN_1488; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2023 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_399 : _GEN_1489; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2024 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_400 : _GEN_1490; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2025 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_401 : _GEN_1491; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2026 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_402 : _GEN_1492; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2027 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_403 : _GEN_1493; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2028 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_404 : _GEN_1494; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2029 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_405 : _GEN_1495; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2030 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_406 : _GEN_1496; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2031 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_407 : _GEN_1497; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2032 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_408 : _GEN_1498; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2033 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_409 : _GEN_1499; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2034 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_410 : _GEN_1500; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2035 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_411 : _GEN_1501; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2036 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_412 : _GEN_1502; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2037 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_413 : _GEN_1503; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2038 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_414 : _GEN_1504; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2039 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_415 : _GEN_1505; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2040 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_416 : _GEN_1506; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2041 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_417 : _GEN_1507; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2042 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_418 : _GEN_1508; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2043 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_419 : _GEN_1509; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2044 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_420 : _GEN_1510; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2045 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_421 : _GEN_1511; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2046 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_422 : _GEN_1512; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2047 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_423 : _GEN_1513; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2048 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_424 : _GEN_1514; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2049 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_425 : _GEN_1515; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2050 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_426 : _GEN_1516; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2051 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_427 : _GEN_1517; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2052 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_428 : _GEN_1518; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2053 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_429 : _GEN_1519; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2054 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_430 : _GEN_1520; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2055 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_431 : _GEN_1521; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2056 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_432 : _GEN_1522; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2057 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_433 : _GEN_1523; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2058 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_434 : _GEN_1524; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2059 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_435 : _GEN_1525; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2060 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_436 : _GEN_1526; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2061 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_437 : _GEN_1527; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2062 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_438 : _GEN_1528; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2063 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_439 : _GEN_1529; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2064 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_440 : _GEN_1530; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2065 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_441 : _GEN_1531; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2066 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_442 : _GEN_1532; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2067 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_443 : _GEN_1533; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2068 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_444 : _GEN_1534; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2069 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_445 : _GEN_1535; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2070 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_446 : _GEN_1536; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2071 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_447 : _GEN_1537; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2072 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_448 : _GEN_1538; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2073 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_449 : _GEN_1539; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2074 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_450 : _GEN_1540; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2075 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_451 : _GEN_1541; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2076 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_452 : _GEN_1542; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2077 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_453 : _GEN_1543; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2078 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_454 : _GEN_1544; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2079 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_455 : _GEN_1545; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2080 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_456 : _GEN_1546; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2081 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_457 : _GEN_1547; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2082 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_458 : _GEN_1548; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2083 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_459 : _GEN_1549; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2084 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_460 : _GEN_1550; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2085 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_461 : _GEN_1551; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2086 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_462 : _GEN_1552; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2087 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_463 : _GEN_1553; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2088 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_464 : _GEN_1554; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2089 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_465 : _GEN_1555; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2090 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_466 : _GEN_1556; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2091 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_467 : _GEN_1557; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2092 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_468 : _GEN_1558; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2093 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_469 : _GEN_1559; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2094 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_470 : _GEN_1560; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2095 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_471 : _GEN_1561; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2096 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_472 : _GEN_1562; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2097 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_473 : _GEN_1563; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2098 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_474 : _GEN_1564; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2099 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_475 : _GEN_1565; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2100 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_476 : _GEN_1566; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2101 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_477 : _GEN_1567; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2102 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_478 : _GEN_1568; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2103 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_479 : _GEN_1569; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2104 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_480 : _GEN_1570; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2105 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_481 : _GEN_1571; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2106 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_482 : _GEN_1572; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2107 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_483 : _GEN_1573; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2108 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_484 : _GEN_1574; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2109 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_485 : _GEN_1575; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2110 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_486 : _GEN_1576; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2111 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_487 : _GEN_1577; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2112 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_488 : _GEN_1578; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2113 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_489 : _GEN_1579; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2114 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_490 : _GEN_1580; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2115 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_491 : _GEN_1581; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2116 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_492 : _GEN_1582; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2117 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_493 : _GEN_1583; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2118 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_494 : _GEN_1584; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2119 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_495 : _GEN_1585; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2120 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_496 : _GEN_1586; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2121 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_497 : _GEN_1587; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2122 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_498 : _GEN_1588; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2123 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_499 : _GEN_1589; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2124 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_500 : _GEN_1590; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2125 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_501 : _GEN_1591; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2126 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_502 : _GEN_1592; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2127 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_503 : _GEN_1593; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2128 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_504 : _GEN_1594; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2129 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_505 : _GEN_1595; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2130 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_506 : _GEN_1596; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2131 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_507 : _GEN_1597; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2132 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_508 : _GEN_1598; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2133 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_509 : _GEN_1599; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2134 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_510 : _GEN_1600; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2135 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_511 : _GEN_1601; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire  _GEN_2137 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_next_config_id : _GEN_1603; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [3:0] _GEN_2138 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_next_processor_id : _GEN_1604; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2158 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_0 : _GEN_1624; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2159 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_1 : _GEN_1625; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2160 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_2 : _GEN_1626; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2161 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_3 : _GEN_1627; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2162 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_4 : _GEN_1628; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2163 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_5 : _GEN_1629; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2164 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_6 : _GEN_1630; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2165 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_7 : _GEN_1631; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2166 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_8 : _GEN_1632; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2167 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_9 : _GEN_1633; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2168 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_10 : _GEN_1634; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2169 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_11 : _GEN_1635; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2170 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_12 : _GEN_1636; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2171 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_13 : _GEN_1637; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2172 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_14 : _GEN_1638; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2173 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_15 : _GEN_1639; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2174 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_16 : _GEN_1640; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2175 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_17 : _GEN_1641; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2176 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_18 : _GEN_1642; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2177 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_19 : _GEN_1643; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2178 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_20 : _GEN_1644; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2179 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_21 : _GEN_1645; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2180 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_22 : _GEN_1646; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2181 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_23 : _GEN_1647; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2182 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_24 : _GEN_1648; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2183 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_25 : _GEN_1649; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2184 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_26 : _GEN_1650; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2185 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_27 : _GEN_1651; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2186 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_28 : _GEN_1652; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2187 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_29 : _GEN_1653; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2188 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_30 : _GEN_1654; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2189 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_31 : _GEN_1655; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2190 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_32 : _GEN_1656; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2191 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_33 : _GEN_1657; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2192 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_34 : _GEN_1658; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2193 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_35 : _GEN_1659; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2194 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_36 : _GEN_1660; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2195 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_37 : _GEN_1661; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2196 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_38 : _GEN_1662; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2197 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_39 : _GEN_1663; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2198 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_40 : _GEN_1664; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2199 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_41 : _GEN_1665; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2200 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_42 : _GEN_1666; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2201 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_43 : _GEN_1667; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2202 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_44 : _GEN_1668; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2203 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_45 : _GEN_1669; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2204 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_46 : _GEN_1670; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2205 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_47 : _GEN_1671; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2206 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_48 : _GEN_1672; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2207 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_49 : _GEN_1673; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2208 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_50 : _GEN_1674; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2209 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_51 : _GEN_1675; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2210 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_52 : _GEN_1676; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2211 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_53 : _GEN_1677; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2212 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_54 : _GEN_1678; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2213 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_55 : _GEN_1679; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2214 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_56 : _GEN_1680; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2215 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_57 : _GEN_1681; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2216 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_58 : _GEN_1682; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2217 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_59 : _GEN_1683; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2218 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_60 : _GEN_1684; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2219 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_61 : _GEN_1685; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2220 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_62 : _GEN_1686; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2221 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_63 : _GEN_1687; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2222 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_64 : _GEN_1688; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2223 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_65 : _GEN_1689; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2224 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_66 : _GEN_1690; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2225 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_67 : _GEN_1691; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2226 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_68 : _GEN_1692; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2227 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_69 : _GEN_1693; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2228 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_70 : _GEN_1694; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2229 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_71 : _GEN_1695; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2230 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_72 : _GEN_1696; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2231 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_73 : _GEN_1697; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2232 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_74 : _GEN_1698; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2233 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_75 : _GEN_1699; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2234 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_76 : _GEN_1700; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2235 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_77 : _GEN_1701; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2236 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_78 : _GEN_1702; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2237 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_79 : _GEN_1703; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2238 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_80 : _GEN_1704; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2239 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_81 : _GEN_1705; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2240 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_82 : _GEN_1706; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2241 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_83 : _GEN_1707; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2242 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_84 : _GEN_1708; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2243 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_85 : _GEN_1709; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2244 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_86 : _GEN_1710; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2245 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_87 : _GEN_1711; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2246 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_88 : _GEN_1712; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2247 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_89 : _GEN_1713; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2248 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_90 : _GEN_1714; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2249 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_91 : _GEN_1715; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2250 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_92 : _GEN_1716; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2251 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_93 : _GEN_1717; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2252 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_94 : _GEN_1718; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2253 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_95 : _GEN_1719; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2254 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_96 : _GEN_1720; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2255 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_97 : _GEN_1721; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2256 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_98 : _GEN_1722; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2257 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_99 : _GEN_1723; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2258 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_100 : _GEN_1724; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2259 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_101 : _GEN_1725; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2260 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_102 : _GEN_1726; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2261 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_103 : _GEN_1727; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2262 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_104 : _GEN_1728; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2263 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_105 : _GEN_1729; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2264 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_106 : _GEN_1730; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2265 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_107 : _GEN_1731; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2266 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_108 : _GEN_1732; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2267 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_109 : _GEN_1733; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2268 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_110 : _GEN_1734; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2269 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_111 : _GEN_1735; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2270 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_112 : _GEN_1736; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2271 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_113 : _GEN_1737; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2272 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_114 : _GEN_1738; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2273 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_115 : _GEN_1739; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2274 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_116 : _GEN_1740; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2275 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_117 : _GEN_1741; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2276 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_118 : _GEN_1742; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2277 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_119 : _GEN_1743; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2278 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_120 : _GEN_1744; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2279 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_121 : _GEN_1745; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2280 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_122 : _GEN_1746; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2281 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_123 : _GEN_1747; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2282 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_124 : _GEN_1748; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2283 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_125 : _GEN_1749; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2284 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_126 : _GEN_1750; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2285 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_127 : _GEN_1751; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2286 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_128 : _GEN_1752; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2287 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_129 : _GEN_1753; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2288 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_130 : _GEN_1754; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2289 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_131 : _GEN_1755; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2290 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_132 : _GEN_1756; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2291 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_133 : _GEN_1757; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2292 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_134 : _GEN_1758; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2293 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_135 : _GEN_1759; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2294 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_136 : _GEN_1760; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2295 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_137 : _GEN_1761; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2296 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_138 : _GEN_1762; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2297 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_139 : _GEN_1763; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2298 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_140 : _GEN_1764; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2299 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_141 : _GEN_1765; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2300 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_142 : _GEN_1766; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2301 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_143 : _GEN_1767; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2302 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_144 : _GEN_1768; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2303 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_145 : _GEN_1769; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2304 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_146 : _GEN_1770; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2305 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_147 : _GEN_1771; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2306 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_148 : _GEN_1772; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2307 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_149 : _GEN_1773; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2308 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_150 : _GEN_1774; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2309 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_151 : _GEN_1775; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2310 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_152 : _GEN_1776; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2311 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_153 : _GEN_1777; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2312 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_154 : _GEN_1778; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2313 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_155 : _GEN_1779; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2314 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_156 : _GEN_1780; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2315 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_157 : _GEN_1781; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2316 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_158 : _GEN_1782; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2317 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_159 : _GEN_1783; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2318 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_160 : _GEN_1784; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2319 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_161 : _GEN_1785; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2320 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_162 : _GEN_1786; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2321 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_163 : _GEN_1787; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2322 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_164 : _GEN_1788; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2323 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_165 : _GEN_1789; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2324 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_166 : _GEN_1790; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2325 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_167 : _GEN_1791; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2326 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_168 : _GEN_1792; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2327 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_169 : _GEN_1793; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2328 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_170 : _GEN_1794; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2329 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_171 : _GEN_1795; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2330 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_172 : _GEN_1796; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2331 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_173 : _GEN_1797; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2332 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_174 : _GEN_1798; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2333 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_175 : _GEN_1799; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2334 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_176 : _GEN_1800; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2335 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_177 : _GEN_1801; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2336 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_178 : _GEN_1802; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2337 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_179 : _GEN_1803; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2338 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_180 : _GEN_1804; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2339 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_181 : _GEN_1805; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2340 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_182 : _GEN_1806; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2341 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_183 : _GEN_1807; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2342 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_184 : _GEN_1808; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2343 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_185 : _GEN_1809; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2344 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_186 : _GEN_1810; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2345 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_187 : _GEN_1811; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2346 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_188 : _GEN_1812; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2347 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_189 : _GEN_1813; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2348 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_190 : _GEN_1814; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2349 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_191 : _GEN_1815; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2350 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_192 : _GEN_1816; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2351 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_193 : _GEN_1817; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2352 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_194 : _GEN_1818; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2353 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_195 : _GEN_1819; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2354 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_196 : _GEN_1820; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2355 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_197 : _GEN_1821; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2356 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_198 : _GEN_1822; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2357 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_199 : _GEN_1823; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2358 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_200 : _GEN_1824; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2359 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_201 : _GEN_1825; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2360 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_202 : _GEN_1826; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2361 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_203 : _GEN_1827; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2362 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_204 : _GEN_1828; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2363 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_205 : _GEN_1829; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2364 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_206 : _GEN_1830; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2365 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_207 : _GEN_1831; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2366 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_208 : _GEN_1832; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2367 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_209 : _GEN_1833; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2368 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_210 : _GEN_1834; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2369 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_211 : _GEN_1835; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2370 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_212 : _GEN_1836; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2371 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_213 : _GEN_1837; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2372 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_214 : _GEN_1838; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2373 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_215 : _GEN_1839; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2374 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_216 : _GEN_1840; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2375 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_217 : _GEN_1841; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2376 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_218 : _GEN_1842; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2377 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_219 : _GEN_1843; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2378 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_220 : _GEN_1844; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2379 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_221 : _GEN_1845; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2380 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_222 : _GEN_1846; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2381 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_223 : _GEN_1847; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2382 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_224 : _GEN_1848; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2383 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_225 : _GEN_1849; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2384 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_226 : _GEN_1850; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2385 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_227 : _GEN_1851; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2386 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_228 : _GEN_1852; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2387 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_229 : _GEN_1853; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2388 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_230 : _GEN_1854; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2389 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_231 : _GEN_1855; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2390 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_232 : _GEN_1856; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2391 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_233 : _GEN_1857; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2392 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_234 : _GEN_1858; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2393 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_235 : _GEN_1859; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2394 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_236 : _GEN_1860; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2395 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_237 : _GEN_1861; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2396 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_238 : _GEN_1862; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2397 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_239 : _GEN_1863; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2398 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_240 : _GEN_1864; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2399 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_241 : _GEN_1865; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2400 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_242 : _GEN_1866; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2401 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_243 : _GEN_1867; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2402 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_244 : _GEN_1868; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2403 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_245 : _GEN_1869; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2404 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_246 : _GEN_1870; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2405 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_247 : _GEN_1871; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2406 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_248 : _GEN_1872; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2407 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_249 : _GEN_1873; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2408 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_250 : _GEN_1874; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2409 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_251 : _GEN_1875; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2410 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_252 : _GEN_1876; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2411 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_253 : _GEN_1877; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2412 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_254 : _GEN_1878; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2413 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_255 : _GEN_1879; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2414 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_256 : _GEN_1880; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2415 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_257 : _GEN_1881; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2416 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_258 : _GEN_1882; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2417 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_259 : _GEN_1883; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2418 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_260 : _GEN_1884; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2419 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_261 : _GEN_1885; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2420 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_262 : _GEN_1886; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2421 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_263 : _GEN_1887; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2422 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_264 : _GEN_1888; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2423 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_265 : _GEN_1889; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2424 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_266 : _GEN_1890; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2425 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_267 : _GEN_1891; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2426 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_268 : _GEN_1892; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2427 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_269 : _GEN_1893; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2428 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_270 : _GEN_1894; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2429 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_271 : _GEN_1895; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2430 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_272 : _GEN_1896; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2431 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_273 : _GEN_1897; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2432 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_274 : _GEN_1898; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2433 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_275 : _GEN_1899; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2434 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_276 : _GEN_1900; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2435 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_277 : _GEN_1901; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2436 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_278 : _GEN_1902; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2437 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_279 : _GEN_1903; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2438 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_280 : _GEN_1904; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2439 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_281 : _GEN_1905; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2440 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_282 : _GEN_1906; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2441 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_283 : _GEN_1907; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2442 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_284 : _GEN_1908; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2443 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_285 : _GEN_1909; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2444 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_286 : _GEN_1910; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2445 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_287 : _GEN_1911; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2446 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_288 : _GEN_1912; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2447 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_289 : _GEN_1913; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2448 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_290 : _GEN_1914; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2449 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_291 : _GEN_1915; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2450 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_292 : _GEN_1916; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2451 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_293 : _GEN_1917; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2452 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_294 : _GEN_1918; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2453 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_295 : _GEN_1919; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2454 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_296 : _GEN_1920; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2455 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_297 : _GEN_1921; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2456 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_298 : _GEN_1922; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2457 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_299 : _GEN_1923; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2458 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_300 : _GEN_1924; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2459 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_301 : _GEN_1925; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2460 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_302 : _GEN_1926; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2461 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_303 : _GEN_1927; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2462 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_304 : _GEN_1928; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2463 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_305 : _GEN_1929; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2464 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_306 : _GEN_1930; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2465 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_307 : _GEN_1931; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2466 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_308 : _GEN_1932; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2467 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_309 : _GEN_1933; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2468 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_310 : _GEN_1934; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2469 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_311 : _GEN_1935; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2470 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_312 : _GEN_1936; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2471 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_313 : _GEN_1937; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2472 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_314 : _GEN_1938; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2473 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_315 : _GEN_1939; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2474 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_316 : _GEN_1940; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2475 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_317 : _GEN_1941; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2476 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_318 : _GEN_1942; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2477 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_319 : _GEN_1943; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2478 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_320 : _GEN_1944; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2479 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_321 : _GEN_1945; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2480 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_322 : _GEN_1946; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2481 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_323 : _GEN_1947; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2482 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_324 : _GEN_1948; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2483 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_325 : _GEN_1949; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2484 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_326 : _GEN_1950; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2485 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_327 : _GEN_1951; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2486 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_328 : _GEN_1952; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2487 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_329 : _GEN_1953; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2488 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_330 : _GEN_1954; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2489 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_331 : _GEN_1955; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2490 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_332 : _GEN_1956; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2491 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_333 : _GEN_1957; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2492 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_334 : _GEN_1958; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2493 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_335 : _GEN_1959; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2494 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_336 : _GEN_1960; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2495 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_337 : _GEN_1961; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2496 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_338 : _GEN_1962; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2497 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_339 : _GEN_1963; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2498 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_340 : _GEN_1964; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2499 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_341 : _GEN_1965; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2500 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_342 : _GEN_1966; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2501 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_343 : _GEN_1967; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2502 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_344 : _GEN_1968; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2503 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_345 : _GEN_1969; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2504 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_346 : _GEN_1970; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2505 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_347 : _GEN_1971; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2506 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_348 : _GEN_1972; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2507 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_349 : _GEN_1973; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2508 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_350 : _GEN_1974; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2509 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_351 : _GEN_1975; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2510 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_352 : _GEN_1976; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2511 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_353 : _GEN_1977; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2512 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_354 : _GEN_1978; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2513 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_355 : _GEN_1979; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2514 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_356 : _GEN_1980; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2515 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_357 : _GEN_1981; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2516 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_358 : _GEN_1982; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2517 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_359 : _GEN_1983; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2518 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_360 : _GEN_1984; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2519 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_361 : _GEN_1985; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2520 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_362 : _GEN_1986; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2521 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_363 : _GEN_1987; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2522 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_364 : _GEN_1988; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2523 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_365 : _GEN_1989; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2524 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_366 : _GEN_1990; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2525 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_367 : _GEN_1991; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2526 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_368 : _GEN_1992; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2527 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_369 : _GEN_1993; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2528 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_370 : _GEN_1994; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2529 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_371 : _GEN_1995; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2530 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_372 : _GEN_1996; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2531 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_373 : _GEN_1997; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2532 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_374 : _GEN_1998; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2533 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_375 : _GEN_1999; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2534 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_376 : _GEN_2000; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2535 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_377 : _GEN_2001; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2536 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_378 : _GEN_2002; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2537 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_379 : _GEN_2003; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2538 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_380 : _GEN_2004; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2539 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_381 : _GEN_2005; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2540 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_382 : _GEN_2006; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2541 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_383 : _GEN_2007; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2542 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_384 : _GEN_2008; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2543 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_385 : _GEN_2009; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2544 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_386 : _GEN_2010; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2545 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_387 : _GEN_2011; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2546 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_388 : _GEN_2012; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2547 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_389 : _GEN_2013; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2548 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_390 : _GEN_2014; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2549 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_391 : _GEN_2015; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2550 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_392 : _GEN_2016; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2551 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_393 : _GEN_2017; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2552 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_394 : _GEN_2018; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2553 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_395 : _GEN_2019; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2554 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_396 : _GEN_2020; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2555 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_397 : _GEN_2021; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2556 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_398 : _GEN_2022; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2557 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_399 : _GEN_2023; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2558 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_400 : _GEN_2024; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2559 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_401 : _GEN_2025; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2560 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_402 : _GEN_2026; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2561 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_403 : _GEN_2027; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2562 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_404 : _GEN_2028; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2563 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_405 : _GEN_2029; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2564 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_406 : _GEN_2030; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2565 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_407 : _GEN_2031; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2566 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_408 : _GEN_2032; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2567 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_409 : _GEN_2033; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2568 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_410 : _GEN_2034; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2569 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_411 : _GEN_2035; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2570 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_412 : _GEN_2036; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2571 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_413 : _GEN_2037; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2572 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_414 : _GEN_2038; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2573 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_415 : _GEN_2039; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2574 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_416 : _GEN_2040; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2575 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_417 : _GEN_2041; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2576 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_418 : _GEN_2042; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2577 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_419 : _GEN_2043; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2578 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_420 : _GEN_2044; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2579 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_421 : _GEN_2045; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2580 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_422 : _GEN_2046; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2581 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_423 : _GEN_2047; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2582 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_424 : _GEN_2048; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2583 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_425 : _GEN_2049; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2584 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_426 : _GEN_2050; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2585 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_427 : _GEN_2051; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2586 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_428 : _GEN_2052; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2587 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_429 : _GEN_2053; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2588 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_430 : _GEN_2054; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2589 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_431 : _GEN_2055; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2590 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_432 : _GEN_2056; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2591 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_433 : _GEN_2057; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2592 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_434 : _GEN_2058; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2593 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_435 : _GEN_2059; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2594 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_436 : _GEN_2060; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2595 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_437 : _GEN_2061; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2596 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_438 : _GEN_2062; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2597 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_439 : _GEN_2063; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2598 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_440 : _GEN_2064; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2599 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_441 : _GEN_2065; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2600 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_442 : _GEN_2066; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2601 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_443 : _GEN_2067; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2602 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_444 : _GEN_2068; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2603 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_445 : _GEN_2069; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2604 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_446 : _GEN_2070; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2605 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_447 : _GEN_2071; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2606 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_448 : _GEN_2072; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2607 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_449 : _GEN_2073; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2608 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_450 : _GEN_2074; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2609 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_451 : _GEN_2075; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2610 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_452 : _GEN_2076; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2611 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_453 : _GEN_2077; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2612 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_454 : _GEN_2078; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2613 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_455 : _GEN_2079; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2614 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_456 : _GEN_2080; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2615 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_457 : _GEN_2081; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2616 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_458 : _GEN_2082; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2617 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_459 : _GEN_2083; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2618 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_460 : _GEN_2084; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2619 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_461 : _GEN_2085; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2620 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_462 : _GEN_2086; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2621 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_463 : _GEN_2087; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2622 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_464 : _GEN_2088; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2623 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_465 : _GEN_2089; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2624 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_466 : _GEN_2090; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2625 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_467 : _GEN_2091; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2626 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_468 : _GEN_2092; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2627 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_469 : _GEN_2093; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2628 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_470 : _GEN_2094; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2629 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_471 : _GEN_2095; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2630 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_472 : _GEN_2096; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2631 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_473 : _GEN_2097; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2632 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_474 : _GEN_2098; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2633 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_475 : _GEN_2099; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2634 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_476 : _GEN_2100; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2635 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_477 : _GEN_2101; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2636 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_478 : _GEN_2102; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2637 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_479 : _GEN_2103; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2638 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_480 : _GEN_2104; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2639 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_481 : _GEN_2105; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2640 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_482 : _GEN_2106; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2641 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_483 : _GEN_2107; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2642 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_484 : _GEN_2108; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2643 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_485 : _GEN_2109; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2644 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_486 : _GEN_2110; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2645 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_487 : _GEN_2111; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2646 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_488 : _GEN_2112; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2647 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_489 : _GEN_2113; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2648 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_490 : _GEN_2114; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2649 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_491 : _GEN_2115; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2650 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_492 : _GEN_2116; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2651 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_493 : _GEN_2117; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2652 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_494 : _GEN_2118; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2653 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_495 : _GEN_2119; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2654 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_496 : _GEN_2120; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2655 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_497 : _GEN_2121; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2656 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_498 : _GEN_2122; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2657 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_499 : _GEN_2123; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2658 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_500 : _GEN_2124; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2659 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_501 : _GEN_2125; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2660 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_502 : _GEN_2126; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2661 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_503 : _GEN_2127; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2662 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_504 : _GEN_2128; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2663 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_505 : _GEN_2129; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2664 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_506 : _GEN_2130; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2665 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_507 : _GEN_2131; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2666 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_508 : _GEN_2132; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2667 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_509 : _GEN_2133; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2668 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_510 : _GEN_2134; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2669 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_511 : _GEN_2135; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire  _GEN_2671 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_next_config_id : _GEN_2137; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [3:0] _GEN_2672 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_next_processor_id : _GEN_2138; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2692 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_0 : _GEN_2158; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2693 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_1 : _GEN_2159; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2694 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_2 : _GEN_2160; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2695 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_3 : _GEN_2161; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2696 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_4 : _GEN_2162; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2697 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_5 : _GEN_2163; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2698 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_6 : _GEN_2164; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2699 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_7 : _GEN_2165; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2700 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_8 : _GEN_2166; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2701 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_9 : _GEN_2167; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2702 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_10 : _GEN_2168; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2703 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_11 : _GEN_2169; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2704 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_12 : _GEN_2170; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2705 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_13 : _GEN_2171; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2706 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_14 : _GEN_2172; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2707 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_15 : _GEN_2173; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2708 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_16 : _GEN_2174; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2709 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_17 : _GEN_2175; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2710 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_18 : _GEN_2176; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2711 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_19 : _GEN_2177; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2712 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_20 : _GEN_2178; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2713 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_21 : _GEN_2179; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2714 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_22 : _GEN_2180; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2715 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_23 : _GEN_2181; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2716 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_24 : _GEN_2182; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2717 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_25 : _GEN_2183; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2718 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_26 : _GEN_2184; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2719 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_27 : _GEN_2185; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2720 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_28 : _GEN_2186; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2721 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_29 : _GEN_2187; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2722 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_30 : _GEN_2188; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2723 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_31 : _GEN_2189; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2724 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_32 : _GEN_2190; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2725 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_33 : _GEN_2191; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2726 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_34 : _GEN_2192; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2727 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_35 : _GEN_2193; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2728 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_36 : _GEN_2194; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2729 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_37 : _GEN_2195; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2730 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_38 : _GEN_2196; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2731 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_39 : _GEN_2197; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2732 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_40 : _GEN_2198; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2733 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_41 : _GEN_2199; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2734 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_42 : _GEN_2200; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2735 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_43 : _GEN_2201; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2736 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_44 : _GEN_2202; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2737 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_45 : _GEN_2203; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2738 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_46 : _GEN_2204; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2739 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_47 : _GEN_2205; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2740 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_48 : _GEN_2206; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2741 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_49 : _GEN_2207; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2742 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_50 : _GEN_2208; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2743 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_51 : _GEN_2209; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2744 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_52 : _GEN_2210; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2745 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_53 : _GEN_2211; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2746 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_54 : _GEN_2212; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2747 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_55 : _GEN_2213; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2748 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_56 : _GEN_2214; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2749 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_57 : _GEN_2215; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2750 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_58 : _GEN_2216; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2751 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_59 : _GEN_2217; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2752 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_60 : _GEN_2218; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2753 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_61 : _GEN_2219; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2754 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_62 : _GEN_2220; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2755 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_63 : _GEN_2221; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2756 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_64 : _GEN_2222; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2757 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_65 : _GEN_2223; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2758 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_66 : _GEN_2224; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2759 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_67 : _GEN_2225; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2760 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_68 : _GEN_2226; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2761 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_69 : _GEN_2227; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2762 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_70 : _GEN_2228; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2763 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_71 : _GEN_2229; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2764 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_72 : _GEN_2230; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2765 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_73 : _GEN_2231; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2766 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_74 : _GEN_2232; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2767 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_75 : _GEN_2233; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2768 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_76 : _GEN_2234; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2769 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_77 : _GEN_2235; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2770 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_78 : _GEN_2236; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2771 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_79 : _GEN_2237; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2772 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_80 : _GEN_2238; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2773 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_81 : _GEN_2239; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2774 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_82 : _GEN_2240; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2775 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_83 : _GEN_2241; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2776 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_84 : _GEN_2242; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2777 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_85 : _GEN_2243; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2778 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_86 : _GEN_2244; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2779 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_87 : _GEN_2245; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2780 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_88 : _GEN_2246; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2781 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_89 : _GEN_2247; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2782 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_90 : _GEN_2248; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2783 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_91 : _GEN_2249; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2784 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_92 : _GEN_2250; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2785 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_93 : _GEN_2251; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2786 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_94 : _GEN_2252; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2787 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_95 : _GEN_2253; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2788 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_96 : _GEN_2254; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2789 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_97 : _GEN_2255; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2790 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_98 : _GEN_2256; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2791 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_99 : _GEN_2257; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2792 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_100 : _GEN_2258; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2793 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_101 : _GEN_2259; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2794 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_102 : _GEN_2260; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2795 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_103 : _GEN_2261; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2796 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_104 : _GEN_2262; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2797 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_105 : _GEN_2263; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2798 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_106 : _GEN_2264; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2799 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_107 : _GEN_2265; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2800 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_108 : _GEN_2266; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2801 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_109 : _GEN_2267; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2802 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_110 : _GEN_2268; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2803 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_111 : _GEN_2269; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2804 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_112 : _GEN_2270; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2805 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_113 : _GEN_2271; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2806 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_114 : _GEN_2272; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2807 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_115 : _GEN_2273; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2808 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_116 : _GEN_2274; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2809 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_117 : _GEN_2275; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2810 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_118 : _GEN_2276; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2811 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_119 : _GEN_2277; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2812 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_120 : _GEN_2278; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2813 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_121 : _GEN_2279; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2814 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_122 : _GEN_2280; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2815 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_123 : _GEN_2281; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2816 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_124 : _GEN_2282; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2817 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_125 : _GEN_2283; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2818 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_126 : _GEN_2284; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2819 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_127 : _GEN_2285; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2820 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_128 : _GEN_2286; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2821 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_129 : _GEN_2287; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2822 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_130 : _GEN_2288; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2823 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_131 : _GEN_2289; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2824 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_132 : _GEN_2290; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2825 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_133 : _GEN_2291; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2826 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_134 : _GEN_2292; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2827 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_135 : _GEN_2293; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2828 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_136 : _GEN_2294; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2829 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_137 : _GEN_2295; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2830 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_138 : _GEN_2296; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2831 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_139 : _GEN_2297; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2832 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_140 : _GEN_2298; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2833 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_141 : _GEN_2299; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2834 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_142 : _GEN_2300; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2835 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_143 : _GEN_2301; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2836 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_144 : _GEN_2302; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2837 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_145 : _GEN_2303; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2838 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_146 : _GEN_2304; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2839 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_147 : _GEN_2305; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2840 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_148 : _GEN_2306; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2841 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_149 : _GEN_2307; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2842 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_150 : _GEN_2308; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2843 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_151 : _GEN_2309; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2844 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_152 : _GEN_2310; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2845 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_153 : _GEN_2311; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2846 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_154 : _GEN_2312; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2847 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_155 : _GEN_2313; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2848 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_156 : _GEN_2314; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2849 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_157 : _GEN_2315; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2850 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_158 : _GEN_2316; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2851 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_159 : _GEN_2317; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2852 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_160 : _GEN_2318; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2853 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_161 : _GEN_2319; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2854 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_162 : _GEN_2320; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2855 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_163 : _GEN_2321; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2856 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_164 : _GEN_2322; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2857 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_165 : _GEN_2323; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2858 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_166 : _GEN_2324; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2859 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_167 : _GEN_2325; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2860 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_168 : _GEN_2326; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2861 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_169 : _GEN_2327; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2862 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_170 : _GEN_2328; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2863 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_171 : _GEN_2329; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2864 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_172 : _GEN_2330; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2865 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_173 : _GEN_2331; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2866 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_174 : _GEN_2332; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2867 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_175 : _GEN_2333; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2868 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_176 : _GEN_2334; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2869 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_177 : _GEN_2335; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2870 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_178 : _GEN_2336; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2871 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_179 : _GEN_2337; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2872 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_180 : _GEN_2338; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2873 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_181 : _GEN_2339; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2874 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_182 : _GEN_2340; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2875 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_183 : _GEN_2341; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2876 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_184 : _GEN_2342; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2877 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_185 : _GEN_2343; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2878 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_186 : _GEN_2344; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2879 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_187 : _GEN_2345; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2880 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_188 : _GEN_2346; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2881 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_189 : _GEN_2347; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2882 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_190 : _GEN_2348; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2883 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_191 : _GEN_2349; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2884 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_192 : _GEN_2350; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2885 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_193 : _GEN_2351; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2886 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_194 : _GEN_2352; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2887 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_195 : _GEN_2353; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2888 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_196 : _GEN_2354; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2889 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_197 : _GEN_2355; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2890 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_198 : _GEN_2356; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2891 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_199 : _GEN_2357; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2892 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_200 : _GEN_2358; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2893 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_201 : _GEN_2359; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2894 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_202 : _GEN_2360; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2895 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_203 : _GEN_2361; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2896 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_204 : _GEN_2362; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2897 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_205 : _GEN_2363; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2898 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_206 : _GEN_2364; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2899 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_207 : _GEN_2365; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2900 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_208 : _GEN_2366; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2901 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_209 : _GEN_2367; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2902 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_210 : _GEN_2368; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2903 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_211 : _GEN_2369; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2904 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_212 : _GEN_2370; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2905 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_213 : _GEN_2371; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2906 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_214 : _GEN_2372; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2907 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_215 : _GEN_2373; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2908 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_216 : _GEN_2374; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2909 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_217 : _GEN_2375; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2910 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_218 : _GEN_2376; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2911 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_219 : _GEN_2377; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2912 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_220 : _GEN_2378; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2913 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_221 : _GEN_2379; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2914 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_222 : _GEN_2380; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2915 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_223 : _GEN_2381; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2916 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_224 : _GEN_2382; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2917 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_225 : _GEN_2383; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2918 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_226 : _GEN_2384; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2919 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_227 : _GEN_2385; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2920 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_228 : _GEN_2386; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2921 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_229 : _GEN_2387; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2922 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_230 : _GEN_2388; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2923 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_231 : _GEN_2389; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2924 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_232 : _GEN_2390; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2925 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_233 : _GEN_2391; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2926 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_234 : _GEN_2392; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2927 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_235 : _GEN_2393; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2928 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_236 : _GEN_2394; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2929 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_237 : _GEN_2395; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2930 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_238 : _GEN_2396; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2931 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_239 : _GEN_2397; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2932 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_240 : _GEN_2398; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2933 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_241 : _GEN_2399; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2934 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_242 : _GEN_2400; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2935 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_243 : _GEN_2401; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2936 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_244 : _GEN_2402; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2937 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_245 : _GEN_2403; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2938 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_246 : _GEN_2404; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2939 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_247 : _GEN_2405; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2940 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_248 : _GEN_2406; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2941 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_249 : _GEN_2407; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2942 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_250 : _GEN_2408; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2943 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_251 : _GEN_2409; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2944 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_252 : _GEN_2410; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2945 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_253 : _GEN_2411; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2946 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_254 : _GEN_2412; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2947 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_255 : _GEN_2413; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2948 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_256 : _GEN_2414; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2949 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_257 : _GEN_2415; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2950 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_258 : _GEN_2416; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2951 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_259 : _GEN_2417; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2952 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_260 : _GEN_2418; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2953 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_261 : _GEN_2419; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2954 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_262 : _GEN_2420; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2955 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_263 : _GEN_2421; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2956 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_264 : _GEN_2422; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2957 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_265 : _GEN_2423; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2958 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_266 : _GEN_2424; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2959 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_267 : _GEN_2425; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2960 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_268 : _GEN_2426; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2961 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_269 : _GEN_2427; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2962 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_270 : _GEN_2428; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2963 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_271 : _GEN_2429; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2964 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_272 : _GEN_2430; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2965 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_273 : _GEN_2431; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2966 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_274 : _GEN_2432; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2967 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_275 : _GEN_2433; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2968 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_276 : _GEN_2434; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2969 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_277 : _GEN_2435; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2970 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_278 : _GEN_2436; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2971 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_279 : _GEN_2437; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2972 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_280 : _GEN_2438; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2973 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_281 : _GEN_2439; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2974 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_282 : _GEN_2440; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2975 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_283 : _GEN_2441; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2976 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_284 : _GEN_2442; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2977 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_285 : _GEN_2443; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2978 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_286 : _GEN_2444; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2979 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_287 : _GEN_2445; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2980 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_288 : _GEN_2446; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2981 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_289 : _GEN_2447; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2982 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_290 : _GEN_2448; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2983 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_291 : _GEN_2449; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2984 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_292 : _GEN_2450; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2985 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_293 : _GEN_2451; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2986 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_294 : _GEN_2452; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2987 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_295 : _GEN_2453; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2988 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_296 : _GEN_2454; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2989 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_297 : _GEN_2455; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2990 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_298 : _GEN_2456; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2991 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_299 : _GEN_2457; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2992 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_300 : _GEN_2458; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2993 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_301 : _GEN_2459; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2994 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_302 : _GEN_2460; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2995 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_303 : _GEN_2461; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2996 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_304 : _GEN_2462; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2997 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_305 : _GEN_2463; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2998 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_306 : _GEN_2464; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_2999 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_307 : _GEN_2465; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3000 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_308 : _GEN_2466; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3001 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_309 : _GEN_2467; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3002 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_310 : _GEN_2468; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3003 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_311 : _GEN_2469; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3004 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_312 : _GEN_2470; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3005 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_313 : _GEN_2471; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3006 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_314 : _GEN_2472; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3007 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_315 : _GEN_2473; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3008 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_316 : _GEN_2474; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3009 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_317 : _GEN_2475; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3010 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_318 : _GEN_2476; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3011 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_319 : _GEN_2477; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3012 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_320 : _GEN_2478; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3013 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_321 : _GEN_2479; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3014 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_322 : _GEN_2480; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3015 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_323 : _GEN_2481; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3016 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_324 : _GEN_2482; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3017 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_325 : _GEN_2483; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3018 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_326 : _GEN_2484; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3019 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_327 : _GEN_2485; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3020 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_328 : _GEN_2486; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3021 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_329 : _GEN_2487; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3022 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_330 : _GEN_2488; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3023 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_331 : _GEN_2489; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3024 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_332 : _GEN_2490; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3025 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_333 : _GEN_2491; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3026 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_334 : _GEN_2492; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3027 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_335 : _GEN_2493; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3028 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_336 : _GEN_2494; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3029 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_337 : _GEN_2495; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3030 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_338 : _GEN_2496; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3031 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_339 : _GEN_2497; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3032 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_340 : _GEN_2498; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3033 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_341 : _GEN_2499; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3034 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_342 : _GEN_2500; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3035 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_343 : _GEN_2501; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3036 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_344 : _GEN_2502; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3037 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_345 : _GEN_2503; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3038 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_346 : _GEN_2504; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3039 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_347 : _GEN_2505; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3040 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_348 : _GEN_2506; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3041 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_349 : _GEN_2507; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3042 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_350 : _GEN_2508; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3043 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_351 : _GEN_2509; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3044 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_352 : _GEN_2510; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3045 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_353 : _GEN_2511; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3046 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_354 : _GEN_2512; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3047 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_355 : _GEN_2513; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3048 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_356 : _GEN_2514; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3049 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_357 : _GEN_2515; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3050 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_358 : _GEN_2516; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3051 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_359 : _GEN_2517; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3052 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_360 : _GEN_2518; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3053 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_361 : _GEN_2519; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3054 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_362 : _GEN_2520; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3055 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_363 : _GEN_2521; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3056 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_364 : _GEN_2522; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3057 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_365 : _GEN_2523; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3058 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_366 : _GEN_2524; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3059 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_367 : _GEN_2525; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3060 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_368 : _GEN_2526; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3061 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_369 : _GEN_2527; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3062 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_370 : _GEN_2528; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3063 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_371 : _GEN_2529; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3064 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_372 : _GEN_2530; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3065 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_373 : _GEN_2531; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3066 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_374 : _GEN_2532; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3067 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_375 : _GEN_2533; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3068 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_376 : _GEN_2534; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3069 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_377 : _GEN_2535; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3070 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_378 : _GEN_2536; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3071 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_379 : _GEN_2537; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3072 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_380 : _GEN_2538; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3073 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_381 : _GEN_2539; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3074 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_382 : _GEN_2540; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3075 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_383 : _GEN_2541; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3076 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_384 : _GEN_2542; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3077 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_385 : _GEN_2543; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3078 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_386 : _GEN_2544; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3079 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_387 : _GEN_2545; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3080 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_388 : _GEN_2546; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3081 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_389 : _GEN_2547; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3082 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_390 : _GEN_2548; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3083 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_391 : _GEN_2549; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3084 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_392 : _GEN_2550; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3085 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_393 : _GEN_2551; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3086 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_394 : _GEN_2552; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3087 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_395 : _GEN_2553; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3088 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_396 : _GEN_2554; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3089 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_397 : _GEN_2555; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3090 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_398 : _GEN_2556; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3091 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_399 : _GEN_2557; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3092 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_400 : _GEN_2558; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3093 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_401 : _GEN_2559; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3094 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_402 : _GEN_2560; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3095 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_403 : _GEN_2561; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3096 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_404 : _GEN_2562; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3097 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_405 : _GEN_2563; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3098 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_406 : _GEN_2564; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3099 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_407 : _GEN_2565; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3100 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_408 : _GEN_2566; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3101 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_409 : _GEN_2567; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3102 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_410 : _GEN_2568; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3103 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_411 : _GEN_2569; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3104 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_412 : _GEN_2570; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3105 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_413 : _GEN_2571; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3106 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_414 : _GEN_2572; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3107 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_415 : _GEN_2573; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3108 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_416 : _GEN_2574; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3109 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_417 : _GEN_2575; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3110 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_418 : _GEN_2576; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3111 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_419 : _GEN_2577; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3112 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_420 : _GEN_2578; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3113 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_421 : _GEN_2579; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3114 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_422 : _GEN_2580; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3115 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_423 : _GEN_2581; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3116 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_424 : _GEN_2582; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3117 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_425 : _GEN_2583; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3118 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_426 : _GEN_2584; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3119 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_427 : _GEN_2585; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3120 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_428 : _GEN_2586; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3121 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_429 : _GEN_2587; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3122 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_430 : _GEN_2588; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3123 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_431 : _GEN_2589; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3124 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_432 : _GEN_2590; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3125 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_433 : _GEN_2591; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3126 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_434 : _GEN_2592; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3127 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_435 : _GEN_2593; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3128 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_436 : _GEN_2594; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3129 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_437 : _GEN_2595; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3130 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_438 : _GEN_2596; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3131 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_439 : _GEN_2597; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3132 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_440 : _GEN_2598; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3133 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_441 : _GEN_2599; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3134 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_442 : _GEN_2600; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3135 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_443 : _GEN_2601; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3136 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_444 : _GEN_2602; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3137 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_445 : _GEN_2603; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3138 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_446 : _GEN_2604; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3139 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_447 : _GEN_2605; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3140 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_448 : _GEN_2606; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3141 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_449 : _GEN_2607; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3142 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_450 : _GEN_2608; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3143 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_451 : _GEN_2609; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3144 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_452 : _GEN_2610; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3145 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_453 : _GEN_2611; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3146 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_454 : _GEN_2612; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3147 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_455 : _GEN_2613; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3148 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_456 : _GEN_2614; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3149 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_457 : _GEN_2615; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3150 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_458 : _GEN_2616; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3151 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_459 : _GEN_2617; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3152 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_460 : _GEN_2618; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3153 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_461 : _GEN_2619; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3154 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_462 : _GEN_2620; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3155 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_463 : _GEN_2621; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3156 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_464 : _GEN_2622; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3157 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_465 : _GEN_2623; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3158 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_466 : _GEN_2624; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3159 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_467 : _GEN_2625; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3160 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_468 : _GEN_2626; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3161 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_469 : _GEN_2627; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3162 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_470 : _GEN_2628; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3163 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_471 : _GEN_2629; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3164 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_472 : _GEN_2630; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3165 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_473 : _GEN_2631; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3166 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_474 : _GEN_2632; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3167 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_475 : _GEN_2633; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3168 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_476 : _GEN_2634; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3169 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_477 : _GEN_2635; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3170 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_478 : _GEN_2636; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3171 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_479 : _GEN_2637; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3172 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_480 : _GEN_2638; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3173 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_481 : _GEN_2639; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3174 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_482 : _GEN_2640; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3175 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_483 : _GEN_2641; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3176 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_484 : _GEN_2642; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3177 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_485 : _GEN_2643; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3178 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_486 : _GEN_2644; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3179 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_487 : _GEN_2645; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3180 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_488 : _GEN_2646; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3181 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_489 : _GEN_2647; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3182 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_490 : _GEN_2648; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3183 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_491 : _GEN_2649; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3184 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_492 : _GEN_2650; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3185 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_493 : _GEN_2651; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3186 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_494 : _GEN_2652; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3187 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_495 : _GEN_2653; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3188 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_496 : _GEN_2654; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3189 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_497 : _GEN_2655; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3190 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_498 : _GEN_2656; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3191 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_499 : _GEN_2657; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3192 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_500 : _GEN_2658; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3193 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_501 : _GEN_2659; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3194 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_502 : _GEN_2660; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3195 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_503 : _GEN_2661; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3196 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_504 : _GEN_2662; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3197 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_505 : _GEN_2663; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3198 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_506 : _GEN_2664; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3199 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_507 : _GEN_2665; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3200 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_508 : _GEN_2666; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3201 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_509 : _GEN_2667; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3202 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_510 : _GEN_2668; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_3203 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_511 : _GEN_2669; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire  mod_j = io_mod_cs == 3'h0; // @[parser_pisa.scala 56:35]
  wire  mod_j_1 = io_mod_cs == 3'h1; // @[parser_pisa.scala 56:35]
  wire  mod_j_2 = io_mod_cs == 3'h2; // @[parser_pisa.scala 56:35]
  wire  mod_j_3 = io_mod_cs == 3'h3; // @[parser_pisa.scala 56:35]
  wire  mod_j_4 = io_mod_cs == 3'h4; // @[parser_pisa.scala 56:35]
  wire  mod_j_5 = io_mod_cs == 3'h5; // @[parser_pisa.scala 56:35]
  wire  mod_j_6 = io_mod_cs == 3'h6; // @[parser_pisa.scala 56:35]
  wire  mod_j_7 = io_mod_cs == 3'h7; // @[parser_pisa.scala 56:35]
  ParseModule mau_0 ( // @[parser_pisa.scala 31:25]
    .clock(mau_0_clock),
    .io_pipe_phv_in_data_0(mau_0_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(mau_0_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(mau_0_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(mau_0_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(mau_0_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(mau_0_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(mau_0_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(mau_0_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(mau_0_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(mau_0_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(mau_0_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(mau_0_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(mau_0_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(mau_0_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(mau_0_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(mau_0_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(mau_0_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(mau_0_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(mau_0_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(mau_0_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(mau_0_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(mau_0_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(mau_0_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(mau_0_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(mau_0_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(mau_0_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(mau_0_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(mau_0_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(mau_0_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(mau_0_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(mau_0_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(mau_0_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(mau_0_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(mau_0_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(mau_0_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(mau_0_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(mau_0_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(mau_0_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(mau_0_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(mau_0_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(mau_0_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(mau_0_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(mau_0_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(mau_0_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(mau_0_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(mau_0_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(mau_0_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(mau_0_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(mau_0_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(mau_0_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(mau_0_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(mau_0_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(mau_0_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(mau_0_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(mau_0_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(mau_0_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(mau_0_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(mau_0_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(mau_0_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(mau_0_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(mau_0_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(mau_0_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(mau_0_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(mau_0_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(mau_0_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(mau_0_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(mau_0_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(mau_0_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(mau_0_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(mau_0_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(mau_0_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(mau_0_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(mau_0_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(mau_0_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(mau_0_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(mau_0_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(mau_0_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(mau_0_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(mau_0_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(mau_0_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(mau_0_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(mau_0_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(mau_0_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(mau_0_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(mau_0_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(mau_0_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(mau_0_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(mau_0_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(mau_0_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(mau_0_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(mau_0_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(mau_0_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(mau_0_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(mau_0_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(mau_0_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(mau_0_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(mau_0_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(mau_0_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(mau_0_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(mau_0_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(mau_0_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(mau_0_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(mau_0_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(mau_0_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(mau_0_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(mau_0_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(mau_0_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(mau_0_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(mau_0_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(mau_0_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(mau_0_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(mau_0_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(mau_0_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(mau_0_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(mau_0_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(mau_0_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(mau_0_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(mau_0_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(mau_0_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(mau_0_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(mau_0_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(mau_0_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(mau_0_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(mau_0_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(mau_0_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(mau_0_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(mau_0_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(mau_0_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(mau_0_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(mau_0_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(mau_0_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(mau_0_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(mau_0_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(mau_0_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(mau_0_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(mau_0_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(mau_0_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(mau_0_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(mau_0_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(mau_0_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(mau_0_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(mau_0_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(mau_0_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(mau_0_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(mau_0_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(mau_0_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(mau_0_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(mau_0_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(mau_0_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(mau_0_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(mau_0_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(mau_0_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(mau_0_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(mau_0_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(mau_0_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(mau_0_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(mau_0_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(mau_0_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(mau_0_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(mau_0_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(mau_0_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(mau_0_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(mau_0_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(mau_0_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(mau_0_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(mau_0_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(mau_0_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(mau_0_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(mau_0_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(mau_0_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(mau_0_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(mau_0_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(mau_0_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(mau_0_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(mau_0_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(mau_0_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(mau_0_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(mau_0_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(mau_0_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(mau_0_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(mau_0_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(mau_0_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(mau_0_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(mau_0_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(mau_0_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(mau_0_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(mau_0_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(mau_0_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(mau_0_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(mau_0_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(mau_0_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(mau_0_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(mau_0_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(mau_0_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(mau_0_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(mau_0_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(mau_0_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(mau_0_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(mau_0_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(mau_0_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(mau_0_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(mau_0_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(mau_0_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(mau_0_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(mau_0_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(mau_0_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(mau_0_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(mau_0_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(mau_0_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(mau_0_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(mau_0_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(mau_0_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(mau_0_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(mau_0_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(mau_0_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(mau_0_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(mau_0_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(mau_0_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(mau_0_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(mau_0_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(mau_0_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(mau_0_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(mau_0_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(mau_0_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(mau_0_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(mau_0_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(mau_0_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(mau_0_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(mau_0_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(mau_0_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(mau_0_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(mau_0_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(mau_0_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(mau_0_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(mau_0_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(mau_0_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(mau_0_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(mau_0_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(mau_0_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(mau_0_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(mau_0_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(mau_0_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(mau_0_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(mau_0_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(mau_0_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(mau_0_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(mau_0_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(mau_0_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(mau_0_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(mau_0_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(mau_0_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(mau_0_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(mau_0_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(mau_0_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(mau_0_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(mau_0_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_data_256(mau_0_io_pipe_phv_in_data_256),
    .io_pipe_phv_in_data_257(mau_0_io_pipe_phv_in_data_257),
    .io_pipe_phv_in_data_258(mau_0_io_pipe_phv_in_data_258),
    .io_pipe_phv_in_data_259(mau_0_io_pipe_phv_in_data_259),
    .io_pipe_phv_in_data_260(mau_0_io_pipe_phv_in_data_260),
    .io_pipe_phv_in_data_261(mau_0_io_pipe_phv_in_data_261),
    .io_pipe_phv_in_data_262(mau_0_io_pipe_phv_in_data_262),
    .io_pipe_phv_in_data_263(mau_0_io_pipe_phv_in_data_263),
    .io_pipe_phv_in_data_264(mau_0_io_pipe_phv_in_data_264),
    .io_pipe_phv_in_data_265(mau_0_io_pipe_phv_in_data_265),
    .io_pipe_phv_in_data_266(mau_0_io_pipe_phv_in_data_266),
    .io_pipe_phv_in_data_267(mau_0_io_pipe_phv_in_data_267),
    .io_pipe_phv_in_data_268(mau_0_io_pipe_phv_in_data_268),
    .io_pipe_phv_in_data_269(mau_0_io_pipe_phv_in_data_269),
    .io_pipe_phv_in_data_270(mau_0_io_pipe_phv_in_data_270),
    .io_pipe_phv_in_data_271(mau_0_io_pipe_phv_in_data_271),
    .io_pipe_phv_in_data_272(mau_0_io_pipe_phv_in_data_272),
    .io_pipe_phv_in_data_273(mau_0_io_pipe_phv_in_data_273),
    .io_pipe_phv_in_data_274(mau_0_io_pipe_phv_in_data_274),
    .io_pipe_phv_in_data_275(mau_0_io_pipe_phv_in_data_275),
    .io_pipe_phv_in_data_276(mau_0_io_pipe_phv_in_data_276),
    .io_pipe_phv_in_data_277(mau_0_io_pipe_phv_in_data_277),
    .io_pipe_phv_in_data_278(mau_0_io_pipe_phv_in_data_278),
    .io_pipe_phv_in_data_279(mau_0_io_pipe_phv_in_data_279),
    .io_pipe_phv_in_data_280(mau_0_io_pipe_phv_in_data_280),
    .io_pipe_phv_in_data_281(mau_0_io_pipe_phv_in_data_281),
    .io_pipe_phv_in_data_282(mau_0_io_pipe_phv_in_data_282),
    .io_pipe_phv_in_data_283(mau_0_io_pipe_phv_in_data_283),
    .io_pipe_phv_in_data_284(mau_0_io_pipe_phv_in_data_284),
    .io_pipe_phv_in_data_285(mau_0_io_pipe_phv_in_data_285),
    .io_pipe_phv_in_data_286(mau_0_io_pipe_phv_in_data_286),
    .io_pipe_phv_in_data_287(mau_0_io_pipe_phv_in_data_287),
    .io_pipe_phv_in_data_288(mau_0_io_pipe_phv_in_data_288),
    .io_pipe_phv_in_data_289(mau_0_io_pipe_phv_in_data_289),
    .io_pipe_phv_in_data_290(mau_0_io_pipe_phv_in_data_290),
    .io_pipe_phv_in_data_291(mau_0_io_pipe_phv_in_data_291),
    .io_pipe_phv_in_data_292(mau_0_io_pipe_phv_in_data_292),
    .io_pipe_phv_in_data_293(mau_0_io_pipe_phv_in_data_293),
    .io_pipe_phv_in_data_294(mau_0_io_pipe_phv_in_data_294),
    .io_pipe_phv_in_data_295(mau_0_io_pipe_phv_in_data_295),
    .io_pipe_phv_in_data_296(mau_0_io_pipe_phv_in_data_296),
    .io_pipe_phv_in_data_297(mau_0_io_pipe_phv_in_data_297),
    .io_pipe_phv_in_data_298(mau_0_io_pipe_phv_in_data_298),
    .io_pipe_phv_in_data_299(mau_0_io_pipe_phv_in_data_299),
    .io_pipe_phv_in_data_300(mau_0_io_pipe_phv_in_data_300),
    .io_pipe_phv_in_data_301(mau_0_io_pipe_phv_in_data_301),
    .io_pipe_phv_in_data_302(mau_0_io_pipe_phv_in_data_302),
    .io_pipe_phv_in_data_303(mau_0_io_pipe_phv_in_data_303),
    .io_pipe_phv_in_data_304(mau_0_io_pipe_phv_in_data_304),
    .io_pipe_phv_in_data_305(mau_0_io_pipe_phv_in_data_305),
    .io_pipe_phv_in_data_306(mau_0_io_pipe_phv_in_data_306),
    .io_pipe_phv_in_data_307(mau_0_io_pipe_phv_in_data_307),
    .io_pipe_phv_in_data_308(mau_0_io_pipe_phv_in_data_308),
    .io_pipe_phv_in_data_309(mau_0_io_pipe_phv_in_data_309),
    .io_pipe_phv_in_data_310(mau_0_io_pipe_phv_in_data_310),
    .io_pipe_phv_in_data_311(mau_0_io_pipe_phv_in_data_311),
    .io_pipe_phv_in_data_312(mau_0_io_pipe_phv_in_data_312),
    .io_pipe_phv_in_data_313(mau_0_io_pipe_phv_in_data_313),
    .io_pipe_phv_in_data_314(mau_0_io_pipe_phv_in_data_314),
    .io_pipe_phv_in_data_315(mau_0_io_pipe_phv_in_data_315),
    .io_pipe_phv_in_data_316(mau_0_io_pipe_phv_in_data_316),
    .io_pipe_phv_in_data_317(mau_0_io_pipe_phv_in_data_317),
    .io_pipe_phv_in_data_318(mau_0_io_pipe_phv_in_data_318),
    .io_pipe_phv_in_data_319(mau_0_io_pipe_phv_in_data_319),
    .io_pipe_phv_in_data_320(mau_0_io_pipe_phv_in_data_320),
    .io_pipe_phv_in_data_321(mau_0_io_pipe_phv_in_data_321),
    .io_pipe_phv_in_data_322(mau_0_io_pipe_phv_in_data_322),
    .io_pipe_phv_in_data_323(mau_0_io_pipe_phv_in_data_323),
    .io_pipe_phv_in_data_324(mau_0_io_pipe_phv_in_data_324),
    .io_pipe_phv_in_data_325(mau_0_io_pipe_phv_in_data_325),
    .io_pipe_phv_in_data_326(mau_0_io_pipe_phv_in_data_326),
    .io_pipe_phv_in_data_327(mau_0_io_pipe_phv_in_data_327),
    .io_pipe_phv_in_data_328(mau_0_io_pipe_phv_in_data_328),
    .io_pipe_phv_in_data_329(mau_0_io_pipe_phv_in_data_329),
    .io_pipe_phv_in_data_330(mau_0_io_pipe_phv_in_data_330),
    .io_pipe_phv_in_data_331(mau_0_io_pipe_phv_in_data_331),
    .io_pipe_phv_in_data_332(mau_0_io_pipe_phv_in_data_332),
    .io_pipe_phv_in_data_333(mau_0_io_pipe_phv_in_data_333),
    .io_pipe_phv_in_data_334(mau_0_io_pipe_phv_in_data_334),
    .io_pipe_phv_in_data_335(mau_0_io_pipe_phv_in_data_335),
    .io_pipe_phv_in_data_336(mau_0_io_pipe_phv_in_data_336),
    .io_pipe_phv_in_data_337(mau_0_io_pipe_phv_in_data_337),
    .io_pipe_phv_in_data_338(mau_0_io_pipe_phv_in_data_338),
    .io_pipe_phv_in_data_339(mau_0_io_pipe_phv_in_data_339),
    .io_pipe_phv_in_data_340(mau_0_io_pipe_phv_in_data_340),
    .io_pipe_phv_in_data_341(mau_0_io_pipe_phv_in_data_341),
    .io_pipe_phv_in_data_342(mau_0_io_pipe_phv_in_data_342),
    .io_pipe_phv_in_data_343(mau_0_io_pipe_phv_in_data_343),
    .io_pipe_phv_in_data_344(mau_0_io_pipe_phv_in_data_344),
    .io_pipe_phv_in_data_345(mau_0_io_pipe_phv_in_data_345),
    .io_pipe_phv_in_data_346(mau_0_io_pipe_phv_in_data_346),
    .io_pipe_phv_in_data_347(mau_0_io_pipe_phv_in_data_347),
    .io_pipe_phv_in_data_348(mau_0_io_pipe_phv_in_data_348),
    .io_pipe_phv_in_data_349(mau_0_io_pipe_phv_in_data_349),
    .io_pipe_phv_in_data_350(mau_0_io_pipe_phv_in_data_350),
    .io_pipe_phv_in_data_351(mau_0_io_pipe_phv_in_data_351),
    .io_pipe_phv_in_data_352(mau_0_io_pipe_phv_in_data_352),
    .io_pipe_phv_in_data_353(mau_0_io_pipe_phv_in_data_353),
    .io_pipe_phv_in_data_354(mau_0_io_pipe_phv_in_data_354),
    .io_pipe_phv_in_data_355(mau_0_io_pipe_phv_in_data_355),
    .io_pipe_phv_in_data_356(mau_0_io_pipe_phv_in_data_356),
    .io_pipe_phv_in_data_357(mau_0_io_pipe_phv_in_data_357),
    .io_pipe_phv_in_data_358(mau_0_io_pipe_phv_in_data_358),
    .io_pipe_phv_in_data_359(mau_0_io_pipe_phv_in_data_359),
    .io_pipe_phv_in_data_360(mau_0_io_pipe_phv_in_data_360),
    .io_pipe_phv_in_data_361(mau_0_io_pipe_phv_in_data_361),
    .io_pipe_phv_in_data_362(mau_0_io_pipe_phv_in_data_362),
    .io_pipe_phv_in_data_363(mau_0_io_pipe_phv_in_data_363),
    .io_pipe_phv_in_data_364(mau_0_io_pipe_phv_in_data_364),
    .io_pipe_phv_in_data_365(mau_0_io_pipe_phv_in_data_365),
    .io_pipe_phv_in_data_366(mau_0_io_pipe_phv_in_data_366),
    .io_pipe_phv_in_data_367(mau_0_io_pipe_phv_in_data_367),
    .io_pipe_phv_in_data_368(mau_0_io_pipe_phv_in_data_368),
    .io_pipe_phv_in_data_369(mau_0_io_pipe_phv_in_data_369),
    .io_pipe_phv_in_data_370(mau_0_io_pipe_phv_in_data_370),
    .io_pipe_phv_in_data_371(mau_0_io_pipe_phv_in_data_371),
    .io_pipe_phv_in_data_372(mau_0_io_pipe_phv_in_data_372),
    .io_pipe_phv_in_data_373(mau_0_io_pipe_phv_in_data_373),
    .io_pipe_phv_in_data_374(mau_0_io_pipe_phv_in_data_374),
    .io_pipe_phv_in_data_375(mau_0_io_pipe_phv_in_data_375),
    .io_pipe_phv_in_data_376(mau_0_io_pipe_phv_in_data_376),
    .io_pipe_phv_in_data_377(mau_0_io_pipe_phv_in_data_377),
    .io_pipe_phv_in_data_378(mau_0_io_pipe_phv_in_data_378),
    .io_pipe_phv_in_data_379(mau_0_io_pipe_phv_in_data_379),
    .io_pipe_phv_in_data_380(mau_0_io_pipe_phv_in_data_380),
    .io_pipe_phv_in_data_381(mau_0_io_pipe_phv_in_data_381),
    .io_pipe_phv_in_data_382(mau_0_io_pipe_phv_in_data_382),
    .io_pipe_phv_in_data_383(mau_0_io_pipe_phv_in_data_383),
    .io_pipe_phv_in_data_384(mau_0_io_pipe_phv_in_data_384),
    .io_pipe_phv_in_data_385(mau_0_io_pipe_phv_in_data_385),
    .io_pipe_phv_in_data_386(mau_0_io_pipe_phv_in_data_386),
    .io_pipe_phv_in_data_387(mau_0_io_pipe_phv_in_data_387),
    .io_pipe_phv_in_data_388(mau_0_io_pipe_phv_in_data_388),
    .io_pipe_phv_in_data_389(mau_0_io_pipe_phv_in_data_389),
    .io_pipe_phv_in_data_390(mau_0_io_pipe_phv_in_data_390),
    .io_pipe_phv_in_data_391(mau_0_io_pipe_phv_in_data_391),
    .io_pipe_phv_in_data_392(mau_0_io_pipe_phv_in_data_392),
    .io_pipe_phv_in_data_393(mau_0_io_pipe_phv_in_data_393),
    .io_pipe_phv_in_data_394(mau_0_io_pipe_phv_in_data_394),
    .io_pipe_phv_in_data_395(mau_0_io_pipe_phv_in_data_395),
    .io_pipe_phv_in_data_396(mau_0_io_pipe_phv_in_data_396),
    .io_pipe_phv_in_data_397(mau_0_io_pipe_phv_in_data_397),
    .io_pipe_phv_in_data_398(mau_0_io_pipe_phv_in_data_398),
    .io_pipe_phv_in_data_399(mau_0_io_pipe_phv_in_data_399),
    .io_pipe_phv_in_data_400(mau_0_io_pipe_phv_in_data_400),
    .io_pipe_phv_in_data_401(mau_0_io_pipe_phv_in_data_401),
    .io_pipe_phv_in_data_402(mau_0_io_pipe_phv_in_data_402),
    .io_pipe_phv_in_data_403(mau_0_io_pipe_phv_in_data_403),
    .io_pipe_phv_in_data_404(mau_0_io_pipe_phv_in_data_404),
    .io_pipe_phv_in_data_405(mau_0_io_pipe_phv_in_data_405),
    .io_pipe_phv_in_data_406(mau_0_io_pipe_phv_in_data_406),
    .io_pipe_phv_in_data_407(mau_0_io_pipe_phv_in_data_407),
    .io_pipe_phv_in_data_408(mau_0_io_pipe_phv_in_data_408),
    .io_pipe_phv_in_data_409(mau_0_io_pipe_phv_in_data_409),
    .io_pipe_phv_in_data_410(mau_0_io_pipe_phv_in_data_410),
    .io_pipe_phv_in_data_411(mau_0_io_pipe_phv_in_data_411),
    .io_pipe_phv_in_data_412(mau_0_io_pipe_phv_in_data_412),
    .io_pipe_phv_in_data_413(mau_0_io_pipe_phv_in_data_413),
    .io_pipe_phv_in_data_414(mau_0_io_pipe_phv_in_data_414),
    .io_pipe_phv_in_data_415(mau_0_io_pipe_phv_in_data_415),
    .io_pipe_phv_in_data_416(mau_0_io_pipe_phv_in_data_416),
    .io_pipe_phv_in_data_417(mau_0_io_pipe_phv_in_data_417),
    .io_pipe_phv_in_data_418(mau_0_io_pipe_phv_in_data_418),
    .io_pipe_phv_in_data_419(mau_0_io_pipe_phv_in_data_419),
    .io_pipe_phv_in_data_420(mau_0_io_pipe_phv_in_data_420),
    .io_pipe_phv_in_data_421(mau_0_io_pipe_phv_in_data_421),
    .io_pipe_phv_in_data_422(mau_0_io_pipe_phv_in_data_422),
    .io_pipe_phv_in_data_423(mau_0_io_pipe_phv_in_data_423),
    .io_pipe_phv_in_data_424(mau_0_io_pipe_phv_in_data_424),
    .io_pipe_phv_in_data_425(mau_0_io_pipe_phv_in_data_425),
    .io_pipe_phv_in_data_426(mau_0_io_pipe_phv_in_data_426),
    .io_pipe_phv_in_data_427(mau_0_io_pipe_phv_in_data_427),
    .io_pipe_phv_in_data_428(mau_0_io_pipe_phv_in_data_428),
    .io_pipe_phv_in_data_429(mau_0_io_pipe_phv_in_data_429),
    .io_pipe_phv_in_data_430(mau_0_io_pipe_phv_in_data_430),
    .io_pipe_phv_in_data_431(mau_0_io_pipe_phv_in_data_431),
    .io_pipe_phv_in_data_432(mau_0_io_pipe_phv_in_data_432),
    .io_pipe_phv_in_data_433(mau_0_io_pipe_phv_in_data_433),
    .io_pipe_phv_in_data_434(mau_0_io_pipe_phv_in_data_434),
    .io_pipe_phv_in_data_435(mau_0_io_pipe_phv_in_data_435),
    .io_pipe_phv_in_data_436(mau_0_io_pipe_phv_in_data_436),
    .io_pipe_phv_in_data_437(mau_0_io_pipe_phv_in_data_437),
    .io_pipe_phv_in_data_438(mau_0_io_pipe_phv_in_data_438),
    .io_pipe_phv_in_data_439(mau_0_io_pipe_phv_in_data_439),
    .io_pipe_phv_in_data_440(mau_0_io_pipe_phv_in_data_440),
    .io_pipe_phv_in_data_441(mau_0_io_pipe_phv_in_data_441),
    .io_pipe_phv_in_data_442(mau_0_io_pipe_phv_in_data_442),
    .io_pipe_phv_in_data_443(mau_0_io_pipe_phv_in_data_443),
    .io_pipe_phv_in_data_444(mau_0_io_pipe_phv_in_data_444),
    .io_pipe_phv_in_data_445(mau_0_io_pipe_phv_in_data_445),
    .io_pipe_phv_in_data_446(mau_0_io_pipe_phv_in_data_446),
    .io_pipe_phv_in_data_447(mau_0_io_pipe_phv_in_data_447),
    .io_pipe_phv_in_data_448(mau_0_io_pipe_phv_in_data_448),
    .io_pipe_phv_in_data_449(mau_0_io_pipe_phv_in_data_449),
    .io_pipe_phv_in_data_450(mau_0_io_pipe_phv_in_data_450),
    .io_pipe_phv_in_data_451(mau_0_io_pipe_phv_in_data_451),
    .io_pipe_phv_in_data_452(mau_0_io_pipe_phv_in_data_452),
    .io_pipe_phv_in_data_453(mau_0_io_pipe_phv_in_data_453),
    .io_pipe_phv_in_data_454(mau_0_io_pipe_phv_in_data_454),
    .io_pipe_phv_in_data_455(mau_0_io_pipe_phv_in_data_455),
    .io_pipe_phv_in_data_456(mau_0_io_pipe_phv_in_data_456),
    .io_pipe_phv_in_data_457(mau_0_io_pipe_phv_in_data_457),
    .io_pipe_phv_in_data_458(mau_0_io_pipe_phv_in_data_458),
    .io_pipe_phv_in_data_459(mau_0_io_pipe_phv_in_data_459),
    .io_pipe_phv_in_data_460(mau_0_io_pipe_phv_in_data_460),
    .io_pipe_phv_in_data_461(mau_0_io_pipe_phv_in_data_461),
    .io_pipe_phv_in_data_462(mau_0_io_pipe_phv_in_data_462),
    .io_pipe_phv_in_data_463(mau_0_io_pipe_phv_in_data_463),
    .io_pipe_phv_in_data_464(mau_0_io_pipe_phv_in_data_464),
    .io_pipe_phv_in_data_465(mau_0_io_pipe_phv_in_data_465),
    .io_pipe_phv_in_data_466(mau_0_io_pipe_phv_in_data_466),
    .io_pipe_phv_in_data_467(mau_0_io_pipe_phv_in_data_467),
    .io_pipe_phv_in_data_468(mau_0_io_pipe_phv_in_data_468),
    .io_pipe_phv_in_data_469(mau_0_io_pipe_phv_in_data_469),
    .io_pipe_phv_in_data_470(mau_0_io_pipe_phv_in_data_470),
    .io_pipe_phv_in_data_471(mau_0_io_pipe_phv_in_data_471),
    .io_pipe_phv_in_data_472(mau_0_io_pipe_phv_in_data_472),
    .io_pipe_phv_in_data_473(mau_0_io_pipe_phv_in_data_473),
    .io_pipe_phv_in_data_474(mau_0_io_pipe_phv_in_data_474),
    .io_pipe_phv_in_data_475(mau_0_io_pipe_phv_in_data_475),
    .io_pipe_phv_in_data_476(mau_0_io_pipe_phv_in_data_476),
    .io_pipe_phv_in_data_477(mau_0_io_pipe_phv_in_data_477),
    .io_pipe_phv_in_data_478(mau_0_io_pipe_phv_in_data_478),
    .io_pipe_phv_in_data_479(mau_0_io_pipe_phv_in_data_479),
    .io_pipe_phv_in_data_480(mau_0_io_pipe_phv_in_data_480),
    .io_pipe_phv_in_data_481(mau_0_io_pipe_phv_in_data_481),
    .io_pipe_phv_in_data_482(mau_0_io_pipe_phv_in_data_482),
    .io_pipe_phv_in_data_483(mau_0_io_pipe_phv_in_data_483),
    .io_pipe_phv_in_data_484(mau_0_io_pipe_phv_in_data_484),
    .io_pipe_phv_in_data_485(mau_0_io_pipe_phv_in_data_485),
    .io_pipe_phv_in_data_486(mau_0_io_pipe_phv_in_data_486),
    .io_pipe_phv_in_data_487(mau_0_io_pipe_phv_in_data_487),
    .io_pipe_phv_in_data_488(mau_0_io_pipe_phv_in_data_488),
    .io_pipe_phv_in_data_489(mau_0_io_pipe_phv_in_data_489),
    .io_pipe_phv_in_data_490(mau_0_io_pipe_phv_in_data_490),
    .io_pipe_phv_in_data_491(mau_0_io_pipe_phv_in_data_491),
    .io_pipe_phv_in_data_492(mau_0_io_pipe_phv_in_data_492),
    .io_pipe_phv_in_data_493(mau_0_io_pipe_phv_in_data_493),
    .io_pipe_phv_in_data_494(mau_0_io_pipe_phv_in_data_494),
    .io_pipe_phv_in_data_495(mau_0_io_pipe_phv_in_data_495),
    .io_pipe_phv_in_data_496(mau_0_io_pipe_phv_in_data_496),
    .io_pipe_phv_in_data_497(mau_0_io_pipe_phv_in_data_497),
    .io_pipe_phv_in_data_498(mau_0_io_pipe_phv_in_data_498),
    .io_pipe_phv_in_data_499(mau_0_io_pipe_phv_in_data_499),
    .io_pipe_phv_in_data_500(mau_0_io_pipe_phv_in_data_500),
    .io_pipe_phv_in_data_501(mau_0_io_pipe_phv_in_data_501),
    .io_pipe_phv_in_data_502(mau_0_io_pipe_phv_in_data_502),
    .io_pipe_phv_in_data_503(mau_0_io_pipe_phv_in_data_503),
    .io_pipe_phv_in_data_504(mau_0_io_pipe_phv_in_data_504),
    .io_pipe_phv_in_data_505(mau_0_io_pipe_phv_in_data_505),
    .io_pipe_phv_in_data_506(mau_0_io_pipe_phv_in_data_506),
    .io_pipe_phv_in_data_507(mau_0_io_pipe_phv_in_data_507),
    .io_pipe_phv_in_data_508(mau_0_io_pipe_phv_in_data_508),
    .io_pipe_phv_in_data_509(mau_0_io_pipe_phv_in_data_509),
    .io_pipe_phv_in_data_510(mau_0_io_pipe_phv_in_data_510),
    .io_pipe_phv_in_data_511(mau_0_io_pipe_phv_in_data_511),
    .io_pipe_phv_in_header_0(mau_0_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(mau_0_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(mau_0_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(mau_0_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(mau_0_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(mau_0_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(mau_0_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(mau_0_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(mau_0_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(mau_0_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(mau_0_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(mau_0_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(mau_0_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(mau_0_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(mau_0_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(mau_0_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(mau_0_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(mau_0_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(mau_0_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(mau_0_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(mau_0_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(mau_0_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(mau_0_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(mau_0_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(mau_0_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(mau_0_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(mau_0_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(mau_0_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(mau_0_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(mau_0_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(mau_0_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(mau_0_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(mau_0_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(mau_0_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(mau_0_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(mau_0_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(mau_0_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(mau_0_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(mau_0_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(mau_0_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(mau_0_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(mau_0_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(mau_0_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(mau_0_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(mau_0_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(mau_0_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(mau_0_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(mau_0_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(mau_0_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(mau_0_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(mau_0_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(mau_0_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(mau_0_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(mau_0_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(mau_0_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(mau_0_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(mau_0_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(mau_0_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(mau_0_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(mau_0_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(mau_0_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(mau_0_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(mau_0_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(mau_0_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(mau_0_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(mau_0_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(mau_0_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(mau_0_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(mau_0_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(mau_0_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(mau_0_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(mau_0_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(mau_0_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(mau_0_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(mau_0_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(mau_0_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(mau_0_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(mau_0_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(mau_0_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(mau_0_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(mau_0_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(mau_0_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(mau_0_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(mau_0_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(mau_0_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(mau_0_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(mau_0_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(mau_0_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(mau_0_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(mau_0_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(mau_0_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(mau_0_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(mau_0_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(mau_0_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(mau_0_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(mau_0_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(mau_0_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(mau_0_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(mau_0_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(mau_0_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(mau_0_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(mau_0_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(mau_0_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(mau_0_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(mau_0_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(mau_0_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(mau_0_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(mau_0_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(mau_0_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(mau_0_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(mau_0_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(mau_0_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(mau_0_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(mau_0_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(mau_0_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(mau_0_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(mau_0_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(mau_0_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(mau_0_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(mau_0_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(mau_0_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(mau_0_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(mau_0_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(mau_0_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(mau_0_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(mau_0_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(mau_0_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(mau_0_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(mau_0_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(mau_0_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(mau_0_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(mau_0_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(mau_0_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(mau_0_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(mau_0_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(mau_0_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(mau_0_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(mau_0_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(mau_0_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(mau_0_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(mau_0_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(mau_0_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(mau_0_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(mau_0_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(mau_0_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(mau_0_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(mau_0_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(mau_0_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(mau_0_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(mau_0_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(mau_0_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(mau_0_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(mau_0_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(mau_0_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(mau_0_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(mau_0_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(mau_0_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(mau_0_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(mau_0_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(mau_0_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(mau_0_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(mau_0_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(mau_0_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(mau_0_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(mau_0_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(mau_0_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(mau_0_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(mau_0_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(mau_0_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(mau_0_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(mau_0_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(mau_0_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(mau_0_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(mau_0_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(mau_0_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(mau_0_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(mau_0_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(mau_0_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(mau_0_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(mau_0_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(mau_0_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(mau_0_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(mau_0_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(mau_0_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(mau_0_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(mau_0_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(mau_0_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(mau_0_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(mau_0_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(mau_0_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(mau_0_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(mau_0_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(mau_0_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(mau_0_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(mau_0_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(mau_0_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(mau_0_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(mau_0_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(mau_0_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(mau_0_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(mau_0_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(mau_0_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(mau_0_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(mau_0_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(mau_0_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(mau_0_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(mau_0_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(mau_0_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(mau_0_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(mau_0_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(mau_0_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(mau_0_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(mau_0_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(mau_0_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(mau_0_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(mau_0_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(mau_0_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(mau_0_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(mau_0_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(mau_0_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(mau_0_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(mau_0_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(mau_0_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(mau_0_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(mau_0_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(mau_0_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(mau_0_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(mau_0_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(mau_0_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(mau_0_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(mau_0_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(mau_0_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(mau_0_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(mau_0_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(mau_0_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(mau_0_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(mau_0_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(mau_0_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(mau_0_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(mau_0_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(mau_0_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(mau_0_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(mau_0_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(mau_0_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(mau_0_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(mau_0_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(mau_0_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(mau_0_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(mau_0_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(mau_0_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(mau_0_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(mau_0_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(mau_0_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(mau_0_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(mau_0_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(mau_0_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(mau_0_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(mau_0_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(mau_0_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(mau_0_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(mau_0_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(mau_0_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(mau_0_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(mau_0_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(mau_0_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(mau_0_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(mau_0_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(mau_0_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(mau_0_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(mau_0_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(mau_0_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(mau_0_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(mau_0_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(mau_0_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(mau_0_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(mau_0_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(mau_0_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(mau_0_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_data_256(mau_0_io_pipe_phv_out_data_256),
    .io_pipe_phv_out_data_257(mau_0_io_pipe_phv_out_data_257),
    .io_pipe_phv_out_data_258(mau_0_io_pipe_phv_out_data_258),
    .io_pipe_phv_out_data_259(mau_0_io_pipe_phv_out_data_259),
    .io_pipe_phv_out_data_260(mau_0_io_pipe_phv_out_data_260),
    .io_pipe_phv_out_data_261(mau_0_io_pipe_phv_out_data_261),
    .io_pipe_phv_out_data_262(mau_0_io_pipe_phv_out_data_262),
    .io_pipe_phv_out_data_263(mau_0_io_pipe_phv_out_data_263),
    .io_pipe_phv_out_data_264(mau_0_io_pipe_phv_out_data_264),
    .io_pipe_phv_out_data_265(mau_0_io_pipe_phv_out_data_265),
    .io_pipe_phv_out_data_266(mau_0_io_pipe_phv_out_data_266),
    .io_pipe_phv_out_data_267(mau_0_io_pipe_phv_out_data_267),
    .io_pipe_phv_out_data_268(mau_0_io_pipe_phv_out_data_268),
    .io_pipe_phv_out_data_269(mau_0_io_pipe_phv_out_data_269),
    .io_pipe_phv_out_data_270(mau_0_io_pipe_phv_out_data_270),
    .io_pipe_phv_out_data_271(mau_0_io_pipe_phv_out_data_271),
    .io_pipe_phv_out_data_272(mau_0_io_pipe_phv_out_data_272),
    .io_pipe_phv_out_data_273(mau_0_io_pipe_phv_out_data_273),
    .io_pipe_phv_out_data_274(mau_0_io_pipe_phv_out_data_274),
    .io_pipe_phv_out_data_275(mau_0_io_pipe_phv_out_data_275),
    .io_pipe_phv_out_data_276(mau_0_io_pipe_phv_out_data_276),
    .io_pipe_phv_out_data_277(mau_0_io_pipe_phv_out_data_277),
    .io_pipe_phv_out_data_278(mau_0_io_pipe_phv_out_data_278),
    .io_pipe_phv_out_data_279(mau_0_io_pipe_phv_out_data_279),
    .io_pipe_phv_out_data_280(mau_0_io_pipe_phv_out_data_280),
    .io_pipe_phv_out_data_281(mau_0_io_pipe_phv_out_data_281),
    .io_pipe_phv_out_data_282(mau_0_io_pipe_phv_out_data_282),
    .io_pipe_phv_out_data_283(mau_0_io_pipe_phv_out_data_283),
    .io_pipe_phv_out_data_284(mau_0_io_pipe_phv_out_data_284),
    .io_pipe_phv_out_data_285(mau_0_io_pipe_phv_out_data_285),
    .io_pipe_phv_out_data_286(mau_0_io_pipe_phv_out_data_286),
    .io_pipe_phv_out_data_287(mau_0_io_pipe_phv_out_data_287),
    .io_pipe_phv_out_data_288(mau_0_io_pipe_phv_out_data_288),
    .io_pipe_phv_out_data_289(mau_0_io_pipe_phv_out_data_289),
    .io_pipe_phv_out_data_290(mau_0_io_pipe_phv_out_data_290),
    .io_pipe_phv_out_data_291(mau_0_io_pipe_phv_out_data_291),
    .io_pipe_phv_out_data_292(mau_0_io_pipe_phv_out_data_292),
    .io_pipe_phv_out_data_293(mau_0_io_pipe_phv_out_data_293),
    .io_pipe_phv_out_data_294(mau_0_io_pipe_phv_out_data_294),
    .io_pipe_phv_out_data_295(mau_0_io_pipe_phv_out_data_295),
    .io_pipe_phv_out_data_296(mau_0_io_pipe_phv_out_data_296),
    .io_pipe_phv_out_data_297(mau_0_io_pipe_phv_out_data_297),
    .io_pipe_phv_out_data_298(mau_0_io_pipe_phv_out_data_298),
    .io_pipe_phv_out_data_299(mau_0_io_pipe_phv_out_data_299),
    .io_pipe_phv_out_data_300(mau_0_io_pipe_phv_out_data_300),
    .io_pipe_phv_out_data_301(mau_0_io_pipe_phv_out_data_301),
    .io_pipe_phv_out_data_302(mau_0_io_pipe_phv_out_data_302),
    .io_pipe_phv_out_data_303(mau_0_io_pipe_phv_out_data_303),
    .io_pipe_phv_out_data_304(mau_0_io_pipe_phv_out_data_304),
    .io_pipe_phv_out_data_305(mau_0_io_pipe_phv_out_data_305),
    .io_pipe_phv_out_data_306(mau_0_io_pipe_phv_out_data_306),
    .io_pipe_phv_out_data_307(mau_0_io_pipe_phv_out_data_307),
    .io_pipe_phv_out_data_308(mau_0_io_pipe_phv_out_data_308),
    .io_pipe_phv_out_data_309(mau_0_io_pipe_phv_out_data_309),
    .io_pipe_phv_out_data_310(mau_0_io_pipe_phv_out_data_310),
    .io_pipe_phv_out_data_311(mau_0_io_pipe_phv_out_data_311),
    .io_pipe_phv_out_data_312(mau_0_io_pipe_phv_out_data_312),
    .io_pipe_phv_out_data_313(mau_0_io_pipe_phv_out_data_313),
    .io_pipe_phv_out_data_314(mau_0_io_pipe_phv_out_data_314),
    .io_pipe_phv_out_data_315(mau_0_io_pipe_phv_out_data_315),
    .io_pipe_phv_out_data_316(mau_0_io_pipe_phv_out_data_316),
    .io_pipe_phv_out_data_317(mau_0_io_pipe_phv_out_data_317),
    .io_pipe_phv_out_data_318(mau_0_io_pipe_phv_out_data_318),
    .io_pipe_phv_out_data_319(mau_0_io_pipe_phv_out_data_319),
    .io_pipe_phv_out_data_320(mau_0_io_pipe_phv_out_data_320),
    .io_pipe_phv_out_data_321(mau_0_io_pipe_phv_out_data_321),
    .io_pipe_phv_out_data_322(mau_0_io_pipe_phv_out_data_322),
    .io_pipe_phv_out_data_323(mau_0_io_pipe_phv_out_data_323),
    .io_pipe_phv_out_data_324(mau_0_io_pipe_phv_out_data_324),
    .io_pipe_phv_out_data_325(mau_0_io_pipe_phv_out_data_325),
    .io_pipe_phv_out_data_326(mau_0_io_pipe_phv_out_data_326),
    .io_pipe_phv_out_data_327(mau_0_io_pipe_phv_out_data_327),
    .io_pipe_phv_out_data_328(mau_0_io_pipe_phv_out_data_328),
    .io_pipe_phv_out_data_329(mau_0_io_pipe_phv_out_data_329),
    .io_pipe_phv_out_data_330(mau_0_io_pipe_phv_out_data_330),
    .io_pipe_phv_out_data_331(mau_0_io_pipe_phv_out_data_331),
    .io_pipe_phv_out_data_332(mau_0_io_pipe_phv_out_data_332),
    .io_pipe_phv_out_data_333(mau_0_io_pipe_phv_out_data_333),
    .io_pipe_phv_out_data_334(mau_0_io_pipe_phv_out_data_334),
    .io_pipe_phv_out_data_335(mau_0_io_pipe_phv_out_data_335),
    .io_pipe_phv_out_data_336(mau_0_io_pipe_phv_out_data_336),
    .io_pipe_phv_out_data_337(mau_0_io_pipe_phv_out_data_337),
    .io_pipe_phv_out_data_338(mau_0_io_pipe_phv_out_data_338),
    .io_pipe_phv_out_data_339(mau_0_io_pipe_phv_out_data_339),
    .io_pipe_phv_out_data_340(mau_0_io_pipe_phv_out_data_340),
    .io_pipe_phv_out_data_341(mau_0_io_pipe_phv_out_data_341),
    .io_pipe_phv_out_data_342(mau_0_io_pipe_phv_out_data_342),
    .io_pipe_phv_out_data_343(mau_0_io_pipe_phv_out_data_343),
    .io_pipe_phv_out_data_344(mau_0_io_pipe_phv_out_data_344),
    .io_pipe_phv_out_data_345(mau_0_io_pipe_phv_out_data_345),
    .io_pipe_phv_out_data_346(mau_0_io_pipe_phv_out_data_346),
    .io_pipe_phv_out_data_347(mau_0_io_pipe_phv_out_data_347),
    .io_pipe_phv_out_data_348(mau_0_io_pipe_phv_out_data_348),
    .io_pipe_phv_out_data_349(mau_0_io_pipe_phv_out_data_349),
    .io_pipe_phv_out_data_350(mau_0_io_pipe_phv_out_data_350),
    .io_pipe_phv_out_data_351(mau_0_io_pipe_phv_out_data_351),
    .io_pipe_phv_out_data_352(mau_0_io_pipe_phv_out_data_352),
    .io_pipe_phv_out_data_353(mau_0_io_pipe_phv_out_data_353),
    .io_pipe_phv_out_data_354(mau_0_io_pipe_phv_out_data_354),
    .io_pipe_phv_out_data_355(mau_0_io_pipe_phv_out_data_355),
    .io_pipe_phv_out_data_356(mau_0_io_pipe_phv_out_data_356),
    .io_pipe_phv_out_data_357(mau_0_io_pipe_phv_out_data_357),
    .io_pipe_phv_out_data_358(mau_0_io_pipe_phv_out_data_358),
    .io_pipe_phv_out_data_359(mau_0_io_pipe_phv_out_data_359),
    .io_pipe_phv_out_data_360(mau_0_io_pipe_phv_out_data_360),
    .io_pipe_phv_out_data_361(mau_0_io_pipe_phv_out_data_361),
    .io_pipe_phv_out_data_362(mau_0_io_pipe_phv_out_data_362),
    .io_pipe_phv_out_data_363(mau_0_io_pipe_phv_out_data_363),
    .io_pipe_phv_out_data_364(mau_0_io_pipe_phv_out_data_364),
    .io_pipe_phv_out_data_365(mau_0_io_pipe_phv_out_data_365),
    .io_pipe_phv_out_data_366(mau_0_io_pipe_phv_out_data_366),
    .io_pipe_phv_out_data_367(mau_0_io_pipe_phv_out_data_367),
    .io_pipe_phv_out_data_368(mau_0_io_pipe_phv_out_data_368),
    .io_pipe_phv_out_data_369(mau_0_io_pipe_phv_out_data_369),
    .io_pipe_phv_out_data_370(mau_0_io_pipe_phv_out_data_370),
    .io_pipe_phv_out_data_371(mau_0_io_pipe_phv_out_data_371),
    .io_pipe_phv_out_data_372(mau_0_io_pipe_phv_out_data_372),
    .io_pipe_phv_out_data_373(mau_0_io_pipe_phv_out_data_373),
    .io_pipe_phv_out_data_374(mau_0_io_pipe_phv_out_data_374),
    .io_pipe_phv_out_data_375(mau_0_io_pipe_phv_out_data_375),
    .io_pipe_phv_out_data_376(mau_0_io_pipe_phv_out_data_376),
    .io_pipe_phv_out_data_377(mau_0_io_pipe_phv_out_data_377),
    .io_pipe_phv_out_data_378(mau_0_io_pipe_phv_out_data_378),
    .io_pipe_phv_out_data_379(mau_0_io_pipe_phv_out_data_379),
    .io_pipe_phv_out_data_380(mau_0_io_pipe_phv_out_data_380),
    .io_pipe_phv_out_data_381(mau_0_io_pipe_phv_out_data_381),
    .io_pipe_phv_out_data_382(mau_0_io_pipe_phv_out_data_382),
    .io_pipe_phv_out_data_383(mau_0_io_pipe_phv_out_data_383),
    .io_pipe_phv_out_data_384(mau_0_io_pipe_phv_out_data_384),
    .io_pipe_phv_out_data_385(mau_0_io_pipe_phv_out_data_385),
    .io_pipe_phv_out_data_386(mau_0_io_pipe_phv_out_data_386),
    .io_pipe_phv_out_data_387(mau_0_io_pipe_phv_out_data_387),
    .io_pipe_phv_out_data_388(mau_0_io_pipe_phv_out_data_388),
    .io_pipe_phv_out_data_389(mau_0_io_pipe_phv_out_data_389),
    .io_pipe_phv_out_data_390(mau_0_io_pipe_phv_out_data_390),
    .io_pipe_phv_out_data_391(mau_0_io_pipe_phv_out_data_391),
    .io_pipe_phv_out_data_392(mau_0_io_pipe_phv_out_data_392),
    .io_pipe_phv_out_data_393(mau_0_io_pipe_phv_out_data_393),
    .io_pipe_phv_out_data_394(mau_0_io_pipe_phv_out_data_394),
    .io_pipe_phv_out_data_395(mau_0_io_pipe_phv_out_data_395),
    .io_pipe_phv_out_data_396(mau_0_io_pipe_phv_out_data_396),
    .io_pipe_phv_out_data_397(mau_0_io_pipe_phv_out_data_397),
    .io_pipe_phv_out_data_398(mau_0_io_pipe_phv_out_data_398),
    .io_pipe_phv_out_data_399(mau_0_io_pipe_phv_out_data_399),
    .io_pipe_phv_out_data_400(mau_0_io_pipe_phv_out_data_400),
    .io_pipe_phv_out_data_401(mau_0_io_pipe_phv_out_data_401),
    .io_pipe_phv_out_data_402(mau_0_io_pipe_phv_out_data_402),
    .io_pipe_phv_out_data_403(mau_0_io_pipe_phv_out_data_403),
    .io_pipe_phv_out_data_404(mau_0_io_pipe_phv_out_data_404),
    .io_pipe_phv_out_data_405(mau_0_io_pipe_phv_out_data_405),
    .io_pipe_phv_out_data_406(mau_0_io_pipe_phv_out_data_406),
    .io_pipe_phv_out_data_407(mau_0_io_pipe_phv_out_data_407),
    .io_pipe_phv_out_data_408(mau_0_io_pipe_phv_out_data_408),
    .io_pipe_phv_out_data_409(mau_0_io_pipe_phv_out_data_409),
    .io_pipe_phv_out_data_410(mau_0_io_pipe_phv_out_data_410),
    .io_pipe_phv_out_data_411(mau_0_io_pipe_phv_out_data_411),
    .io_pipe_phv_out_data_412(mau_0_io_pipe_phv_out_data_412),
    .io_pipe_phv_out_data_413(mau_0_io_pipe_phv_out_data_413),
    .io_pipe_phv_out_data_414(mau_0_io_pipe_phv_out_data_414),
    .io_pipe_phv_out_data_415(mau_0_io_pipe_phv_out_data_415),
    .io_pipe_phv_out_data_416(mau_0_io_pipe_phv_out_data_416),
    .io_pipe_phv_out_data_417(mau_0_io_pipe_phv_out_data_417),
    .io_pipe_phv_out_data_418(mau_0_io_pipe_phv_out_data_418),
    .io_pipe_phv_out_data_419(mau_0_io_pipe_phv_out_data_419),
    .io_pipe_phv_out_data_420(mau_0_io_pipe_phv_out_data_420),
    .io_pipe_phv_out_data_421(mau_0_io_pipe_phv_out_data_421),
    .io_pipe_phv_out_data_422(mau_0_io_pipe_phv_out_data_422),
    .io_pipe_phv_out_data_423(mau_0_io_pipe_phv_out_data_423),
    .io_pipe_phv_out_data_424(mau_0_io_pipe_phv_out_data_424),
    .io_pipe_phv_out_data_425(mau_0_io_pipe_phv_out_data_425),
    .io_pipe_phv_out_data_426(mau_0_io_pipe_phv_out_data_426),
    .io_pipe_phv_out_data_427(mau_0_io_pipe_phv_out_data_427),
    .io_pipe_phv_out_data_428(mau_0_io_pipe_phv_out_data_428),
    .io_pipe_phv_out_data_429(mau_0_io_pipe_phv_out_data_429),
    .io_pipe_phv_out_data_430(mau_0_io_pipe_phv_out_data_430),
    .io_pipe_phv_out_data_431(mau_0_io_pipe_phv_out_data_431),
    .io_pipe_phv_out_data_432(mau_0_io_pipe_phv_out_data_432),
    .io_pipe_phv_out_data_433(mau_0_io_pipe_phv_out_data_433),
    .io_pipe_phv_out_data_434(mau_0_io_pipe_phv_out_data_434),
    .io_pipe_phv_out_data_435(mau_0_io_pipe_phv_out_data_435),
    .io_pipe_phv_out_data_436(mau_0_io_pipe_phv_out_data_436),
    .io_pipe_phv_out_data_437(mau_0_io_pipe_phv_out_data_437),
    .io_pipe_phv_out_data_438(mau_0_io_pipe_phv_out_data_438),
    .io_pipe_phv_out_data_439(mau_0_io_pipe_phv_out_data_439),
    .io_pipe_phv_out_data_440(mau_0_io_pipe_phv_out_data_440),
    .io_pipe_phv_out_data_441(mau_0_io_pipe_phv_out_data_441),
    .io_pipe_phv_out_data_442(mau_0_io_pipe_phv_out_data_442),
    .io_pipe_phv_out_data_443(mau_0_io_pipe_phv_out_data_443),
    .io_pipe_phv_out_data_444(mau_0_io_pipe_phv_out_data_444),
    .io_pipe_phv_out_data_445(mau_0_io_pipe_phv_out_data_445),
    .io_pipe_phv_out_data_446(mau_0_io_pipe_phv_out_data_446),
    .io_pipe_phv_out_data_447(mau_0_io_pipe_phv_out_data_447),
    .io_pipe_phv_out_data_448(mau_0_io_pipe_phv_out_data_448),
    .io_pipe_phv_out_data_449(mau_0_io_pipe_phv_out_data_449),
    .io_pipe_phv_out_data_450(mau_0_io_pipe_phv_out_data_450),
    .io_pipe_phv_out_data_451(mau_0_io_pipe_phv_out_data_451),
    .io_pipe_phv_out_data_452(mau_0_io_pipe_phv_out_data_452),
    .io_pipe_phv_out_data_453(mau_0_io_pipe_phv_out_data_453),
    .io_pipe_phv_out_data_454(mau_0_io_pipe_phv_out_data_454),
    .io_pipe_phv_out_data_455(mau_0_io_pipe_phv_out_data_455),
    .io_pipe_phv_out_data_456(mau_0_io_pipe_phv_out_data_456),
    .io_pipe_phv_out_data_457(mau_0_io_pipe_phv_out_data_457),
    .io_pipe_phv_out_data_458(mau_0_io_pipe_phv_out_data_458),
    .io_pipe_phv_out_data_459(mau_0_io_pipe_phv_out_data_459),
    .io_pipe_phv_out_data_460(mau_0_io_pipe_phv_out_data_460),
    .io_pipe_phv_out_data_461(mau_0_io_pipe_phv_out_data_461),
    .io_pipe_phv_out_data_462(mau_0_io_pipe_phv_out_data_462),
    .io_pipe_phv_out_data_463(mau_0_io_pipe_phv_out_data_463),
    .io_pipe_phv_out_data_464(mau_0_io_pipe_phv_out_data_464),
    .io_pipe_phv_out_data_465(mau_0_io_pipe_phv_out_data_465),
    .io_pipe_phv_out_data_466(mau_0_io_pipe_phv_out_data_466),
    .io_pipe_phv_out_data_467(mau_0_io_pipe_phv_out_data_467),
    .io_pipe_phv_out_data_468(mau_0_io_pipe_phv_out_data_468),
    .io_pipe_phv_out_data_469(mau_0_io_pipe_phv_out_data_469),
    .io_pipe_phv_out_data_470(mau_0_io_pipe_phv_out_data_470),
    .io_pipe_phv_out_data_471(mau_0_io_pipe_phv_out_data_471),
    .io_pipe_phv_out_data_472(mau_0_io_pipe_phv_out_data_472),
    .io_pipe_phv_out_data_473(mau_0_io_pipe_phv_out_data_473),
    .io_pipe_phv_out_data_474(mau_0_io_pipe_phv_out_data_474),
    .io_pipe_phv_out_data_475(mau_0_io_pipe_phv_out_data_475),
    .io_pipe_phv_out_data_476(mau_0_io_pipe_phv_out_data_476),
    .io_pipe_phv_out_data_477(mau_0_io_pipe_phv_out_data_477),
    .io_pipe_phv_out_data_478(mau_0_io_pipe_phv_out_data_478),
    .io_pipe_phv_out_data_479(mau_0_io_pipe_phv_out_data_479),
    .io_pipe_phv_out_data_480(mau_0_io_pipe_phv_out_data_480),
    .io_pipe_phv_out_data_481(mau_0_io_pipe_phv_out_data_481),
    .io_pipe_phv_out_data_482(mau_0_io_pipe_phv_out_data_482),
    .io_pipe_phv_out_data_483(mau_0_io_pipe_phv_out_data_483),
    .io_pipe_phv_out_data_484(mau_0_io_pipe_phv_out_data_484),
    .io_pipe_phv_out_data_485(mau_0_io_pipe_phv_out_data_485),
    .io_pipe_phv_out_data_486(mau_0_io_pipe_phv_out_data_486),
    .io_pipe_phv_out_data_487(mau_0_io_pipe_phv_out_data_487),
    .io_pipe_phv_out_data_488(mau_0_io_pipe_phv_out_data_488),
    .io_pipe_phv_out_data_489(mau_0_io_pipe_phv_out_data_489),
    .io_pipe_phv_out_data_490(mau_0_io_pipe_phv_out_data_490),
    .io_pipe_phv_out_data_491(mau_0_io_pipe_phv_out_data_491),
    .io_pipe_phv_out_data_492(mau_0_io_pipe_phv_out_data_492),
    .io_pipe_phv_out_data_493(mau_0_io_pipe_phv_out_data_493),
    .io_pipe_phv_out_data_494(mau_0_io_pipe_phv_out_data_494),
    .io_pipe_phv_out_data_495(mau_0_io_pipe_phv_out_data_495),
    .io_pipe_phv_out_data_496(mau_0_io_pipe_phv_out_data_496),
    .io_pipe_phv_out_data_497(mau_0_io_pipe_phv_out_data_497),
    .io_pipe_phv_out_data_498(mau_0_io_pipe_phv_out_data_498),
    .io_pipe_phv_out_data_499(mau_0_io_pipe_phv_out_data_499),
    .io_pipe_phv_out_data_500(mau_0_io_pipe_phv_out_data_500),
    .io_pipe_phv_out_data_501(mau_0_io_pipe_phv_out_data_501),
    .io_pipe_phv_out_data_502(mau_0_io_pipe_phv_out_data_502),
    .io_pipe_phv_out_data_503(mau_0_io_pipe_phv_out_data_503),
    .io_pipe_phv_out_data_504(mau_0_io_pipe_phv_out_data_504),
    .io_pipe_phv_out_data_505(mau_0_io_pipe_phv_out_data_505),
    .io_pipe_phv_out_data_506(mau_0_io_pipe_phv_out_data_506),
    .io_pipe_phv_out_data_507(mau_0_io_pipe_phv_out_data_507),
    .io_pipe_phv_out_data_508(mau_0_io_pipe_phv_out_data_508),
    .io_pipe_phv_out_data_509(mau_0_io_pipe_phv_out_data_509),
    .io_pipe_phv_out_data_510(mau_0_io_pipe_phv_out_data_510),
    .io_pipe_phv_out_data_511(mau_0_io_pipe_phv_out_data_511),
    .io_pipe_phv_out_header_0(mau_0_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(mau_0_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(mau_0_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(mau_0_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(mau_0_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(mau_0_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(mau_0_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(mau_0_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(mau_0_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(mau_0_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(mau_0_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(mau_0_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(mau_0_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(mau_0_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(mau_0_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(mau_0_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(mau_0_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(mau_0_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(mau_0_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(mau_0_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(mau_0_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(mau_0_io_pipe_phv_out_is_valid_processor),
    .io_mod_state_id_mod(mau_0_io_mod_state_id_mod),
    .io_mod_state_id(mau_0_io_mod_state_id),
    .io_mod_sram_w_cs(mau_0_io_mod_sram_w_cs),
    .io_mod_sram_w_en(mau_0_io_mod_sram_w_en),
    .io_mod_sram_w_addr(mau_0_io_mod_sram_w_addr),
    .io_mod_sram_w_data(mau_0_io_mod_sram_w_data)
  );
  ParseModule mau_1 ( // @[parser_pisa.scala 31:25]
    .clock(mau_1_clock),
    .io_pipe_phv_in_data_0(mau_1_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(mau_1_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(mau_1_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(mau_1_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(mau_1_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(mau_1_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(mau_1_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(mau_1_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(mau_1_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(mau_1_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(mau_1_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(mau_1_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(mau_1_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(mau_1_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(mau_1_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(mau_1_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(mau_1_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(mau_1_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(mau_1_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(mau_1_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(mau_1_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(mau_1_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(mau_1_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(mau_1_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(mau_1_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(mau_1_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(mau_1_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(mau_1_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(mau_1_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(mau_1_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(mau_1_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(mau_1_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(mau_1_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(mau_1_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(mau_1_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(mau_1_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(mau_1_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(mau_1_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(mau_1_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(mau_1_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(mau_1_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(mau_1_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(mau_1_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(mau_1_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(mau_1_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(mau_1_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(mau_1_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(mau_1_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(mau_1_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(mau_1_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(mau_1_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(mau_1_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(mau_1_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(mau_1_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(mau_1_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(mau_1_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(mau_1_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(mau_1_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(mau_1_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(mau_1_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(mau_1_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(mau_1_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(mau_1_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(mau_1_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(mau_1_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(mau_1_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(mau_1_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(mau_1_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(mau_1_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(mau_1_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(mau_1_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(mau_1_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(mau_1_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(mau_1_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(mau_1_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(mau_1_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(mau_1_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(mau_1_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(mau_1_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(mau_1_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(mau_1_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(mau_1_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(mau_1_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(mau_1_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(mau_1_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(mau_1_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(mau_1_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(mau_1_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(mau_1_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(mau_1_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(mau_1_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(mau_1_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(mau_1_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(mau_1_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(mau_1_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(mau_1_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(mau_1_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(mau_1_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(mau_1_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(mau_1_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(mau_1_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(mau_1_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(mau_1_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(mau_1_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(mau_1_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(mau_1_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(mau_1_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(mau_1_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(mau_1_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(mau_1_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(mau_1_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(mau_1_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(mau_1_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(mau_1_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(mau_1_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(mau_1_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(mau_1_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(mau_1_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(mau_1_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(mau_1_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(mau_1_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(mau_1_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(mau_1_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(mau_1_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(mau_1_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(mau_1_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(mau_1_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(mau_1_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(mau_1_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(mau_1_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(mau_1_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(mau_1_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(mau_1_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(mau_1_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(mau_1_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(mau_1_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(mau_1_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(mau_1_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(mau_1_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(mau_1_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(mau_1_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(mau_1_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(mau_1_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(mau_1_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(mau_1_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(mau_1_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(mau_1_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(mau_1_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(mau_1_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(mau_1_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(mau_1_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(mau_1_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(mau_1_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(mau_1_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(mau_1_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(mau_1_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(mau_1_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(mau_1_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(mau_1_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(mau_1_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(mau_1_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(mau_1_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(mau_1_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(mau_1_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(mau_1_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(mau_1_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(mau_1_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(mau_1_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(mau_1_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(mau_1_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(mau_1_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(mau_1_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(mau_1_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(mau_1_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(mau_1_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(mau_1_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(mau_1_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(mau_1_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(mau_1_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(mau_1_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(mau_1_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(mau_1_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(mau_1_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(mau_1_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(mau_1_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(mau_1_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(mau_1_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(mau_1_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(mau_1_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(mau_1_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(mau_1_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(mau_1_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(mau_1_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(mau_1_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(mau_1_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(mau_1_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(mau_1_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(mau_1_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(mau_1_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(mau_1_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(mau_1_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(mau_1_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(mau_1_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(mau_1_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(mau_1_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(mau_1_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(mau_1_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(mau_1_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(mau_1_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(mau_1_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(mau_1_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(mau_1_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(mau_1_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(mau_1_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(mau_1_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(mau_1_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(mau_1_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(mau_1_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(mau_1_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(mau_1_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(mau_1_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(mau_1_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(mau_1_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(mau_1_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(mau_1_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(mau_1_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(mau_1_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(mau_1_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(mau_1_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(mau_1_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(mau_1_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(mau_1_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(mau_1_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(mau_1_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(mau_1_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(mau_1_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(mau_1_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(mau_1_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(mau_1_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(mau_1_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(mau_1_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(mau_1_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(mau_1_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(mau_1_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(mau_1_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(mau_1_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(mau_1_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(mau_1_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(mau_1_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(mau_1_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(mau_1_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(mau_1_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(mau_1_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(mau_1_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(mau_1_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(mau_1_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_data_256(mau_1_io_pipe_phv_in_data_256),
    .io_pipe_phv_in_data_257(mau_1_io_pipe_phv_in_data_257),
    .io_pipe_phv_in_data_258(mau_1_io_pipe_phv_in_data_258),
    .io_pipe_phv_in_data_259(mau_1_io_pipe_phv_in_data_259),
    .io_pipe_phv_in_data_260(mau_1_io_pipe_phv_in_data_260),
    .io_pipe_phv_in_data_261(mau_1_io_pipe_phv_in_data_261),
    .io_pipe_phv_in_data_262(mau_1_io_pipe_phv_in_data_262),
    .io_pipe_phv_in_data_263(mau_1_io_pipe_phv_in_data_263),
    .io_pipe_phv_in_data_264(mau_1_io_pipe_phv_in_data_264),
    .io_pipe_phv_in_data_265(mau_1_io_pipe_phv_in_data_265),
    .io_pipe_phv_in_data_266(mau_1_io_pipe_phv_in_data_266),
    .io_pipe_phv_in_data_267(mau_1_io_pipe_phv_in_data_267),
    .io_pipe_phv_in_data_268(mau_1_io_pipe_phv_in_data_268),
    .io_pipe_phv_in_data_269(mau_1_io_pipe_phv_in_data_269),
    .io_pipe_phv_in_data_270(mau_1_io_pipe_phv_in_data_270),
    .io_pipe_phv_in_data_271(mau_1_io_pipe_phv_in_data_271),
    .io_pipe_phv_in_data_272(mau_1_io_pipe_phv_in_data_272),
    .io_pipe_phv_in_data_273(mau_1_io_pipe_phv_in_data_273),
    .io_pipe_phv_in_data_274(mau_1_io_pipe_phv_in_data_274),
    .io_pipe_phv_in_data_275(mau_1_io_pipe_phv_in_data_275),
    .io_pipe_phv_in_data_276(mau_1_io_pipe_phv_in_data_276),
    .io_pipe_phv_in_data_277(mau_1_io_pipe_phv_in_data_277),
    .io_pipe_phv_in_data_278(mau_1_io_pipe_phv_in_data_278),
    .io_pipe_phv_in_data_279(mau_1_io_pipe_phv_in_data_279),
    .io_pipe_phv_in_data_280(mau_1_io_pipe_phv_in_data_280),
    .io_pipe_phv_in_data_281(mau_1_io_pipe_phv_in_data_281),
    .io_pipe_phv_in_data_282(mau_1_io_pipe_phv_in_data_282),
    .io_pipe_phv_in_data_283(mau_1_io_pipe_phv_in_data_283),
    .io_pipe_phv_in_data_284(mau_1_io_pipe_phv_in_data_284),
    .io_pipe_phv_in_data_285(mau_1_io_pipe_phv_in_data_285),
    .io_pipe_phv_in_data_286(mau_1_io_pipe_phv_in_data_286),
    .io_pipe_phv_in_data_287(mau_1_io_pipe_phv_in_data_287),
    .io_pipe_phv_in_data_288(mau_1_io_pipe_phv_in_data_288),
    .io_pipe_phv_in_data_289(mau_1_io_pipe_phv_in_data_289),
    .io_pipe_phv_in_data_290(mau_1_io_pipe_phv_in_data_290),
    .io_pipe_phv_in_data_291(mau_1_io_pipe_phv_in_data_291),
    .io_pipe_phv_in_data_292(mau_1_io_pipe_phv_in_data_292),
    .io_pipe_phv_in_data_293(mau_1_io_pipe_phv_in_data_293),
    .io_pipe_phv_in_data_294(mau_1_io_pipe_phv_in_data_294),
    .io_pipe_phv_in_data_295(mau_1_io_pipe_phv_in_data_295),
    .io_pipe_phv_in_data_296(mau_1_io_pipe_phv_in_data_296),
    .io_pipe_phv_in_data_297(mau_1_io_pipe_phv_in_data_297),
    .io_pipe_phv_in_data_298(mau_1_io_pipe_phv_in_data_298),
    .io_pipe_phv_in_data_299(mau_1_io_pipe_phv_in_data_299),
    .io_pipe_phv_in_data_300(mau_1_io_pipe_phv_in_data_300),
    .io_pipe_phv_in_data_301(mau_1_io_pipe_phv_in_data_301),
    .io_pipe_phv_in_data_302(mau_1_io_pipe_phv_in_data_302),
    .io_pipe_phv_in_data_303(mau_1_io_pipe_phv_in_data_303),
    .io_pipe_phv_in_data_304(mau_1_io_pipe_phv_in_data_304),
    .io_pipe_phv_in_data_305(mau_1_io_pipe_phv_in_data_305),
    .io_pipe_phv_in_data_306(mau_1_io_pipe_phv_in_data_306),
    .io_pipe_phv_in_data_307(mau_1_io_pipe_phv_in_data_307),
    .io_pipe_phv_in_data_308(mau_1_io_pipe_phv_in_data_308),
    .io_pipe_phv_in_data_309(mau_1_io_pipe_phv_in_data_309),
    .io_pipe_phv_in_data_310(mau_1_io_pipe_phv_in_data_310),
    .io_pipe_phv_in_data_311(mau_1_io_pipe_phv_in_data_311),
    .io_pipe_phv_in_data_312(mau_1_io_pipe_phv_in_data_312),
    .io_pipe_phv_in_data_313(mau_1_io_pipe_phv_in_data_313),
    .io_pipe_phv_in_data_314(mau_1_io_pipe_phv_in_data_314),
    .io_pipe_phv_in_data_315(mau_1_io_pipe_phv_in_data_315),
    .io_pipe_phv_in_data_316(mau_1_io_pipe_phv_in_data_316),
    .io_pipe_phv_in_data_317(mau_1_io_pipe_phv_in_data_317),
    .io_pipe_phv_in_data_318(mau_1_io_pipe_phv_in_data_318),
    .io_pipe_phv_in_data_319(mau_1_io_pipe_phv_in_data_319),
    .io_pipe_phv_in_data_320(mau_1_io_pipe_phv_in_data_320),
    .io_pipe_phv_in_data_321(mau_1_io_pipe_phv_in_data_321),
    .io_pipe_phv_in_data_322(mau_1_io_pipe_phv_in_data_322),
    .io_pipe_phv_in_data_323(mau_1_io_pipe_phv_in_data_323),
    .io_pipe_phv_in_data_324(mau_1_io_pipe_phv_in_data_324),
    .io_pipe_phv_in_data_325(mau_1_io_pipe_phv_in_data_325),
    .io_pipe_phv_in_data_326(mau_1_io_pipe_phv_in_data_326),
    .io_pipe_phv_in_data_327(mau_1_io_pipe_phv_in_data_327),
    .io_pipe_phv_in_data_328(mau_1_io_pipe_phv_in_data_328),
    .io_pipe_phv_in_data_329(mau_1_io_pipe_phv_in_data_329),
    .io_pipe_phv_in_data_330(mau_1_io_pipe_phv_in_data_330),
    .io_pipe_phv_in_data_331(mau_1_io_pipe_phv_in_data_331),
    .io_pipe_phv_in_data_332(mau_1_io_pipe_phv_in_data_332),
    .io_pipe_phv_in_data_333(mau_1_io_pipe_phv_in_data_333),
    .io_pipe_phv_in_data_334(mau_1_io_pipe_phv_in_data_334),
    .io_pipe_phv_in_data_335(mau_1_io_pipe_phv_in_data_335),
    .io_pipe_phv_in_data_336(mau_1_io_pipe_phv_in_data_336),
    .io_pipe_phv_in_data_337(mau_1_io_pipe_phv_in_data_337),
    .io_pipe_phv_in_data_338(mau_1_io_pipe_phv_in_data_338),
    .io_pipe_phv_in_data_339(mau_1_io_pipe_phv_in_data_339),
    .io_pipe_phv_in_data_340(mau_1_io_pipe_phv_in_data_340),
    .io_pipe_phv_in_data_341(mau_1_io_pipe_phv_in_data_341),
    .io_pipe_phv_in_data_342(mau_1_io_pipe_phv_in_data_342),
    .io_pipe_phv_in_data_343(mau_1_io_pipe_phv_in_data_343),
    .io_pipe_phv_in_data_344(mau_1_io_pipe_phv_in_data_344),
    .io_pipe_phv_in_data_345(mau_1_io_pipe_phv_in_data_345),
    .io_pipe_phv_in_data_346(mau_1_io_pipe_phv_in_data_346),
    .io_pipe_phv_in_data_347(mau_1_io_pipe_phv_in_data_347),
    .io_pipe_phv_in_data_348(mau_1_io_pipe_phv_in_data_348),
    .io_pipe_phv_in_data_349(mau_1_io_pipe_phv_in_data_349),
    .io_pipe_phv_in_data_350(mau_1_io_pipe_phv_in_data_350),
    .io_pipe_phv_in_data_351(mau_1_io_pipe_phv_in_data_351),
    .io_pipe_phv_in_data_352(mau_1_io_pipe_phv_in_data_352),
    .io_pipe_phv_in_data_353(mau_1_io_pipe_phv_in_data_353),
    .io_pipe_phv_in_data_354(mau_1_io_pipe_phv_in_data_354),
    .io_pipe_phv_in_data_355(mau_1_io_pipe_phv_in_data_355),
    .io_pipe_phv_in_data_356(mau_1_io_pipe_phv_in_data_356),
    .io_pipe_phv_in_data_357(mau_1_io_pipe_phv_in_data_357),
    .io_pipe_phv_in_data_358(mau_1_io_pipe_phv_in_data_358),
    .io_pipe_phv_in_data_359(mau_1_io_pipe_phv_in_data_359),
    .io_pipe_phv_in_data_360(mau_1_io_pipe_phv_in_data_360),
    .io_pipe_phv_in_data_361(mau_1_io_pipe_phv_in_data_361),
    .io_pipe_phv_in_data_362(mau_1_io_pipe_phv_in_data_362),
    .io_pipe_phv_in_data_363(mau_1_io_pipe_phv_in_data_363),
    .io_pipe_phv_in_data_364(mau_1_io_pipe_phv_in_data_364),
    .io_pipe_phv_in_data_365(mau_1_io_pipe_phv_in_data_365),
    .io_pipe_phv_in_data_366(mau_1_io_pipe_phv_in_data_366),
    .io_pipe_phv_in_data_367(mau_1_io_pipe_phv_in_data_367),
    .io_pipe_phv_in_data_368(mau_1_io_pipe_phv_in_data_368),
    .io_pipe_phv_in_data_369(mau_1_io_pipe_phv_in_data_369),
    .io_pipe_phv_in_data_370(mau_1_io_pipe_phv_in_data_370),
    .io_pipe_phv_in_data_371(mau_1_io_pipe_phv_in_data_371),
    .io_pipe_phv_in_data_372(mau_1_io_pipe_phv_in_data_372),
    .io_pipe_phv_in_data_373(mau_1_io_pipe_phv_in_data_373),
    .io_pipe_phv_in_data_374(mau_1_io_pipe_phv_in_data_374),
    .io_pipe_phv_in_data_375(mau_1_io_pipe_phv_in_data_375),
    .io_pipe_phv_in_data_376(mau_1_io_pipe_phv_in_data_376),
    .io_pipe_phv_in_data_377(mau_1_io_pipe_phv_in_data_377),
    .io_pipe_phv_in_data_378(mau_1_io_pipe_phv_in_data_378),
    .io_pipe_phv_in_data_379(mau_1_io_pipe_phv_in_data_379),
    .io_pipe_phv_in_data_380(mau_1_io_pipe_phv_in_data_380),
    .io_pipe_phv_in_data_381(mau_1_io_pipe_phv_in_data_381),
    .io_pipe_phv_in_data_382(mau_1_io_pipe_phv_in_data_382),
    .io_pipe_phv_in_data_383(mau_1_io_pipe_phv_in_data_383),
    .io_pipe_phv_in_data_384(mau_1_io_pipe_phv_in_data_384),
    .io_pipe_phv_in_data_385(mau_1_io_pipe_phv_in_data_385),
    .io_pipe_phv_in_data_386(mau_1_io_pipe_phv_in_data_386),
    .io_pipe_phv_in_data_387(mau_1_io_pipe_phv_in_data_387),
    .io_pipe_phv_in_data_388(mau_1_io_pipe_phv_in_data_388),
    .io_pipe_phv_in_data_389(mau_1_io_pipe_phv_in_data_389),
    .io_pipe_phv_in_data_390(mau_1_io_pipe_phv_in_data_390),
    .io_pipe_phv_in_data_391(mau_1_io_pipe_phv_in_data_391),
    .io_pipe_phv_in_data_392(mau_1_io_pipe_phv_in_data_392),
    .io_pipe_phv_in_data_393(mau_1_io_pipe_phv_in_data_393),
    .io_pipe_phv_in_data_394(mau_1_io_pipe_phv_in_data_394),
    .io_pipe_phv_in_data_395(mau_1_io_pipe_phv_in_data_395),
    .io_pipe_phv_in_data_396(mau_1_io_pipe_phv_in_data_396),
    .io_pipe_phv_in_data_397(mau_1_io_pipe_phv_in_data_397),
    .io_pipe_phv_in_data_398(mau_1_io_pipe_phv_in_data_398),
    .io_pipe_phv_in_data_399(mau_1_io_pipe_phv_in_data_399),
    .io_pipe_phv_in_data_400(mau_1_io_pipe_phv_in_data_400),
    .io_pipe_phv_in_data_401(mau_1_io_pipe_phv_in_data_401),
    .io_pipe_phv_in_data_402(mau_1_io_pipe_phv_in_data_402),
    .io_pipe_phv_in_data_403(mau_1_io_pipe_phv_in_data_403),
    .io_pipe_phv_in_data_404(mau_1_io_pipe_phv_in_data_404),
    .io_pipe_phv_in_data_405(mau_1_io_pipe_phv_in_data_405),
    .io_pipe_phv_in_data_406(mau_1_io_pipe_phv_in_data_406),
    .io_pipe_phv_in_data_407(mau_1_io_pipe_phv_in_data_407),
    .io_pipe_phv_in_data_408(mau_1_io_pipe_phv_in_data_408),
    .io_pipe_phv_in_data_409(mau_1_io_pipe_phv_in_data_409),
    .io_pipe_phv_in_data_410(mau_1_io_pipe_phv_in_data_410),
    .io_pipe_phv_in_data_411(mau_1_io_pipe_phv_in_data_411),
    .io_pipe_phv_in_data_412(mau_1_io_pipe_phv_in_data_412),
    .io_pipe_phv_in_data_413(mau_1_io_pipe_phv_in_data_413),
    .io_pipe_phv_in_data_414(mau_1_io_pipe_phv_in_data_414),
    .io_pipe_phv_in_data_415(mau_1_io_pipe_phv_in_data_415),
    .io_pipe_phv_in_data_416(mau_1_io_pipe_phv_in_data_416),
    .io_pipe_phv_in_data_417(mau_1_io_pipe_phv_in_data_417),
    .io_pipe_phv_in_data_418(mau_1_io_pipe_phv_in_data_418),
    .io_pipe_phv_in_data_419(mau_1_io_pipe_phv_in_data_419),
    .io_pipe_phv_in_data_420(mau_1_io_pipe_phv_in_data_420),
    .io_pipe_phv_in_data_421(mau_1_io_pipe_phv_in_data_421),
    .io_pipe_phv_in_data_422(mau_1_io_pipe_phv_in_data_422),
    .io_pipe_phv_in_data_423(mau_1_io_pipe_phv_in_data_423),
    .io_pipe_phv_in_data_424(mau_1_io_pipe_phv_in_data_424),
    .io_pipe_phv_in_data_425(mau_1_io_pipe_phv_in_data_425),
    .io_pipe_phv_in_data_426(mau_1_io_pipe_phv_in_data_426),
    .io_pipe_phv_in_data_427(mau_1_io_pipe_phv_in_data_427),
    .io_pipe_phv_in_data_428(mau_1_io_pipe_phv_in_data_428),
    .io_pipe_phv_in_data_429(mau_1_io_pipe_phv_in_data_429),
    .io_pipe_phv_in_data_430(mau_1_io_pipe_phv_in_data_430),
    .io_pipe_phv_in_data_431(mau_1_io_pipe_phv_in_data_431),
    .io_pipe_phv_in_data_432(mau_1_io_pipe_phv_in_data_432),
    .io_pipe_phv_in_data_433(mau_1_io_pipe_phv_in_data_433),
    .io_pipe_phv_in_data_434(mau_1_io_pipe_phv_in_data_434),
    .io_pipe_phv_in_data_435(mau_1_io_pipe_phv_in_data_435),
    .io_pipe_phv_in_data_436(mau_1_io_pipe_phv_in_data_436),
    .io_pipe_phv_in_data_437(mau_1_io_pipe_phv_in_data_437),
    .io_pipe_phv_in_data_438(mau_1_io_pipe_phv_in_data_438),
    .io_pipe_phv_in_data_439(mau_1_io_pipe_phv_in_data_439),
    .io_pipe_phv_in_data_440(mau_1_io_pipe_phv_in_data_440),
    .io_pipe_phv_in_data_441(mau_1_io_pipe_phv_in_data_441),
    .io_pipe_phv_in_data_442(mau_1_io_pipe_phv_in_data_442),
    .io_pipe_phv_in_data_443(mau_1_io_pipe_phv_in_data_443),
    .io_pipe_phv_in_data_444(mau_1_io_pipe_phv_in_data_444),
    .io_pipe_phv_in_data_445(mau_1_io_pipe_phv_in_data_445),
    .io_pipe_phv_in_data_446(mau_1_io_pipe_phv_in_data_446),
    .io_pipe_phv_in_data_447(mau_1_io_pipe_phv_in_data_447),
    .io_pipe_phv_in_data_448(mau_1_io_pipe_phv_in_data_448),
    .io_pipe_phv_in_data_449(mau_1_io_pipe_phv_in_data_449),
    .io_pipe_phv_in_data_450(mau_1_io_pipe_phv_in_data_450),
    .io_pipe_phv_in_data_451(mau_1_io_pipe_phv_in_data_451),
    .io_pipe_phv_in_data_452(mau_1_io_pipe_phv_in_data_452),
    .io_pipe_phv_in_data_453(mau_1_io_pipe_phv_in_data_453),
    .io_pipe_phv_in_data_454(mau_1_io_pipe_phv_in_data_454),
    .io_pipe_phv_in_data_455(mau_1_io_pipe_phv_in_data_455),
    .io_pipe_phv_in_data_456(mau_1_io_pipe_phv_in_data_456),
    .io_pipe_phv_in_data_457(mau_1_io_pipe_phv_in_data_457),
    .io_pipe_phv_in_data_458(mau_1_io_pipe_phv_in_data_458),
    .io_pipe_phv_in_data_459(mau_1_io_pipe_phv_in_data_459),
    .io_pipe_phv_in_data_460(mau_1_io_pipe_phv_in_data_460),
    .io_pipe_phv_in_data_461(mau_1_io_pipe_phv_in_data_461),
    .io_pipe_phv_in_data_462(mau_1_io_pipe_phv_in_data_462),
    .io_pipe_phv_in_data_463(mau_1_io_pipe_phv_in_data_463),
    .io_pipe_phv_in_data_464(mau_1_io_pipe_phv_in_data_464),
    .io_pipe_phv_in_data_465(mau_1_io_pipe_phv_in_data_465),
    .io_pipe_phv_in_data_466(mau_1_io_pipe_phv_in_data_466),
    .io_pipe_phv_in_data_467(mau_1_io_pipe_phv_in_data_467),
    .io_pipe_phv_in_data_468(mau_1_io_pipe_phv_in_data_468),
    .io_pipe_phv_in_data_469(mau_1_io_pipe_phv_in_data_469),
    .io_pipe_phv_in_data_470(mau_1_io_pipe_phv_in_data_470),
    .io_pipe_phv_in_data_471(mau_1_io_pipe_phv_in_data_471),
    .io_pipe_phv_in_data_472(mau_1_io_pipe_phv_in_data_472),
    .io_pipe_phv_in_data_473(mau_1_io_pipe_phv_in_data_473),
    .io_pipe_phv_in_data_474(mau_1_io_pipe_phv_in_data_474),
    .io_pipe_phv_in_data_475(mau_1_io_pipe_phv_in_data_475),
    .io_pipe_phv_in_data_476(mau_1_io_pipe_phv_in_data_476),
    .io_pipe_phv_in_data_477(mau_1_io_pipe_phv_in_data_477),
    .io_pipe_phv_in_data_478(mau_1_io_pipe_phv_in_data_478),
    .io_pipe_phv_in_data_479(mau_1_io_pipe_phv_in_data_479),
    .io_pipe_phv_in_data_480(mau_1_io_pipe_phv_in_data_480),
    .io_pipe_phv_in_data_481(mau_1_io_pipe_phv_in_data_481),
    .io_pipe_phv_in_data_482(mau_1_io_pipe_phv_in_data_482),
    .io_pipe_phv_in_data_483(mau_1_io_pipe_phv_in_data_483),
    .io_pipe_phv_in_data_484(mau_1_io_pipe_phv_in_data_484),
    .io_pipe_phv_in_data_485(mau_1_io_pipe_phv_in_data_485),
    .io_pipe_phv_in_data_486(mau_1_io_pipe_phv_in_data_486),
    .io_pipe_phv_in_data_487(mau_1_io_pipe_phv_in_data_487),
    .io_pipe_phv_in_data_488(mau_1_io_pipe_phv_in_data_488),
    .io_pipe_phv_in_data_489(mau_1_io_pipe_phv_in_data_489),
    .io_pipe_phv_in_data_490(mau_1_io_pipe_phv_in_data_490),
    .io_pipe_phv_in_data_491(mau_1_io_pipe_phv_in_data_491),
    .io_pipe_phv_in_data_492(mau_1_io_pipe_phv_in_data_492),
    .io_pipe_phv_in_data_493(mau_1_io_pipe_phv_in_data_493),
    .io_pipe_phv_in_data_494(mau_1_io_pipe_phv_in_data_494),
    .io_pipe_phv_in_data_495(mau_1_io_pipe_phv_in_data_495),
    .io_pipe_phv_in_data_496(mau_1_io_pipe_phv_in_data_496),
    .io_pipe_phv_in_data_497(mau_1_io_pipe_phv_in_data_497),
    .io_pipe_phv_in_data_498(mau_1_io_pipe_phv_in_data_498),
    .io_pipe_phv_in_data_499(mau_1_io_pipe_phv_in_data_499),
    .io_pipe_phv_in_data_500(mau_1_io_pipe_phv_in_data_500),
    .io_pipe_phv_in_data_501(mau_1_io_pipe_phv_in_data_501),
    .io_pipe_phv_in_data_502(mau_1_io_pipe_phv_in_data_502),
    .io_pipe_phv_in_data_503(mau_1_io_pipe_phv_in_data_503),
    .io_pipe_phv_in_data_504(mau_1_io_pipe_phv_in_data_504),
    .io_pipe_phv_in_data_505(mau_1_io_pipe_phv_in_data_505),
    .io_pipe_phv_in_data_506(mau_1_io_pipe_phv_in_data_506),
    .io_pipe_phv_in_data_507(mau_1_io_pipe_phv_in_data_507),
    .io_pipe_phv_in_data_508(mau_1_io_pipe_phv_in_data_508),
    .io_pipe_phv_in_data_509(mau_1_io_pipe_phv_in_data_509),
    .io_pipe_phv_in_data_510(mau_1_io_pipe_phv_in_data_510),
    .io_pipe_phv_in_data_511(mau_1_io_pipe_phv_in_data_511),
    .io_pipe_phv_in_header_0(mau_1_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(mau_1_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(mau_1_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(mau_1_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(mau_1_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(mau_1_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(mau_1_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(mau_1_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(mau_1_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(mau_1_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(mau_1_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(mau_1_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(mau_1_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(mau_1_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(mau_1_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(mau_1_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(mau_1_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(mau_1_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(mau_1_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(mau_1_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(mau_1_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(mau_1_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(mau_1_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(mau_1_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(mau_1_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(mau_1_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(mau_1_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(mau_1_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(mau_1_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(mau_1_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(mau_1_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(mau_1_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(mau_1_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(mau_1_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(mau_1_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(mau_1_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(mau_1_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(mau_1_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(mau_1_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(mau_1_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(mau_1_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(mau_1_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(mau_1_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(mau_1_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(mau_1_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(mau_1_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(mau_1_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(mau_1_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(mau_1_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(mau_1_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(mau_1_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(mau_1_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(mau_1_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(mau_1_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(mau_1_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(mau_1_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(mau_1_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(mau_1_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(mau_1_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(mau_1_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(mau_1_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(mau_1_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(mau_1_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(mau_1_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(mau_1_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(mau_1_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(mau_1_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(mau_1_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(mau_1_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(mau_1_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(mau_1_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(mau_1_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(mau_1_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(mau_1_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(mau_1_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(mau_1_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(mau_1_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(mau_1_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(mau_1_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(mau_1_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(mau_1_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(mau_1_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(mau_1_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(mau_1_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(mau_1_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(mau_1_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(mau_1_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(mau_1_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(mau_1_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(mau_1_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(mau_1_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(mau_1_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(mau_1_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(mau_1_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(mau_1_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(mau_1_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(mau_1_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(mau_1_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(mau_1_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(mau_1_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(mau_1_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(mau_1_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(mau_1_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(mau_1_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(mau_1_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(mau_1_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(mau_1_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(mau_1_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(mau_1_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(mau_1_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(mau_1_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(mau_1_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(mau_1_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(mau_1_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(mau_1_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(mau_1_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(mau_1_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(mau_1_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(mau_1_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(mau_1_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(mau_1_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(mau_1_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(mau_1_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(mau_1_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(mau_1_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(mau_1_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(mau_1_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(mau_1_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(mau_1_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(mau_1_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(mau_1_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(mau_1_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(mau_1_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(mau_1_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(mau_1_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(mau_1_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(mau_1_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(mau_1_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(mau_1_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(mau_1_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(mau_1_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(mau_1_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(mau_1_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(mau_1_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(mau_1_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(mau_1_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(mau_1_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(mau_1_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(mau_1_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(mau_1_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(mau_1_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(mau_1_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(mau_1_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(mau_1_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(mau_1_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(mau_1_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(mau_1_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(mau_1_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(mau_1_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(mau_1_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(mau_1_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(mau_1_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(mau_1_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(mau_1_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(mau_1_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(mau_1_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(mau_1_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(mau_1_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(mau_1_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(mau_1_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(mau_1_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(mau_1_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(mau_1_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(mau_1_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(mau_1_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(mau_1_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(mau_1_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(mau_1_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(mau_1_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(mau_1_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(mau_1_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(mau_1_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(mau_1_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(mau_1_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(mau_1_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(mau_1_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(mau_1_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(mau_1_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(mau_1_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(mau_1_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(mau_1_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(mau_1_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(mau_1_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(mau_1_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(mau_1_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(mau_1_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(mau_1_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(mau_1_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(mau_1_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(mau_1_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(mau_1_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(mau_1_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(mau_1_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(mau_1_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(mau_1_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(mau_1_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(mau_1_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(mau_1_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(mau_1_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(mau_1_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(mau_1_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(mau_1_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(mau_1_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(mau_1_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(mau_1_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(mau_1_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(mau_1_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(mau_1_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(mau_1_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(mau_1_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(mau_1_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(mau_1_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(mau_1_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(mau_1_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(mau_1_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(mau_1_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(mau_1_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(mau_1_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(mau_1_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(mau_1_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(mau_1_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(mau_1_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(mau_1_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(mau_1_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(mau_1_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(mau_1_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(mau_1_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(mau_1_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(mau_1_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(mau_1_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(mau_1_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(mau_1_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(mau_1_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(mau_1_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(mau_1_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(mau_1_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(mau_1_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(mau_1_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(mau_1_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(mau_1_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(mau_1_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(mau_1_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(mau_1_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(mau_1_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(mau_1_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(mau_1_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(mau_1_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(mau_1_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(mau_1_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(mau_1_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(mau_1_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(mau_1_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(mau_1_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(mau_1_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(mau_1_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(mau_1_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(mau_1_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(mau_1_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(mau_1_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(mau_1_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(mau_1_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(mau_1_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(mau_1_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(mau_1_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(mau_1_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(mau_1_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(mau_1_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(mau_1_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_data_256(mau_1_io_pipe_phv_out_data_256),
    .io_pipe_phv_out_data_257(mau_1_io_pipe_phv_out_data_257),
    .io_pipe_phv_out_data_258(mau_1_io_pipe_phv_out_data_258),
    .io_pipe_phv_out_data_259(mau_1_io_pipe_phv_out_data_259),
    .io_pipe_phv_out_data_260(mau_1_io_pipe_phv_out_data_260),
    .io_pipe_phv_out_data_261(mau_1_io_pipe_phv_out_data_261),
    .io_pipe_phv_out_data_262(mau_1_io_pipe_phv_out_data_262),
    .io_pipe_phv_out_data_263(mau_1_io_pipe_phv_out_data_263),
    .io_pipe_phv_out_data_264(mau_1_io_pipe_phv_out_data_264),
    .io_pipe_phv_out_data_265(mau_1_io_pipe_phv_out_data_265),
    .io_pipe_phv_out_data_266(mau_1_io_pipe_phv_out_data_266),
    .io_pipe_phv_out_data_267(mau_1_io_pipe_phv_out_data_267),
    .io_pipe_phv_out_data_268(mau_1_io_pipe_phv_out_data_268),
    .io_pipe_phv_out_data_269(mau_1_io_pipe_phv_out_data_269),
    .io_pipe_phv_out_data_270(mau_1_io_pipe_phv_out_data_270),
    .io_pipe_phv_out_data_271(mau_1_io_pipe_phv_out_data_271),
    .io_pipe_phv_out_data_272(mau_1_io_pipe_phv_out_data_272),
    .io_pipe_phv_out_data_273(mau_1_io_pipe_phv_out_data_273),
    .io_pipe_phv_out_data_274(mau_1_io_pipe_phv_out_data_274),
    .io_pipe_phv_out_data_275(mau_1_io_pipe_phv_out_data_275),
    .io_pipe_phv_out_data_276(mau_1_io_pipe_phv_out_data_276),
    .io_pipe_phv_out_data_277(mau_1_io_pipe_phv_out_data_277),
    .io_pipe_phv_out_data_278(mau_1_io_pipe_phv_out_data_278),
    .io_pipe_phv_out_data_279(mau_1_io_pipe_phv_out_data_279),
    .io_pipe_phv_out_data_280(mau_1_io_pipe_phv_out_data_280),
    .io_pipe_phv_out_data_281(mau_1_io_pipe_phv_out_data_281),
    .io_pipe_phv_out_data_282(mau_1_io_pipe_phv_out_data_282),
    .io_pipe_phv_out_data_283(mau_1_io_pipe_phv_out_data_283),
    .io_pipe_phv_out_data_284(mau_1_io_pipe_phv_out_data_284),
    .io_pipe_phv_out_data_285(mau_1_io_pipe_phv_out_data_285),
    .io_pipe_phv_out_data_286(mau_1_io_pipe_phv_out_data_286),
    .io_pipe_phv_out_data_287(mau_1_io_pipe_phv_out_data_287),
    .io_pipe_phv_out_data_288(mau_1_io_pipe_phv_out_data_288),
    .io_pipe_phv_out_data_289(mau_1_io_pipe_phv_out_data_289),
    .io_pipe_phv_out_data_290(mau_1_io_pipe_phv_out_data_290),
    .io_pipe_phv_out_data_291(mau_1_io_pipe_phv_out_data_291),
    .io_pipe_phv_out_data_292(mau_1_io_pipe_phv_out_data_292),
    .io_pipe_phv_out_data_293(mau_1_io_pipe_phv_out_data_293),
    .io_pipe_phv_out_data_294(mau_1_io_pipe_phv_out_data_294),
    .io_pipe_phv_out_data_295(mau_1_io_pipe_phv_out_data_295),
    .io_pipe_phv_out_data_296(mau_1_io_pipe_phv_out_data_296),
    .io_pipe_phv_out_data_297(mau_1_io_pipe_phv_out_data_297),
    .io_pipe_phv_out_data_298(mau_1_io_pipe_phv_out_data_298),
    .io_pipe_phv_out_data_299(mau_1_io_pipe_phv_out_data_299),
    .io_pipe_phv_out_data_300(mau_1_io_pipe_phv_out_data_300),
    .io_pipe_phv_out_data_301(mau_1_io_pipe_phv_out_data_301),
    .io_pipe_phv_out_data_302(mau_1_io_pipe_phv_out_data_302),
    .io_pipe_phv_out_data_303(mau_1_io_pipe_phv_out_data_303),
    .io_pipe_phv_out_data_304(mau_1_io_pipe_phv_out_data_304),
    .io_pipe_phv_out_data_305(mau_1_io_pipe_phv_out_data_305),
    .io_pipe_phv_out_data_306(mau_1_io_pipe_phv_out_data_306),
    .io_pipe_phv_out_data_307(mau_1_io_pipe_phv_out_data_307),
    .io_pipe_phv_out_data_308(mau_1_io_pipe_phv_out_data_308),
    .io_pipe_phv_out_data_309(mau_1_io_pipe_phv_out_data_309),
    .io_pipe_phv_out_data_310(mau_1_io_pipe_phv_out_data_310),
    .io_pipe_phv_out_data_311(mau_1_io_pipe_phv_out_data_311),
    .io_pipe_phv_out_data_312(mau_1_io_pipe_phv_out_data_312),
    .io_pipe_phv_out_data_313(mau_1_io_pipe_phv_out_data_313),
    .io_pipe_phv_out_data_314(mau_1_io_pipe_phv_out_data_314),
    .io_pipe_phv_out_data_315(mau_1_io_pipe_phv_out_data_315),
    .io_pipe_phv_out_data_316(mau_1_io_pipe_phv_out_data_316),
    .io_pipe_phv_out_data_317(mau_1_io_pipe_phv_out_data_317),
    .io_pipe_phv_out_data_318(mau_1_io_pipe_phv_out_data_318),
    .io_pipe_phv_out_data_319(mau_1_io_pipe_phv_out_data_319),
    .io_pipe_phv_out_data_320(mau_1_io_pipe_phv_out_data_320),
    .io_pipe_phv_out_data_321(mau_1_io_pipe_phv_out_data_321),
    .io_pipe_phv_out_data_322(mau_1_io_pipe_phv_out_data_322),
    .io_pipe_phv_out_data_323(mau_1_io_pipe_phv_out_data_323),
    .io_pipe_phv_out_data_324(mau_1_io_pipe_phv_out_data_324),
    .io_pipe_phv_out_data_325(mau_1_io_pipe_phv_out_data_325),
    .io_pipe_phv_out_data_326(mau_1_io_pipe_phv_out_data_326),
    .io_pipe_phv_out_data_327(mau_1_io_pipe_phv_out_data_327),
    .io_pipe_phv_out_data_328(mau_1_io_pipe_phv_out_data_328),
    .io_pipe_phv_out_data_329(mau_1_io_pipe_phv_out_data_329),
    .io_pipe_phv_out_data_330(mau_1_io_pipe_phv_out_data_330),
    .io_pipe_phv_out_data_331(mau_1_io_pipe_phv_out_data_331),
    .io_pipe_phv_out_data_332(mau_1_io_pipe_phv_out_data_332),
    .io_pipe_phv_out_data_333(mau_1_io_pipe_phv_out_data_333),
    .io_pipe_phv_out_data_334(mau_1_io_pipe_phv_out_data_334),
    .io_pipe_phv_out_data_335(mau_1_io_pipe_phv_out_data_335),
    .io_pipe_phv_out_data_336(mau_1_io_pipe_phv_out_data_336),
    .io_pipe_phv_out_data_337(mau_1_io_pipe_phv_out_data_337),
    .io_pipe_phv_out_data_338(mau_1_io_pipe_phv_out_data_338),
    .io_pipe_phv_out_data_339(mau_1_io_pipe_phv_out_data_339),
    .io_pipe_phv_out_data_340(mau_1_io_pipe_phv_out_data_340),
    .io_pipe_phv_out_data_341(mau_1_io_pipe_phv_out_data_341),
    .io_pipe_phv_out_data_342(mau_1_io_pipe_phv_out_data_342),
    .io_pipe_phv_out_data_343(mau_1_io_pipe_phv_out_data_343),
    .io_pipe_phv_out_data_344(mau_1_io_pipe_phv_out_data_344),
    .io_pipe_phv_out_data_345(mau_1_io_pipe_phv_out_data_345),
    .io_pipe_phv_out_data_346(mau_1_io_pipe_phv_out_data_346),
    .io_pipe_phv_out_data_347(mau_1_io_pipe_phv_out_data_347),
    .io_pipe_phv_out_data_348(mau_1_io_pipe_phv_out_data_348),
    .io_pipe_phv_out_data_349(mau_1_io_pipe_phv_out_data_349),
    .io_pipe_phv_out_data_350(mau_1_io_pipe_phv_out_data_350),
    .io_pipe_phv_out_data_351(mau_1_io_pipe_phv_out_data_351),
    .io_pipe_phv_out_data_352(mau_1_io_pipe_phv_out_data_352),
    .io_pipe_phv_out_data_353(mau_1_io_pipe_phv_out_data_353),
    .io_pipe_phv_out_data_354(mau_1_io_pipe_phv_out_data_354),
    .io_pipe_phv_out_data_355(mau_1_io_pipe_phv_out_data_355),
    .io_pipe_phv_out_data_356(mau_1_io_pipe_phv_out_data_356),
    .io_pipe_phv_out_data_357(mau_1_io_pipe_phv_out_data_357),
    .io_pipe_phv_out_data_358(mau_1_io_pipe_phv_out_data_358),
    .io_pipe_phv_out_data_359(mau_1_io_pipe_phv_out_data_359),
    .io_pipe_phv_out_data_360(mau_1_io_pipe_phv_out_data_360),
    .io_pipe_phv_out_data_361(mau_1_io_pipe_phv_out_data_361),
    .io_pipe_phv_out_data_362(mau_1_io_pipe_phv_out_data_362),
    .io_pipe_phv_out_data_363(mau_1_io_pipe_phv_out_data_363),
    .io_pipe_phv_out_data_364(mau_1_io_pipe_phv_out_data_364),
    .io_pipe_phv_out_data_365(mau_1_io_pipe_phv_out_data_365),
    .io_pipe_phv_out_data_366(mau_1_io_pipe_phv_out_data_366),
    .io_pipe_phv_out_data_367(mau_1_io_pipe_phv_out_data_367),
    .io_pipe_phv_out_data_368(mau_1_io_pipe_phv_out_data_368),
    .io_pipe_phv_out_data_369(mau_1_io_pipe_phv_out_data_369),
    .io_pipe_phv_out_data_370(mau_1_io_pipe_phv_out_data_370),
    .io_pipe_phv_out_data_371(mau_1_io_pipe_phv_out_data_371),
    .io_pipe_phv_out_data_372(mau_1_io_pipe_phv_out_data_372),
    .io_pipe_phv_out_data_373(mau_1_io_pipe_phv_out_data_373),
    .io_pipe_phv_out_data_374(mau_1_io_pipe_phv_out_data_374),
    .io_pipe_phv_out_data_375(mau_1_io_pipe_phv_out_data_375),
    .io_pipe_phv_out_data_376(mau_1_io_pipe_phv_out_data_376),
    .io_pipe_phv_out_data_377(mau_1_io_pipe_phv_out_data_377),
    .io_pipe_phv_out_data_378(mau_1_io_pipe_phv_out_data_378),
    .io_pipe_phv_out_data_379(mau_1_io_pipe_phv_out_data_379),
    .io_pipe_phv_out_data_380(mau_1_io_pipe_phv_out_data_380),
    .io_pipe_phv_out_data_381(mau_1_io_pipe_phv_out_data_381),
    .io_pipe_phv_out_data_382(mau_1_io_pipe_phv_out_data_382),
    .io_pipe_phv_out_data_383(mau_1_io_pipe_phv_out_data_383),
    .io_pipe_phv_out_data_384(mau_1_io_pipe_phv_out_data_384),
    .io_pipe_phv_out_data_385(mau_1_io_pipe_phv_out_data_385),
    .io_pipe_phv_out_data_386(mau_1_io_pipe_phv_out_data_386),
    .io_pipe_phv_out_data_387(mau_1_io_pipe_phv_out_data_387),
    .io_pipe_phv_out_data_388(mau_1_io_pipe_phv_out_data_388),
    .io_pipe_phv_out_data_389(mau_1_io_pipe_phv_out_data_389),
    .io_pipe_phv_out_data_390(mau_1_io_pipe_phv_out_data_390),
    .io_pipe_phv_out_data_391(mau_1_io_pipe_phv_out_data_391),
    .io_pipe_phv_out_data_392(mau_1_io_pipe_phv_out_data_392),
    .io_pipe_phv_out_data_393(mau_1_io_pipe_phv_out_data_393),
    .io_pipe_phv_out_data_394(mau_1_io_pipe_phv_out_data_394),
    .io_pipe_phv_out_data_395(mau_1_io_pipe_phv_out_data_395),
    .io_pipe_phv_out_data_396(mau_1_io_pipe_phv_out_data_396),
    .io_pipe_phv_out_data_397(mau_1_io_pipe_phv_out_data_397),
    .io_pipe_phv_out_data_398(mau_1_io_pipe_phv_out_data_398),
    .io_pipe_phv_out_data_399(mau_1_io_pipe_phv_out_data_399),
    .io_pipe_phv_out_data_400(mau_1_io_pipe_phv_out_data_400),
    .io_pipe_phv_out_data_401(mau_1_io_pipe_phv_out_data_401),
    .io_pipe_phv_out_data_402(mau_1_io_pipe_phv_out_data_402),
    .io_pipe_phv_out_data_403(mau_1_io_pipe_phv_out_data_403),
    .io_pipe_phv_out_data_404(mau_1_io_pipe_phv_out_data_404),
    .io_pipe_phv_out_data_405(mau_1_io_pipe_phv_out_data_405),
    .io_pipe_phv_out_data_406(mau_1_io_pipe_phv_out_data_406),
    .io_pipe_phv_out_data_407(mau_1_io_pipe_phv_out_data_407),
    .io_pipe_phv_out_data_408(mau_1_io_pipe_phv_out_data_408),
    .io_pipe_phv_out_data_409(mau_1_io_pipe_phv_out_data_409),
    .io_pipe_phv_out_data_410(mau_1_io_pipe_phv_out_data_410),
    .io_pipe_phv_out_data_411(mau_1_io_pipe_phv_out_data_411),
    .io_pipe_phv_out_data_412(mau_1_io_pipe_phv_out_data_412),
    .io_pipe_phv_out_data_413(mau_1_io_pipe_phv_out_data_413),
    .io_pipe_phv_out_data_414(mau_1_io_pipe_phv_out_data_414),
    .io_pipe_phv_out_data_415(mau_1_io_pipe_phv_out_data_415),
    .io_pipe_phv_out_data_416(mau_1_io_pipe_phv_out_data_416),
    .io_pipe_phv_out_data_417(mau_1_io_pipe_phv_out_data_417),
    .io_pipe_phv_out_data_418(mau_1_io_pipe_phv_out_data_418),
    .io_pipe_phv_out_data_419(mau_1_io_pipe_phv_out_data_419),
    .io_pipe_phv_out_data_420(mau_1_io_pipe_phv_out_data_420),
    .io_pipe_phv_out_data_421(mau_1_io_pipe_phv_out_data_421),
    .io_pipe_phv_out_data_422(mau_1_io_pipe_phv_out_data_422),
    .io_pipe_phv_out_data_423(mau_1_io_pipe_phv_out_data_423),
    .io_pipe_phv_out_data_424(mau_1_io_pipe_phv_out_data_424),
    .io_pipe_phv_out_data_425(mau_1_io_pipe_phv_out_data_425),
    .io_pipe_phv_out_data_426(mau_1_io_pipe_phv_out_data_426),
    .io_pipe_phv_out_data_427(mau_1_io_pipe_phv_out_data_427),
    .io_pipe_phv_out_data_428(mau_1_io_pipe_phv_out_data_428),
    .io_pipe_phv_out_data_429(mau_1_io_pipe_phv_out_data_429),
    .io_pipe_phv_out_data_430(mau_1_io_pipe_phv_out_data_430),
    .io_pipe_phv_out_data_431(mau_1_io_pipe_phv_out_data_431),
    .io_pipe_phv_out_data_432(mau_1_io_pipe_phv_out_data_432),
    .io_pipe_phv_out_data_433(mau_1_io_pipe_phv_out_data_433),
    .io_pipe_phv_out_data_434(mau_1_io_pipe_phv_out_data_434),
    .io_pipe_phv_out_data_435(mau_1_io_pipe_phv_out_data_435),
    .io_pipe_phv_out_data_436(mau_1_io_pipe_phv_out_data_436),
    .io_pipe_phv_out_data_437(mau_1_io_pipe_phv_out_data_437),
    .io_pipe_phv_out_data_438(mau_1_io_pipe_phv_out_data_438),
    .io_pipe_phv_out_data_439(mau_1_io_pipe_phv_out_data_439),
    .io_pipe_phv_out_data_440(mau_1_io_pipe_phv_out_data_440),
    .io_pipe_phv_out_data_441(mau_1_io_pipe_phv_out_data_441),
    .io_pipe_phv_out_data_442(mau_1_io_pipe_phv_out_data_442),
    .io_pipe_phv_out_data_443(mau_1_io_pipe_phv_out_data_443),
    .io_pipe_phv_out_data_444(mau_1_io_pipe_phv_out_data_444),
    .io_pipe_phv_out_data_445(mau_1_io_pipe_phv_out_data_445),
    .io_pipe_phv_out_data_446(mau_1_io_pipe_phv_out_data_446),
    .io_pipe_phv_out_data_447(mau_1_io_pipe_phv_out_data_447),
    .io_pipe_phv_out_data_448(mau_1_io_pipe_phv_out_data_448),
    .io_pipe_phv_out_data_449(mau_1_io_pipe_phv_out_data_449),
    .io_pipe_phv_out_data_450(mau_1_io_pipe_phv_out_data_450),
    .io_pipe_phv_out_data_451(mau_1_io_pipe_phv_out_data_451),
    .io_pipe_phv_out_data_452(mau_1_io_pipe_phv_out_data_452),
    .io_pipe_phv_out_data_453(mau_1_io_pipe_phv_out_data_453),
    .io_pipe_phv_out_data_454(mau_1_io_pipe_phv_out_data_454),
    .io_pipe_phv_out_data_455(mau_1_io_pipe_phv_out_data_455),
    .io_pipe_phv_out_data_456(mau_1_io_pipe_phv_out_data_456),
    .io_pipe_phv_out_data_457(mau_1_io_pipe_phv_out_data_457),
    .io_pipe_phv_out_data_458(mau_1_io_pipe_phv_out_data_458),
    .io_pipe_phv_out_data_459(mau_1_io_pipe_phv_out_data_459),
    .io_pipe_phv_out_data_460(mau_1_io_pipe_phv_out_data_460),
    .io_pipe_phv_out_data_461(mau_1_io_pipe_phv_out_data_461),
    .io_pipe_phv_out_data_462(mau_1_io_pipe_phv_out_data_462),
    .io_pipe_phv_out_data_463(mau_1_io_pipe_phv_out_data_463),
    .io_pipe_phv_out_data_464(mau_1_io_pipe_phv_out_data_464),
    .io_pipe_phv_out_data_465(mau_1_io_pipe_phv_out_data_465),
    .io_pipe_phv_out_data_466(mau_1_io_pipe_phv_out_data_466),
    .io_pipe_phv_out_data_467(mau_1_io_pipe_phv_out_data_467),
    .io_pipe_phv_out_data_468(mau_1_io_pipe_phv_out_data_468),
    .io_pipe_phv_out_data_469(mau_1_io_pipe_phv_out_data_469),
    .io_pipe_phv_out_data_470(mau_1_io_pipe_phv_out_data_470),
    .io_pipe_phv_out_data_471(mau_1_io_pipe_phv_out_data_471),
    .io_pipe_phv_out_data_472(mau_1_io_pipe_phv_out_data_472),
    .io_pipe_phv_out_data_473(mau_1_io_pipe_phv_out_data_473),
    .io_pipe_phv_out_data_474(mau_1_io_pipe_phv_out_data_474),
    .io_pipe_phv_out_data_475(mau_1_io_pipe_phv_out_data_475),
    .io_pipe_phv_out_data_476(mau_1_io_pipe_phv_out_data_476),
    .io_pipe_phv_out_data_477(mau_1_io_pipe_phv_out_data_477),
    .io_pipe_phv_out_data_478(mau_1_io_pipe_phv_out_data_478),
    .io_pipe_phv_out_data_479(mau_1_io_pipe_phv_out_data_479),
    .io_pipe_phv_out_data_480(mau_1_io_pipe_phv_out_data_480),
    .io_pipe_phv_out_data_481(mau_1_io_pipe_phv_out_data_481),
    .io_pipe_phv_out_data_482(mau_1_io_pipe_phv_out_data_482),
    .io_pipe_phv_out_data_483(mau_1_io_pipe_phv_out_data_483),
    .io_pipe_phv_out_data_484(mau_1_io_pipe_phv_out_data_484),
    .io_pipe_phv_out_data_485(mau_1_io_pipe_phv_out_data_485),
    .io_pipe_phv_out_data_486(mau_1_io_pipe_phv_out_data_486),
    .io_pipe_phv_out_data_487(mau_1_io_pipe_phv_out_data_487),
    .io_pipe_phv_out_data_488(mau_1_io_pipe_phv_out_data_488),
    .io_pipe_phv_out_data_489(mau_1_io_pipe_phv_out_data_489),
    .io_pipe_phv_out_data_490(mau_1_io_pipe_phv_out_data_490),
    .io_pipe_phv_out_data_491(mau_1_io_pipe_phv_out_data_491),
    .io_pipe_phv_out_data_492(mau_1_io_pipe_phv_out_data_492),
    .io_pipe_phv_out_data_493(mau_1_io_pipe_phv_out_data_493),
    .io_pipe_phv_out_data_494(mau_1_io_pipe_phv_out_data_494),
    .io_pipe_phv_out_data_495(mau_1_io_pipe_phv_out_data_495),
    .io_pipe_phv_out_data_496(mau_1_io_pipe_phv_out_data_496),
    .io_pipe_phv_out_data_497(mau_1_io_pipe_phv_out_data_497),
    .io_pipe_phv_out_data_498(mau_1_io_pipe_phv_out_data_498),
    .io_pipe_phv_out_data_499(mau_1_io_pipe_phv_out_data_499),
    .io_pipe_phv_out_data_500(mau_1_io_pipe_phv_out_data_500),
    .io_pipe_phv_out_data_501(mau_1_io_pipe_phv_out_data_501),
    .io_pipe_phv_out_data_502(mau_1_io_pipe_phv_out_data_502),
    .io_pipe_phv_out_data_503(mau_1_io_pipe_phv_out_data_503),
    .io_pipe_phv_out_data_504(mau_1_io_pipe_phv_out_data_504),
    .io_pipe_phv_out_data_505(mau_1_io_pipe_phv_out_data_505),
    .io_pipe_phv_out_data_506(mau_1_io_pipe_phv_out_data_506),
    .io_pipe_phv_out_data_507(mau_1_io_pipe_phv_out_data_507),
    .io_pipe_phv_out_data_508(mau_1_io_pipe_phv_out_data_508),
    .io_pipe_phv_out_data_509(mau_1_io_pipe_phv_out_data_509),
    .io_pipe_phv_out_data_510(mau_1_io_pipe_phv_out_data_510),
    .io_pipe_phv_out_data_511(mau_1_io_pipe_phv_out_data_511),
    .io_pipe_phv_out_header_0(mau_1_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(mau_1_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(mau_1_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(mau_1_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(mau_1_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(mau_1_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(mau_1_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(mau_1_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(mau_1_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(mau_1_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(mau_1_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(mau_1_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(mau_1_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(mau_1_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(mau_1_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(mau_1_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(mau_1_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(mau_1_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(mau_1_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(mau_1_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(mau_1_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(mau_1_io_pipe_phv_out_is_valid_processor),
    .io_mod_state_id_mod(mau_1_io_mod_state_id_mod),
    .io_mod_state_id(mau_1_io_mod_state_id),
    .io_mod_sram_w_cs(mau_1_io_mod_sram_w_cs),
    .io_mod_sram_w_en(mau_1_io_mod_sram_w_en),
    .io_mod_sram_w_addr(mau_1_io_mod_sram_w_addr),
    .io_mod_sram_w_data(mau_1_io_mod_sram_w_data)
  );
  ParseModule mau_2 ( // @[parser_pisa.scala 31:25]
    .clock(mau_2_clock),
    .io_pipe_phv_in_data_0(mau_2_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(mau_2_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(mau_2_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(mau_2_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(mau_2_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(mau_2_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(mau_2_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(mau_2_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(mau_2_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(mau_2_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(mau_2_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(mau_2_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(mau_2_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(mau_2_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(mau_2_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(mau_2_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(mau_2_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(mau_2_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(mau_2_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(mau_2_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(mau_2_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(mau_2_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(mau_2_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(mau_2_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(mau_2_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(mau_2_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(mau_2_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(mau_2_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(mau_2_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(mau_2_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(mau_2_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(mau_2_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(mau_2_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(mau_2_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(mau_2_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(mau_2_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(mau_2_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(mau_2_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(mau_2_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(mau_2_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(mau_2_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(mau_2_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(mau_2_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(mau_2_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(mau_2_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(mau_2_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(mau_2_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(mau_2_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(mau_2_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(mau_2_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(mau_2_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(mau_2_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(mau_2_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(mau_2_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(mau_2_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(mau_2_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(mau_2_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(mau_2_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(mau_2_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(mau_2_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(mau_2_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(mau_2_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(mau_2_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(mau_2_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(mau_2_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(mau_2_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(mau_2_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(mau_2_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(mau_2_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(mau_2_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(mau_2_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(mau_2_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(mau_2_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(mau_2_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(mau_2_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(mau_2_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(mau_2_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(mau_2_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(mau_2_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(mau_2_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(mau_2_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(mau_2_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(mau_2_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(mau_2_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(mau_2_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(mau_2_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(mau_2_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(mau_2_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(mau_2_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(mau_2_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(mau_2_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(mau_2_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(mau_2_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(mau_2_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(mau_2_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(mau_2_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(mau_2_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(mau_2_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(mau_2_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(mau_2_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(mau_2_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(mau_2_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(mau_2_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(mau_2_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(mau_2_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(mau_2_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(mau_2_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(mau_2_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(mau_2_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(mau_2_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(mau_2_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(mau_2_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(mau_2_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(mau_2_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(mau_2_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(mau_2_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(mau_2_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(mau_2_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(mau_2_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(mau_2_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(mau_2_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(mau_2_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(mau_2_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(mau_2_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(mau_2_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(mau_2_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(mau_2_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(mau_2_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(mau_2_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(mau_2_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(mau_2_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(mau_2_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(mau_2_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(mau_2_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(mau_2_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(mau_2_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(mau_2_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(mau_2_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(mau_2_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(mau_2_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(mau_2_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(mau_2_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(mau_2_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(mau_2_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(mau_2_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(mau_2_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(mau_2_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(mau_2_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(mau_2_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(mau_2_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(mau_2_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(mau_2_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(mau_2_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(mau_2_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(mau_2_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(mau_2_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(mau_2_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(mau_2_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(mau_2_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(mau_2_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(mau_2_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(mau_2_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(mau_2_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(mau_2_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(mau_2_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(mau_2_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(mau_2_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(mau_2_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(mau_2_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(mau_2_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(mau_2_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(mau_2_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(mau_2_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(mau_2_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(mau_2_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(mau_2_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(mau_2_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(mau_2_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(mau_2_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(mau_2_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(mau_2_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(mau_2_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(mau_2_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(mau_2_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(mau_2_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(mau_2_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(mau_2_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(mau_2_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(mau_2_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(mau_2_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(mau_2_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(mau_2_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(mau_2_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(mau_2_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(mau_2_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(mau_2_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(mau_2_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(mau_2_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(mau_2_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(mau_2_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(mau_2_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(mau_2_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(mau_2_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(mau_2_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(mau_2_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(mau_2_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(mau_2_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(mau_2_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(mau_2_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(mau_2_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(mau_2_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(mau_2_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(mau_2_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(mau_2_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(mau_2_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(mau_2_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(mau_2_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(mau_2_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(mau_2_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(mau_2_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(mau_2_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(mau_2_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(mau_2_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(mau_2_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(mau_2_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(mau_2_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(mau_2_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(mau_2_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(mau_2_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(mau_2_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(mau_2_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(mau_2_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(mau_2_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(mau_2_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(mau_2_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(mau_2_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(mau_2_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(mau_2_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(mau_2_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(mau_2_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(mau_2_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(mau_2_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(mau_2_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(mau_2_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(mau_2_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(mau_2_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(mau_2_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(mau_2_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(mau_2_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(mau_2_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(mau_2_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(mau_2_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(mau_2_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(mau_2_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(mau_2_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(mau_2_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_data_256(mau_2_io_pipe_phv_in_data_256),
    .io_pipe_phv_in_data_257(mau_2_io_pipe_phv_in_data_257),
    .io_pipe_phv_in_data_258(mau_2_io_pipe_phv_in_data_258),
    .io_pipe_phv_in_data_259(mau_2_io_pipe_phv_in_data_259),
    .io_pipe_phv_in_data_260(mau_2_io_pipe_phv_in_data_260),
    .io_pipe_phv_in_data_261(mau_2_io_pipe_phv_in_data_261),
    .io_pipe_phv_in_data_262(mau_2_io_pipe_phv_in_data_262),
    .io_pipe_phv_in_data_263(mau_2_io_pipe_phv_in_data_263),
    .io_pipe_phv_in_data_264(mau_2_io_pipe_phv_in_data_264),
    .io_pipe_phv_in_data_265(mau_2_io_pipe_phv_in_data_265),
    .io_pipe_phv_in_data_266(mau_2_io_pipe_phv_in_data_266),
    .io_pipe_phv_in_data_267(mau_2_io_pipe_phv_in_data_267),
    .io_pipe_phv_in_data_268(mau_2_io_pipe_phv_in_data_268),
    .io_pipe_phv_in_data_269(mau_2_io_pipe_phv_in_data_269),
    .io_pipe_phv_in_data_270(mau_2_io_pipe_phv_in_data_270),
    .io_pipe_phv_in_data_271(mau_2_io_pipe_phv_in_data_271),
    .io_pipe_phv_in_data_272(mau_2_io_pipe_phv_in_data_272),
    .io_pipe_phv_in_data_273(mau_2_io_pipe_phv_in_data_273),
    .io_pipe_phv_in_data_274(mau_2_io_pipe_phv_in_data_274),
    .io_pipe_phv_in_data_275(mau_2_io_pipe_phv_in_data_275),
    .io_pipe_phv_in_data_276(mau_2_io_pipe_phv_in_data_276),
    .io_pipe_phv_in_data_277(mau_2_io_pipe_phv_in_data_277),
    .io_pipe_phv_in_data_278(mau_2_io_pipe_phv_in_data_278),
    .io_pipe_phv_in_data_279(mau_2_io_pipe_phv_in_data_279),
    .io_pipe_phv_in_data_280(mau_2_io_pipe_phv_in_data_280),
    .io_pipe_phv_in_data_281(mau_2_io_pipe_phv_in_data_281),
    .io_pipe_phv_in_data_282(mau_2_io_pipe_phv_in_data_282),
    .io_pipe_phv_in_data_283(mau_2_io_pipe_phv_in_data_283),
    .io_pipe_phv_in_data_284(mau_2_io_pipe_phv_in_data_284),
    .io_pipe_phv_in_data_285(mau_2_io_pipe_phv_in_data_285),
    .io_pipe_phv_in_data_286(mau_2_io_pipe_phv_in_data_286),
    .io_pipe_phv_in_data_287(mau_2_io_pipe_phv_in_data_287),
    .io_pipe_phv_in_data_288(mau_2_io_pipe_phv_in_data_288),
    .io_pipe_phv_in_data_289(mau_2_io_pipe_phv_in_data_289),
    .io_pipe_phv_in_data_290(mau_2_io_pipe_phv_in_data_290),
    .io_pipe_phv_in_data_291(mau_2_io_pipe_phv_in_data_291),
    .io_pipe_phv_in_data_292(mau_2_io_pipe_phv_in_data_292),
    .io_pipe_phv_in_data_293(mau_2_io_pipe_phv_in_data_293),
    .io_pipe_phv_in_data_294(mau_2_io_pipe_phv_in_data_294),
    .io_pipe_phv_in_data_295(mau_2_io_pipe_phv_in_data_295),
    .io_pipe_phv_in_data_296(mau_2_io_pipe_phv_in_data_296),
    .io_pipe_phv_in_data_297(mau_2_io_pipe_phv_in_data_297),
    .io_pipe_phv_in_data_298(mau_2_io_pipe_phv_in_data_298),
    .io_pipe_phv_in_data_299(mau_2_io_pipe_phv_in_data_299),
    .io_pipe_phv_in_data_300(mau_2_io_pipe_phv_in_data_300),
    .io_pipe_phv_in_data_301(mau_2_io_pipe_phv_in_data_301),
    .io_pipe_phv_in_data_302(mau_2_io_pipe_phv_in_data_302),
    .io_pipe_phv_in_data_303(mau_2_io_pipe_phv_in_data_303),
    .io_pipe_phv_in_data_304(mau_2_io_pipe_phv_in_data_304),
    .io_pipe_phv_in_data_305(mau_2_io_pipe_phv_in_data_305),
    .io_pipe_phv_in_data_306(mau_2_io_pipe_phv_in_data_306),
    .io_pipe_phv_in_data_307(mau_2_io_pipe_phv_in_data_307),
    .io_pipe_phv_in_data_308(mau_2_io_pipe_phv_in_data_308),
    .io_pipe_phv_in_data_309(mau_2_io_pipe_phv_in_data_309),
    .io_pipe_phv_in_data_310(mau_2_io_pipe_phv_in_data_310),
    .io_pipe_phv_in_data_311(mau_2_io_pipe_phv_in_data_311),
    .io_pipe_phv_in_data_312(mau_2_io_pipe_phv_in_data_312),
    .io_pipe_phv_in_data_313(mau_2_io_pipe_phv_in_data_313),
    .io_pipe_phv_in_data_314(mau_2_io_pipe_phv_in_data_314),
    .io_pipe_phv_in_data_315(mau_2_io_pipe_phv_in_data_315),
    .io_pipe_phv_in_data_316(mau_2_io_pipe_phv_in_data_316),
    .io_pipe_phv_in_data_317(mau_2_io_pipe_phv_in_data_317),
    .io_pipe_phv_in_data_318(mau_2_io_pipe_phv_in_data_318),
    .io_pipe_phv_in_data_319(mau_2_io_pipe_phv_in_data_319),
    .io_pipe_phv_in_data_320(mau_2_io_pipe_phv_in_data_320),
    .io_pipe_phv_in_data_321(mau_2_io_pipe_phv_in_data_321),
    .io_pipe_phv_in_data_322(mau_2_io_pipe_phv_in_data_322),
    .io_pipe_phv_in_data_323(mau_2_io_pipe_phv_in_data_323),
    .io_pipe_phv_in_data_324(mau_2_io_pipe_phv_in_data_324),
    .io_pipe_phv_in_data_325(mau_2_io_pipe_phv_in_data_325),
    .io_pipe_phv_in_data_326(mau_2_io_pipe_phv_in_data_326),
    .io_pipe_phv_in_data_327(mau_2_io_pipe_phv_in_data_327),
    .io_pipe_phv_in_data_328(mau_2_io_pipe_phv_in_data_328),
    .io_pipe_phv_in_data_329(mau_2_io_pipe_phv_in_data_329),
    .io_pipe_phv_in_data_330(mau_2_io_pipe_phv_in_data_330),
    .io_pipe_phv_in_data_331(mau_2_io_pipe_phv_in_data_331),
    .io_pipe_phv_in_data_332(mau_2_io_pipe_phv_in_data_332),
    .io_pipe_phv_in_data_333(mau_2_io_pipe_phv_in_data_333),
    .io_pipe_phv_in_data_334(mau_2_io_pipe_phv_in_data_334),
    .io_pipe_phv_in_data_335(mau_2_io_pipe_phv_in_data_335),
    .io_pipe_phv_in_data_336(mau_2_io_pipe_phv_in_data_336),
    .io_pipe_phv_in_data_337(mau_2_io_pipe_phv_in_data_337),
    .io_pipe_phv_in_data_338(mau_2_io_pipe_phv_in_data_338),
    .io_pipe_phv_in_data_339(mau_2_io_pipe_phv_in_data_339),
    .io_pipe_phv_in_data_340(mau_2_io_pipe_phv_in_data_340),
    .io_pipe_phv_in_data_341(mau_2_io_pipe_phv_in_data_341),
    .io_pipe_phv_in_data_342(mau_2_io_pipe_phv_in_data_342),
    .io_pipe_phv_in_data_343(mau_2_io_pipe_phv_in_data_343),
    .io_pipe_phv_in_data_344(mau_2_io_pipe_phv_in_data_344),
    .io_pipe_phv_in_data_345(mau_2_io_pipe_phv_in_data_345),
    .io_pipe_phv_in_data_346(mau_2_io_pipe_phv_in_data_346),
    .io_pipe_phv_in_data_347(mau_2_io_pipe_phv_in_data_347),
    .io_pipe_phv_in_data_348(mau_2_io_pipe_phv_in_data_348),
    .io_pipe_phv_in_data_349(mau_2_io_pipe_phv_in_data_349),
    .io_pipe_phv_in_data_350(mau_2_io_pipe_phv_in_data_350),
    .io_pipe_phv_in_data_351(mau_2_io_pipe_phv_in_data_351),
    .io_pipe_phv_in_data_352(mau_2_io_pipe_phv_in_data_352),
    .io_pipe_phv_in_data_353(mau_2_io_pipe_phv_in_data_353),
    .io_pipe_phv_in_data_354(mau_2_io_pipe_phv_in_data_354),
    .io_pipe_phv_in_data_355(mau_2_io_pipe_phv_in_data_355),
    .io_pipe_phv_in_data_356(mau_2_io_pipe_phv_in_data_356),
    .io_pipe_phv_in_data_357(mau_2_io_pipe_phv_in_data_357),
    .io_pipe_phv_in_data_358(mau_2_io_pipe_phv_in_data_358),
    .io_pipe_phv_in_data_359(mau_2_io_pipe_phv_in_data_359),
    .io_pipe_phv_in_data_360(mau_2_io_pipe_phv_in_data_360),
    .io_pipe_phv_in_data_361(mau_2_io_pipe_phv_in_data_361),
    .io_pipe_phv_in_data_362(mau_2_io_pipe_phv_in_data_362),
    .io_pipe_phv_in_data_363(mau_2_io_pipe_phv_in_data_363),
    .io_pipe_phv_in_data_364(mau_2_io_pipe_phv_in_data_364),
    .io_pipe_phv_in_data_365(mau_2_io_pipe_phv_in_data_365),
    .io_pipe_phv_in_data_366(mau_2_io_pipe_phv_in_data_366),
    .io_pipe_phv_in_data_367(mau_2_io_pipe_phv_in_data_367),
    .io_pipe_phv_in_data_368(mau_2_io_pipe_phv_in_data_368),
    .io_pipe_phv_in_data_369(mau_2_io_pipe_phv_in_data_369),
    .io_pipe_phv_in_data_370(mau_2_io_pipe_phv_in_data_370),
    .io_pipe_phv_in_data_371(mau_2_io_pipe_phv_in_data_371),
    .io_pipe_phv_in_data_372(mau_2_io_pipe_phv_in_data_372),
    .io_pipe_phv_in_data_373(mau_2_io_pipe_phv_in_data_373),
    .io_pipe_phv_in_data_374(mau_2_io_pipe_phv_in_data_374),
    .io_pipe_phv_in_data_375(mau_2_io_pipe_phv_in_data_375),
    .io_pipe_phv_in_data_376(mau_2_io_pipe_phv_in_data_376),
    .io_pipe_phv_in_data_377(mau_2_io_pipe_phv_in_data_377),
    .io_pipe_phv_in_data_378(mau_2_io_pipe_phv_in_data_378),
    .io_pipe_phv_in_data_379(mau_2_io_pipe_phv_in_data_379),
    .io_pipe_phv_in_data_380(mau_2_io_pipe_phv_in_data_380),
    .io_pipe_phv_in_data_381(mau_2_io_pipe_phv_in_data_381),
    .io_pipe_phv_in_data_382(mau_2_io_pipe_phv_in_data_382),
    .io_pipe_phv_in_data_383(mau_2_io_pipe_phv_in_data_383),
    .io_pipe_phv_in_data_384(mau_2_io_pipe_phv_in_data_384),
    .io_pipe_phv_in_data_385(mau_2_io_pipe_phv_in_data_385),
    .io_pipe_phv_in_data_386(mau_2_io_pipe_phv_in_data_386),
    .io_pipe_phv_in_data_387(mau_2_io_pipe_phv_in_data_387),
    .io_pipe_phv_in_data_388(mau_2_io_pipe_phv_in_data_388),
    .io_pipe_phv_in_data_389(mau_2_io_pipe_phv_in_data_389),
    .io_pipe_phv_in_data_390(mau_2_io_pipe_phv_in_data_390),
    .io_pipe_phv_in_data_391(mau_2_io_pipe_phv_in_data_391),
    .io_pipe_phv_in_data_392(mau_2_io_pipe_phv_in_data_392),
    .io_pipe_phv_in_data_393(mau_2_io_pipe_phv_in_data_393),
    .io_pipe_phv_in_data_394(mau_2_io_pipe_phv_in_data_394),
    .io_pipe_phv_in_data_395(mau_2_io_pipe_phv_in_data_395),
    .io_pipe_phv_in_data_396(mau_2_io_pipe_phv_in_data_396),
    .io_pipe_phv_in_data_397(mau_2_io_pipe_phv_in_data_397),
    .io_pipe_phv_in_data_398(mau_2_io_pipe_phv_in_data_398),
    .io_pipe_phv_in_data_399(mau_2_io_pipe_phv_in_data_399),
    .io_pipe_phv_in_data_400(mau_2_io_pipe_phv_in_data_400),
    .io_pipe_phv_in_data_401(mau_2_io_pipe_phv_in_data_401),
    .io_pipe_phv_in_data_402(mau_2_io_pipe_phv_in_data_402),
    .io_pipe_phv_in_data_403(mau_2_io_pipe_phv_in_data_403),
    .io_pipe_phv_in_data_404(mau_2_io_pipe_phv_in_data_404),
    .io_pipe_phv_in_data_405(mau_2_io_pipe_phv_in_data_405),
    .io_pipe_phv_in_data_406(mau_2_io_pipe_phv_in_data_406),
    .io_pipe_phv_in_data_407(mau_2_io_pipe_phv_in_data_407),
    .io_pipe_phv_in_data_408(mau_2_io_pipe_phv_in_data_408),
    .io_pipe_phv_in_data_409(mau_2_io_pipe_phv_in_data_409),
    .io_pipe_phv_in_data_410(mau_2_io_pipe_phv_in_data_410),
    .io_pipe_phv_in_data_411(mau_2_io_pipe_phv_in_data_411),
    .io_pipe_phv_in_data_412(mau_2_io_pipe_phv_in_data_412),
    .io_pipe_phv_in_data_413(mau_2_io_pipe_phv_in_data_413),
    .io_pipe_phv_in_data_414(mau_2_io_pipe_phv_in_data_414),
    .io_pipe_phv_in_data_415(mau_2_io_pipe_phv_in_data_415),
    .io_pipe_phv_in_data_416(mau_2_io_pipe_phv_in_data_416),
    .io_pipe_phv_in_data_417(mau_2_io_pipe_phv_in_data_417),
    .io_pipe_phv_in_data_418(mau_2_io_pipe_phv_in_data_418),
    .io_pipe_phv_in_data_419(mau_2_io_pipe_phv_in_data_419),
    .io_pipe_phv_in_data_420(mau_2_io_pipe_phv_in_data_420),
    .io_pipe_phv_in_data_421(mau_2_io_pipe_phv_in_data_421),
    .io_pipe_phv_in_data_422(mau_2_io_pipe_phv_in_data_422),
    .io_pipe_phv_in_data_423(mau_2_io_pipe_phv_in_data_423),
    .io_pipe_phv_in_data_424(mau_2_io_pipe_phv_in_data_424),
    .io_pipe_phv_in_data_425(mau_2_io_pipe_phv_in_data_425),
    .io_pipe_phv_in_data_426(mau_2_io_pipe_phv_in_data_426),
    .io_pipe_phv_in_data_427(mau_2_io_pipe_phv_in_data_427),
    .io_pipe_phv_in_data_428(mau_2_io_pipe_phv_in_data_428),
    .io_pipe_phv_in_data_429(mau_2_io_pipe_phv_in_data_429),
    .io_pipe_phv_in_data_430(mau_2_io_pipe_phv_in_data_430),
    .io_pipe_phv_in_data_431(mau_2_io_pipe_phv_in_data_431),
    .io_pipe_phv_in_data_432(mau_2_io_pipe_phv_in_data_432),
    .io_pipe_phv_in_data_433(mau_2_io_pipe_phv_in_data_433),
    .io_pipe_phv_in_data_434(mau_2_io_pipe_phv_in_data_434),
    .io_pipe_phv_in_data_435(mau_2_io_pipe_phv_in_data_435),
    .io_pipe_phv_in_data_436(mau_2_io_pipe_phv_in_data_436),
    .io_pipe_phv_in_data_437(mau_2_io_pipe_phv_in_data_437),
    .io_pipe_phv_in_data_438(mau_2_io_pipe_phv_in_data_438),
    .io_pipe_phv_in_data_439(mau_2_io_pipe_phv_in_data_439),
    .io_pipe_phv_in_data_440(mau_2_io_pipe_phv_in_data_440),
    .io_pipe_phv_in_data_441(mau_2_io_pipe_phv_in_data_441),
    .io_pipe_phv_in_data_442(mau_2_io_pipe_phv_in_data_442),
    .io_pipe_phv_in_data_443(mau_2_io_pipe_phv_in_data_443),
    .io_pipe_phv_in_data_444(mau_2_io_pipe_phv_in_data_444),
    .io_pipe_phv_in_data_445(mau_2_io_pipe_phv_in_data_445),
    .io_pipe_phv_in_data_446(mau_2_io_pipe_phv_in_data_446),
    .io_pipe_phv_in_data_447(mau_2_io_pipe_phv_in_data_447),
    .io_pipe_phv_in_data_448(mau_2_io_pipe_phv_in_data_448),
    .io_pipe_phv_in_data_449(mau_2_io_pipe_phv_in_data_449),
    .io_pipe_phv_in_data_450(mau_2_io_pipe_phv_in_data_450),
    .io_pipe_phv_in_data_451(mau_2_io_pipe_phv_in_data_451),
    .io_pipe_phv_in_data_452(mau_2_io_pipe_phv_in_data_452),
    .io_pipe_phv_in_data_453(mau_2_io_pipe_phv_in_data_453),
    .io_pipe_phv_in_data_454(mau_2_io_pipe_phv_in_data_454),
    .io_pipe_phv_in_data_455(mau_2_io_pipe_phv_in_data_455),
    .io_pipe_phv_in_data_456(mau_2_io_pipe_phv_in_data_456),
    .io_pipe_phv_in_data_457(mau_2_io_pipe_phv_in_data_457),
    .io_pipe_phv_in_data_458(mau_2_io_pipe_phv_in_data_458),
    .io_pipe_phv_in_data_459(mau_2_io_pipe_phv_in_data_459),
    .io_pipe_phv_in_data_460(mau_2_io_pipe_phv_in_data_460),
    .io_pipe_phv_in_data_461(mau_2_io_pipe_phv_in_data_461),
    .io_pipe_phv_in_data_462(mau_2_io_pipe_phv_in_data_462),
    .io_pipe_phv_in_data_463(mau_2_io_pipe_phv_in_data_463),
    .io_pipe_phv_in_data_464(mau_2_io_pipe_phv_in_data_464),
    .io_pipe_phv_in_data_465(mau_2_io_pipe_phv_in_data_465),
    .io_pipe_phv_in_data_466(mau_2_io_pipe_phv_in_data_466),
    .io_pipe_phv_in_data_467(mau_2_io_pipe_phv_in_data_467),
    .io_pipe_phv_in_data_468(mau_2_io_pipe_phv_in_data_468),
    .io_pipe_phv_in_data_469(mau_2_io_pipe_phv_in_data_469),
    .io_pipe_phv_in_data_470(mau_2_io_pipe_phv_in_data_470),
    .io_pipe_phv_in_data_471(mau_2_io_pipe_phv_in_data_471),
    .io_pipe_phv_in_data_472(mau_2_io_pipe_phv_in_data_472),
    .io_pipe_phv_in_data_473(mau_2_io_pipe_phv_in_data_473),
    .io_pipe_phv_in_data_474(mau_2_io_pipe_phv_in_data_474),
    .io_pipe_phv_in_data_475(mau_2_io_pipe_phv_in_data_475),
    .io_pipe_phv_in_data_476(mau_2_io_pipe_phv_in_data_476),
    .io_pipe_phv_in_data_477(mau_2_io_pipe_phv_in_data_477),
    .io_pipe_phv_in_data_478(mau_2_io_pipe_phv_in_data_478),
    .io_pipe_phv_in_data_479(mau_2_io_pipe_phv_in_data_479),
    .io_pipe_phv_in_data_480(mau_2_io_pipe_phv_in_data_480),
    .io_pipe_phv_in_data_481(mau_2_io_pipe_phv_in_data_481),
    .io_pipe_phv_in_data_482(mau_2_io_pipe_phv_in_data_482),
    .io_pipe_phv_in_data_483(mau_2_io_pipe_phv_in_data_483),
    .io_pipe_phv_in_data_484(mau_2_io_pipe_phv_in_data_484),
    .io_pipe_phv_in_data_485(mau_2_io_pipe_phv_in_data_485),
    .io_pipe_phv_in_data_486(mau_2_io_pipe_phv_in_data_486),
    .io_pipe_phv_in_data_487(mau_2_io_pipe_phv_in_data_487),
    .io_pipe_phv_in_data_488(mau_2_io_pipe_phv_in_data_488),
    .io_pipe_phv_in_data_489(mau_2_io_pipe_phv_in_data_489),
    .io_pipe_phv_in_data_490(mau_2_io_pipe_phv_in_data_490),
    .io_pipe_phv_in_data_491(mau_2_io_pipe_phv_in_data_491),
    .io_pipe_phv_in_data_492(mau_2_io_pipe_phv_in_data_492),
    .io_pipe_phv_in_data_493(mau_2_io_pipe_phv_in_data_493),
    .io_pipe_phv_in_data_494(mau_2_io_pipe_phv_in_data_494),
    .io_pipe_phv_in_data_495(mau_2_io_pipe_phv_in_data_495),
    .io_pipe_phv_in_data_496(mau_2_io_pipe_phv_in_data_496),
    .io_pipe_phv_in_data_497(mau_2_io_pipe_phv_in_data_497),
    .io_pipe_phv_in_data_498(mau_2_io_pipe_phv_in_data_498),
    .io_pipe_phv_in_data_499(mau_2_io_pipe_phv_in_data_499),
    .io_pipe_phv_in_data_500(mau_2_io_pipe_phv_in_data_500),
    .io_pipe_phv_in_data_501(mau_2_io_pipe_phv_in_data_501),
    .io_pipe_phv_in_data_502(mau_2_io_pipe_phv_in_data_502),
    .io_pipe_phv_in_data_503(mau_2_io_pipe_phv_in_data_503),
    .io_pipe_phv_in_data_504(mau_2_io_pipe_phv_in_data_504),
    .io_pipe_phv_in_data_505(mau_2_io_pipe_phv_in_data_505),
    .io_pipe_phv_in_data_506(mau_2_io_pipe_phv_in_data_506),
    .io_pipe_phv_in_data_507(mau_2_io_pipe_phv_in_data_507),
    .io_pipe_phv_in_data_508(mau_2_io_pipe_phv_in_data_508),
    .io_pipe_phv_in_data_509(mau_2_io_pipe_phv_in_data_509),
    .io_pipe_phv_in_data_510(mau_2_io_pipe_phv_in_data_510),
    .io_pipe_phv_in_data_511(mau_2_io_pipe_phv_in_data_511),
    .io_pipe_phv_in_header_0(mau_2_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(mau_2_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(mau_2_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(mau_2_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(mau_2_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(mau_2_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(mau_2_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(mau_2_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(mau_2_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(mau_2_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(mau_2_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(mau_2_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(mau_2_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(mau_2_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(mau_2_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(mau_2_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(mau_2_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(mau_2_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(mau_2_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(mau_2_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(mau_2_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(mau_2_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(mau_2_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(mau_2_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(mau_2_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(mau_2_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(mau_2_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(mau_2_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(mau_2_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(mau_2_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(mau_2_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(mau_2_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(mau_2_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(mau_2_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(mau_2_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(mau_2_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(mau_2_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(mau_2_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(mau_2_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(mau_2_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(mau_2_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(mau_2_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(mau_2_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(mau_2_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(mau_2_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(mau_2_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(mau_2_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(mau_2_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(mau_2_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(mau_2_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(mau_2_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(mau_2_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(mau_2_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(mau_2_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(mau_2_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(mau_2_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(mau_2_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(mau_2_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(mau_2_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(mau_2_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(mau_2_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(mau_2_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(mau_2_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(mau_2_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(mau_2_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(mau_2_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(mau_2_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(mau_2_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(mau_2_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(mau_2_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(mau_2_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(mau_2_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(mau_2_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(mau_2_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(mau_2_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(mau_2_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(mau_2_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(mau_2_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(mau_2_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(mau_2_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(mau_2_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(mau_2_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(mau_2_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(mau_2_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(mau_2_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(mau_2_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(mau_2_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(mau_2_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(mau_2_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(mau_2_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(mau_2_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(mau_2_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(mau_2_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(mau_2_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(mau_2_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(mau_2_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(mau_2_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(mau_2_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(mau_2_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(mau_2_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(mau_2_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(mau_2_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(mau_2_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(mau_2_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(mau_2_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(mau_2_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(mau_2_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(mau_2_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(mau_2_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(mau_2_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(mau_2_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(mau_2_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(mau_2_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(mau_2_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(mau_2_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(mau_2_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(mau_2_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(mau_2_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(mau_2_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(mau_2_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(mau_2_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(mau_2_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(mau_2_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(mau_2_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(mau_2_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(mau_2_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(mau_2_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(mau_2_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(mau_2_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(mau_2_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(mau_2_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(mau_2_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(mau_2_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(mau_2_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(mau_2_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(mau_2_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(mau_2_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(mau_2_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(mau_2_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(mau_2_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(mau_2_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(mau_2_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(mau_2_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(mau_2_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(mau_2_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(mau_2_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(mau_2_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(mau_2_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(mau_2_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(mau_2_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(mau_2_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(mau_2_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(mau_2_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(mau_2_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(mau_2_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(mau_2_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(mau_2_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(mau_2_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(mau_2_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(mau_2_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(mau_2_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(mau_2_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(mau_2_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(mau_2_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(mau_2_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(mau_2_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(mau_2_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(mau_2_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(mau_2_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(mau_2_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(mau_2_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(mau_2_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(mau_2_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(mau_2_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(mau_2_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(mau_2_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(mau_2_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(mau_2_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(mau_2_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(mau_2_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(mau_2_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(mau_2_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(mau_2_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(mau_2_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(mau_2_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(mau_2_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(mau_2_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(mau_2_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(mau_2_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(mau_2_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(mau_2_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(mau_2_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(mau_2_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(mau_2_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(mau_2_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(mau_2_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(mau_2_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(mau_2_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(mau_2_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(mau_2_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(mau_2_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(mau_2_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(mau_2_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(mau_2_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(mau_2_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(mau_2_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(mau_2_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(mau_2_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(mau_2_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(mau_2_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(mau_2_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(mau_2_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(mau_2_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(mau_2_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(mau_2_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(mau_2_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(mau_2_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(mau_2_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(mau_2_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(mau_2_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(mau_2_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(mau_2_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(mau_2_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(mau_2_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(mau_2_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(mau_2_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(mau_2_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(mau_2_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(mau_2_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(mau_2_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(mau_2_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(mau_2_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(mau_2_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(mau_2_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(mau_2_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(mau_2_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(mau_2_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(mau_2_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(mau_2_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(mau_2_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(mau_2_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(mau_2_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(mau_2_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(mau_2_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(mau_2_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(mau_2_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(mau_2_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(mau_2_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(mau_2_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(mau_2_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(mau_2_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(mau_2_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(mau_2_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(mau_2_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(mau_2_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(mau_2_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(mau_2_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(mau_2_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(mau_2_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(mau_2_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(mau_2_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(mau_2_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(mau_2_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(mau_2_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(mau_2_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(mau_2_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(mau_2_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(mau_2_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(mau_2_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(mau_2_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(mau_2_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(mau_2_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(mau_2_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(mau_2_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(mau_2_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(mau_2_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(mau_2_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(mau_2_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_data_256(mau_2_io_pipe_phv_out_data_256),
    .io_pipe_phv_out_data_257(mau_2_io_pipe_phv_out_data_257),
    .io_pipe_phv_out_data_258(mau_2_io_pipe_phv_out_data_258),
    .io_pipe_phv_out_data_259(mau_2_io_pipe_phv_out_data_259),
    .io_pipe_phv_out_data_260(mau_2_io_pipe_phv_out_data_260),
    .io_pipe_phv_out_data_261(mau_2_io_pipe_phv_out_data_261),
    .io_pipe_phv_out_data_262(mau_2_io_pipe_phv_out_data_262),
    .io_pipe_phv_out_data_263(mau_2_io_pipe_phv_out_data_263),
    .io_pipe_phv_out_data_264(mau_2_io_pipe_phv_out_data_264),
    .io_pipe_phv_out_data_265(mau_2_io_pipe_phv_out_data_265),
    .io_pipe_phv_out_data_266(mau_2_io_pipe_phv_out_data_266),
    .io_pipe_phv_out_data_267(mau_2_io_pipe_phv_out_data_267),
    .io_pipe_phv_out_data_268(mau_2_io_pipe_phv_out_data_268),
    .io_pipe_phv_out_data_269(mau_2_io_pipe_phv_out_data_269),
    .io_pipe_phv_out_data_270(mau_2_io_pipe_phv_out_data_270),
    .io_pipe_phv_out_data_271(mau_2_io_pipe_phv_out_data_271),
    .io_pipe_phv_out_data_272(mau_2_io_pipe_phv_out_data_272),
    .io_pipe_phv_out_data_273(mau_2_io_pipe_phv_out_data_273),
    .io_pipe_phv_out_data_274(mau_2_io_pipe_phv_out_data_274),
    .io_pipe_phv_out_data_275(mau_2_io_pipe_phv_out_data_275),
    .io_pipe_phv_out_data_276(mau_2_io_pipe_phv_out_data_276),
    .io_pipe_phv_out_data_277(mau_2_io_pipe_phv_out_data_277),
    .io_pipe_phv_out_data_278(mau_2_io_pipe_phv_out_data_278),
    .io_pipe_phv_out_data_279(mau_2_io_pipe_phv_out_data_279),
    .io_pipe_phv_out_data_280(mau_2_io_pipe_phv_out_data_280),
    .io_pipe_phv_out_data_281(mau_2_io_pipe_phv_out_data_281),
    .io_pipe_phv_out_data_282(mau_2_io_pipe_phv_out_data_282),
    .io_pipe_phv_out_data_283(mau_2_io_pipe_phv_out_data_283),
    .io_pipe_phv_out_data_284(mau_2_io_pipe_phv_out_data_284),
    .io_pipe_phv_out_data_285(mau_2_io_pipe_phv_out_data_285),
    .io_pipe_phv_out_data_286(mau_2_io_pipe_phv_out_data_286),
    .io_pipe_phv_out_data_287(mau_2_io_pipe_phv_out_data_287),
    .io_pipe_phv_out_data_288(mau_2_io_pipe_phv_out_data_288),
    .io_pipe_phv_out_data_289(mau_2_io_pipe_phv_out_data_289),
    .io_pipe_phv_out_data_290(mau_2_io_pipe_phv_out_data_290),
    .io_pipe_phv_out_data_291(mau_2_io_pipe_phv_out_data_291),
    .io_pipe_phv_out_data_292(mau_2_io_pipe_phv_out_data_292),
    .io_pipe_phv_out_data_293(mau_2_io_pipe_phv_out_data_293),
    .io_pipe_phv_out_data_294(mau_2_io_pipe_phv_out_data_294),
    .io_pipe_phv_out_data_295(mau_2_io_pipe_phv_out_data_295),
    .io_pipe_phv_out_data_296(mau_2_io_pipe_phv_out_data_296),
    .io_pipe_phv_out_data_297(mau_2_io_pipe_phv_out_data_297),
    .io_pipe_phv_out_data_298(mau_2_io_pipe_phv_out_data_298),
    .io_pipe_phv_out_data_299(mau_2_io_pipe_phv_out_data_299),
    .io_pipe_phv_out_data_300(mau_2_io_pipe_phv_out_data_300),
    .io_pipe_phv_out_data_301(mau_2_io_pipe_phv_out_data_301),
    .io_pipe_phv_out_data_302(mau_2_io_pipe_phv_out_data_302),
    .io_pipe_phv_out_data_303(mau_2_io_pipe_phv_out_data_303),
    .io_pipe_phv_out_data_304(mau_2_io_pipe_phv_out_data_304),
    .io_pipe_phv_out_data_305(mau_2_io_pipe_phv_out_data_305),
    .io_pipe_phv_out_data_306(mau_2_io_pipe_phv_out_data_306),
    .io_pipe_phv_out_data_307(mau_2_io_pipe_phv_out_data_307),
    .io_pipe_phv_out_data_308(mau_2_io_pipe_phv_out_data_308),
    .io_pipe_phv_out_data_309(mau_2_io_pipe_phv_out_data_309),
    .io_pipe_phv_out_data_310(mau_2_io_pipe_phv_out_data_310),
    .io_pipe_phv_out_data_311(mau_2_io_pipe_phv_out_data_311),
    .io_pipe_phv_out_data_312(mau_2_io_pipe_phv_out_data_312),
    .io_pipe_phv_out_data_313(mau_2_io_pipe_phv_out_data_313),
    .io_pipe_phv_out_data_314(mau_2_io_pipe_phv_out_data_314),
    .io_pipe_phv_out_data_315(mau_2_io_pipe_phv_out_data_315),
    .io_pipe_phv_out_data_316(mau_2_io_pipe_phv_out_data_316),
    .io_pipe_phv_out_data_317(mau_2_io_pipe_phv_out_data_317),
    .io_pipe_phv_out_data_318(mau_2_io_pipe_phv_out_data_318),
    .io_pipe_phv_out_data_319(mau_2_io_pipe_phv_out_data_319),
    .io_pipe_phv_out_data_320(mau_2_io_pipe_phv_out_data_320),
    .io_pipe_phv_out_data_321(mau_2_io_pipe_phv_out_data_321),
    .io_pipe_phv_out_data_322(mau_2_io_pipe_phv_out_data_322),
    .io_pipe_phv_out_data_323(mau_2_io_pipe_phv_out_data_323),
    .io_pipe_phv_out_data_324(mau_2_io_pipe_phv_out_data_324),
    .io_pipe_phv_out_data_325(mau_2_io_pipe_phv_out_data_325),
    .io_pipe_phv_out_data_326(mau_2_io_pipe_phv_out_data_326),
    .io_pipe_phv_out_data_327(mau_2_io_pipe_phv_out_data_327),
    .io_pipe_phv_out_data_328(mau_2_io_pipe_phv_out_data_328),
    .io_pipe_phv_out_data_329(mau_2_io_pipe_phv_out_data_329),
    .io_pipe_phv_out_data_330(mau_2_io_pipe_phv_out_data_330),
    .io_pipe_phv_out_data_331(mau_2_io_pipe_phv_out_data_331),
    .io_pipe_phv_out_data_332(mau_2_io_pipe_phv_out_data_332),
    .io_pipe_phv_out_data_333(mau_2_io_pipe_phv_out_data_333),
    .io_pipe_phv_out_data_334(mau_2_io_pipe_phv_out_data_334),
    .io_pipe_phv_out_data_335(mau_2_io_pipe_phv_out_data_335),
    .io_pipe_phv_out_data_336(mau_2_io_pipe_phv_out_data_336),
    .io_pipe_phv_out_data_337(mau_2_io_pipe_phv_out_data_337),
    .io_pipe_phv_out_data_338(mau_2_io_pipe_phv_out_data_338),
    .io_pipe_phv_out_data_339(mau_2_io_pipe_phv_out_data_339),
    .io_pipe_phv_out_data_340(mau_2_io_pipe_phv_out_data_340),
    .io_pipe_phv_out_data_341(mau_2_io_pipe_phv_out_data_341),
    .io_pipe_phv_out_data_342(mau_2_io_pipe_phv_out_data_342),
    .io_pipe_phv_out_data_343(mau_2_io_pipe_phv_out_data_343),
    .io_pipe_phv_out_data_344(mau_2_io_pipe_phv_out_data_344),
    .io_pipe_phv_out_data_345(mau_2_io_pipe_phv_out_data_345),
    .io_pipe_phv_out_data_346(mau_2_io_pipe_phv_out_data_346),
    .io_pipe_phv_out_data_347(mau_2_io_pipe_phv_out_data_347),
    .io_pipe_phv_out_data_348(mau_2_io_pipe_phv_out_data_348),
    .io_pipe_phv_out_data_349(mau_2_io_pipe_phv_out_data_349),
    .io_pipe_phv_out_data_350(mau_2_io_pipe_phv_out_data_350),
    .io_pipe_phv_out_data_351(mau_2_io_pipe_phv_out_data_351),
    .io_pipe_phv_out_data_352(mau_2_io_pipe_phv_out_data_352),
    .io_pipe_phv_out_data_353(mau_2_io_pipe_phv_out_data_353),
    .io_pipe_phv_out_data_354(mau_2_io_pipe_phv_out_data_354),
    .io_pipe_phv_out_data_355(mau_2_io_pipe_phv_out_data_355),
    .io_pipe_phv_out_data_356(mau_2_io_pipe_phv_out_data_356),
    .io_pipe_phv_out_data_357(mau_2_io_pipe_phv_out_data_357),
    .io_pipe_phv_out_data_358(mau_2_io_pipe_phv_out_data_358),
    .io_pipe_phv_out_data_359(mau_2_io_pipe_phv_out_data_359),
    .io_pipe_phv_out_data_360(mau_2_io_pipe_phv_out_data_360),
    .io_pipe_phv_out_data_361(mau_2_io_pipe_phv_out_data_361),
    .io_pipe_phv_out_data_362(mau_2_io_pipe_phv_out_data_362),
    .io_pipe_phv_out_data_363(mau_2_io_pipe_phv_out_data_363),
    .io_pipe_phv_out_data_364(mau_2_io_pipe_phv_out_data_364),
    .io_pipe_phv_out_data_365(mau_2_io_pipe_phv_out_data_365),
    .io_pipe_phv_out_data_366(mau_2_io_pipe_phv_out_data_366),
    .io_pipe_phv_out_data_367(mau_2_io_pipe_phv_out_data_367),
    .io_pipe_phv_out_data_368(mau_2_io_pipe_phv_out_data_368),
    .io_pipe_phv_out_data_369(mau_2_io_pipe_phv_out_data_369),
    .io_pipe_phv_out_data_370(mau_2_io_pipe_phv_out_data_370),
    .io_pipe_phv_out_data_371(mau_2_io_pipe_phv_out_data_371),
    .io_pipe_phv_out_data_372(mau_2_io_pipe_phv_out_data_372),
    .io_pipe_phv_out_data_373(mau_2_io_pipe_phv_out_data_373),
    .io_pipe_phv_out_data_374(mau_2_io_pipe_phv_out_data_374),
    .io_pipe_phv_out_data_375(mau_2_io_pipe_phv_out_data_375),
    .io_pipe_phv_out_data_376(mau_2_io_pipe_phv_out_data_376),
    .io_pipe_phv_out_data_377(mau_2_io_pipe_phv_out_data_377),
    .io_pipe_phv_out_data_378(mau_2_io_pipe_phv_out_data_378),
    .io_pipe_phv_out_data_379(mau_2_io_pipe_phv_out_data_379),
    .io_pipe_phv_out_data_380(mau_2_io_pipe_phv_out_data_380),
    .io_pipe_phv_out_data_381(mau_2_io_pipe_phv_out_data_381),
    .io_pipe_phv_out_data_382(mau_2_io_pipe_phv_out_data_382),
    .io_pipe_phv_out_data_383(mau_2_io_pipe_phv_out_data_383),
    .io_pipe_phv_out_data_384(mau_2_io_pipe_phv_out_data_384),
    .io_pipe_phv_out_data_385(mau_2_io_pipe_phv_out_data_385),
    .io_pipe_phv_out_data_386(mau_2_io_pipe_phv_out_data_386),
    .io_pipe_phv_out_data_387(mau_2_io_pipe_phv_out_data_387),
    .io_pipe_phv_out_data_388(mau_2_io_pipe_phv_out_data_388),
    .io_pipe_phv_out_data_389(mau_2_io_pipe_phv_out_data_389),
    .io_pipe_phv_out_data_390(mau_2_io_pipe_phv_out_data_390),
    .io_pipe_phv_out_data_391(mau_2_io_pipe_phv_out_data_391),
    .io_pipe_phv_out_data_392(mau_2_io_pipe_phv_out_data_392),
    .io_pipe_phv_out_data_393(mau_2_io_pipe_phv_out_data_393),
    .io_pipe_phv_out_data_394(mau_2_io_pipe_phv_out_data_394),
    .io_pipe_phv_out_data_395(mau_2_io_pipe_phv_out_data_395),
    .io_pipe_phv_out_data_396(mau_2_io_pipe_phv_out_data_396),
    .io_pipe_phv_out_data_397(mau_2_io_pipe_phv_out_data_397),
    .io_pipe_phv_out_data_398(mau_2_io_pipe_phv_out_data_398),
    .io_pipe_phv_out_data_399(mau_2_io_pipe_phv_out_data_399),
    .io_pipe_phv_out_data_400(mau_2_io_pipe_phv_out_data_400),
    .io_pipe_phv_out_data_401(mau_2_io_pipe_phv_out_data_401),
    .io_pipe_phv_out_data_402(mau_2_io_pipe_phv_out_data_402),
    .io_pipe_phv_out_data_403(mau_2_io_pipe_phv_out_data_403),
    .io_pipe_phv_out_data_404(mau_2_io_pipe_phv_out_data_404),
    .io_pipe_phv_out_data_405(mau_2_io_pipe_phv_out_data_405),
    .io_pipe_phv_out_data_406(mau_2_io_pipe_phv_out_data_406),
    .io_pipe_phv_out_data_407(mau_2_io_pipe_phv_out_data_407),
    .io_pipe_phv_out_data_408(mau_2_io_pipe_phv_out_data_408),
    .io_pipe_phv_out_data_409(mau_2_io_pipe_phv_out_data_409),
    .io_pipe_phv_out_data_410(mau_2_io_pipe_phv_out_data_410),
    .io_pipe_phv_out_data_411(mau_2_io_pipe_phv_out_data_411),
    .io_pipe_phv_out_data_412(mau_2_io_pipe_phv_out_data_412),
    .io_pipe_phv_out_data_413(mau_2_io_pipe_phv_out_data_413),
    .io_pipe_phv_out_data_414(mau_2_io_pipe_phv_out_data_414),
    .io_pipe_phv_out_data_415(mau_2_io_pipe_phv_out_data_415),
    .io_pipe_phv_out_data_416(mau_2_io_pipe_phv_out_data_416),
    .io_pipe_phv_out_data_417(mau_2_io_pipe_phv_out_data_417),
    .io_pipe_phv_out_data_418(mau_2_io_pipe_phv_out_data_418),
    .io_pipe_phv_out_data_419(mau_2_io_pipe_phv_out_data_419),
    .io_pipe_phv_out_data_420(mau_2_io_pipe_phv_out_data_420),
    .io_pipe_phv_out_data_421(mau_2_io_pipe_phv_out_data_421),
    .io_pipe_phv_out_data_422(mau_2_io_pipe_phv_out_data_422),
    .io_pipe_phv_out_data_423(mau_2_io_pipe_phv_out_data_423),
    .io_pipe_phv_out_data_424(mau_2_io_pipe_phv_out_data_424),
    .io_pipe_phv_out_data_425(mau_2_io_pipe_phv_out_data_425),
    .io_pipe_phv_out_data_426(mau_2_io_pipe_phv_out_data_426),
    .io_pipe_phv_out_data_427(mau_2_io_pipe_phv_out_data_427),
    .io_pipe_phv_out_data_428(mau_2_io_pipe_phv_out_data_428),
    .io_pipe_phv_out_data_429(mau_2_io_pipe_phv_out_data_429),
    .io_pipe_phv_out_data_430(mau_2_io_pipe_phv_out_data_430),
    .io_pipe_phv_out_data_431(mau_2_io_pipe_phv_out_data_431),
    .io_pipe_phv_out_data_432(mau_2_io_pipe_phv_out_data_432),
    .io_pipe_phv_out_data_433(mau_2_io_pipe_phv_out_data_433),
    .io_pipe_phv_out_data_434(mau_2_io_pipe_phv_out_data_434),
    .io_pipe_phv_out_data_435(mau_2_io_pipe_phv_out_data_435),
    .io_pipe_phv_out_data_436(mau_2_io_pipe_phv_out_data_436),
    .io_pipe_phv_out_data_437(mau_2_io_pipe_phv_out_data_437),
    .io_pipe_phv_out_data_438(mau_2_io_pipe_phv_out_data_438),
    .io_pipe_phv_out_data_439(mau_2_io_pipe_phv_out_data_439),
    .io_pipe_phv_out_data_440(mau_2_io_pipe_phv_out_data_440),
    .io_pipe_phv_out_data_441(mau_2_io_pipe_phv_out_data_441),
    .io_pipe_phv_out_data_442(mau_2_io_pipe_phv_out_data_442),
    .io_pipe_phv_out_data_443(mau_2_io_pipe_phv_out_data_443),
    .io_pipe_phv_out_data_444(mau_2_io_pipe_phv_out_data_444),
    .io_pipe_phv_out_data_445(mau_2_io_pipe_phv_out_data_445),
    .io_pipe_phv_out_data_446(mau_2_io_pipe_phv_out_data_446),
    .io_pipe_phv_out_data_447(mau_2_io_pipe_phv_out_data_447),
    .io_pipe_phv_out_data_448(mau_2_io_pipe_phv_out_data_448),
    .io_pipe_phv_out_data_449(mau_2_io_pipe_phv_out_data_449),
    .io_pipe_phv_out_data_450(mau_2_io_pipe_phv_out_data_450),
    .io_pipe_phv_out_data_451(mau_2_io_pipe_phv_out_data_451),
    .io_pipe_phv_out_data_452(mau_2_io_pipe_phv_out_data_452),
    .io_pipe_phv_out_data_453(mau_2_io_pipe_phv_out_data_453),
    .io_pipe_phv_out_data_454(mau_2_io_pipe_phv_out_data_454),
    .io_pipe_phv_out_data_455(mau_2_io_pipe_phv_out_data_455),
    .io_pipe_phv_out_data_456(mau_2_io_pipe_phv_out_data_456),
    .io_pipe_phv_out_data_457(mau_2_io_pipe_phv_out_data_457),
    .io_pipe_phv_out_data_458(mau_2_io_pipe_phv_out_data_458),
    .io_pipe_phv_out_data_459(mau_2_io_pipe_phv_out_data_459),
    .io_pipe_phv_out_data_460(mau_2_io_pipe_phv_out_data_460),
    .io_pipe_phv_out_data_461(mau_2_io_pipe_phv_out_data_461),
    .io_pipe_phv_out_data_462(mau_2_io_pipe_phv_out_data_462),
    .io_pipe_phv_out_data_463(mau_2_io_pipe_phv_out_data_463),
    .io_pipe_phv_out_data_464(mau_2_io_pipe_phv_out_data_464),
    .io_pipe_phv_out_data_465(mau_2_io_pipe_phv_out_data_465),
    .io_pipe_phv_out_data_466(mau_2_io_pipe_phv_out_data_466),
    .io_pipe_phv_out_data_467(mau_2_io_pipe_phv_out_data_467),
    .io_pipe_phv_out_data_468(mau_2_io_pipe_phv_out_data_468),
    .io_pipe_phv_out_data_469(mau_2_io_pipe_phv_out_data_469),
    .io_pipe_phv_out_data_470(mau_2_io_pipe_phv_out_data_470),
    .io_pipe_phv_out_data_471(mau_2_io_pipe_phv_out_data_471),
    .io_pipe_phv_out_data_472(mau_2_io_pipe_phv_out_data_472),
    .io_pipe_phv_out_data_473(mau_2_io_pipe_phv_out_data_473),
    .io_pipe_phv_out_data_474(mau_2_io_pipe_phv_out_data_474),
    .io_pipe_phv_out_data_475(mau_2_io_pipe_phv_out_data_475),
    .io_pipe_phv_out_data_476(mau_2_io_pipe_phv_out_data_476),
    .io_pipe_phv_out_data_477(mau_2_io_pipe_phv_out_data_477),
    .io_pipe_phv_out_data_478(mau_2_io_pipe_phv_out_data_478),
    .io_pipe_phv_out_data_479(mau_2_io_pipe_phv_out_data_479),
    .io_pipe_phv_out_data_480(mau_2_io_pipe_phv_out_data_480),
    .io_pipe_phv_out_data_481(mau_2_io_pipe_phv_out_data_481),
    .io_pipe_phv_out_data_482(mau_2_io_pipe_phv_out_data_482),
    .io_pipe_phv_out_data_483(mau_2_io_pipe_phv_out_data_483),
    .io_pipe_phv_out_data_484(mau_2_io_pipe_phv_out_data_484),
    .io_pipe_phv_out_data_485(mau_2_io_pipe_phv_out_data_485),
    .io_pipe_phv_out_data_486(mau_2_io_pipe_phv_out_data_486),
    .io_pipe_phv_out_data_487(mau_2_io_pipe_phv_out_data_487),
    .io_pipe_phv_out_data_488(mau_2_io_pipe_phv_out_data_488),
    .io_pipe_phv_out_data_489(mau_2_io_pipe_phv_out_data_489),
    .io_pipe_phv_out_data_490(mau_2_io_pipe_phv_out_data_490),
    .io_pipe_phv_out_data_491(mau_2_io_pipe_phv_out_data_491),
    .io_pipe_phv_out_data_492(mau_2_io_pipe_phv_out_data_492),
    .io_pipe_phv_out_data_493(mau_2_io_pipe_phv_out_data_493),
    .io_pipe_phv_out_data_494(mau_2_io_pipe_phv_out_data_494),
    .io_pipe_phv_out_data_495(mau_2_io_pipe_phv_out_data_495),
    .io_pipe_phv_out_data_496(mau_2_io_pipe_phv_out_data_496),
    .io_pipe_phv_out_data_497(mau_2_io_pipe_phv_out_data_497),
    .io_pipe_phv_out_data_498(mau_2_io_pipe_phv_out_data_498),
    .io_pipe_phv_out_data_499(mau_2_io_pipe_phv_out_data_499),
    .io_pipe_phv_out_data_500(mau_2_io_pipe_phv_out_data_500),
    .io_pipe_phv_out_data_501(mau_2_io_pipe_phv_out_data_501),
    .io_pipe_phv_out_data_502(mau_2_io_pipe_phv_out_data_502),
    .io_pipe_phv_out_data_503(mau_2_io_pipe_phv_out_data_503),
    .io_pipe_phv_out_data_504(mau_2_io_pipe_phv_out_data_504),
    .io_pipe_phv_out_data_505(mau_2_io_pipe_phv_out_data_505),
    .io_pipe_phv_out_data_506(mau_2_io_pipe_phv_out_data_506),
    .io_pipe_phv_out_data_507(mau_2_io_pipe_phv_out_data_507),
    .io_pipe_phv_out_data_508(mau_2_io_pipe_phv_out_data_508),
    .io_pipe_phv_out_data_509(mau_2_io_pipe_phv_out_data_509),
    .io_pipe_phv_out_data_510(mau_2_io_pipe_phv_out_data_510),
    .io_pipe_phv_out_data_511(mau_2_io_pipe_phv_out_data_511),
    .io_pipe_phv_out_header_0(mau_2_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(mau_2_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(mau_2_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(mau_2_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(mau_2_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(mau_2_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(mau_2_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(mau_2_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(mau_2_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(mau_2_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(mau_2_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(mau_2_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(mau_2_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(mau_2_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(mau_2_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(mau_2_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(mau_2_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(mau_2_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(mau_2_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(mau_2_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(mau_2_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(mau_2_io_pipe_phv_out_is_valid_processor),
    .io_mod_state_id_mod(mau_2_io_mod_state_id_mod),
    .io_mod_state_id(mau_2_io_mod_state_id),
    .io_mod_sram_w_cs(mau_2_io_mod_sram_w_cs),
    .io_mod_sram_w_en(mau_2_io_mod_sram_w_en),
    .io_mod_sram_w_addr(mau_2_io_mod_sram_w_addr),
    .io_mod_sram_w_data(mau_2_io_mod_sram_w_data)
  );
  ParseModule mau_3 ( // @[parser_pisa.scala 31:25]
    .clock(mau_3_clock),
    .io_pipe_phv_in_data_0(mau_3_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(mau_3_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(mau_3_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(mau_3_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(mau_3_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(mau_3_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(mau_3_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(mau_3_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(mau_3_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(mau_3_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(mau_3_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(mau_3_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(mau_3_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(mau_3_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(mau_3_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(mau_3_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(mau_3_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(mau_3_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(mau_3_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(mau_3_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(mau_3_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(mau_3_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(mau_3_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(mau_3_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(mau_3_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(mau_3_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(mau_3_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(mau_3_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(mau_3_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(mau_3_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(mau_3_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(mau_3_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(mau_3_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(mau_3_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(mau_3_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(mau_3_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(mau_3_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(mau_3_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(mau_3_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(mau_3_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(mau_3_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(mau_3_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(mau_3_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(mau_3_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(mau_3_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(mau_3_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(mau_3_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(mau_3_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(mau_3_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(mau_3_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(mau_3_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(mau_3_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(mau_3_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(mau_3_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(mau_3_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(mau_3_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(mau_3_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(mau_3_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(mau_3_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(mau_3_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(mau_3_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(mau_3_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(mau_3_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(mau_3_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(mau_3_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(mau_3_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(mau_3_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(mau_3_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(mau_3_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(mau_3_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(mau_3_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(mau_3_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(mau_3_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(mau_3_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(mau_3_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(mau_3_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(mau_3_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(mau_3_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(mau_3_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(mau_3_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(mau_3_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(mau_3_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(mau_3_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(mau_3_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(mau_3_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(mau_3_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(mau_3_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(mau_3_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(mau_3_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(mau_3_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(mau_3_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(mau_3_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(mau_3_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(mau_3_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(mau_3_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(mau_3_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(mau_3_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(mau_3_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(mau_3_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(mau_3_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(mau_3_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(mau_3_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(mau_3_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(mau_3_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(mau_3_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(mau_3_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(mau_3_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(mau_3_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(mau_3_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(mau_3_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(mau_3_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(mau_3_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(mau_3_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(mau_3_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(mau_3_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(mau_3_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(mau_3_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(mau_3_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(mau_3_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(mau_3_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(mau_3_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(mau_3_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(mau_3_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(mau_3_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(mau_3_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(mau_3_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(mau_3_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(mau_3_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(mau_3_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(mau_3_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(mau_3_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(mau_3_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(mau_3_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(mau_3_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(mau_3_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(mau_3_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(mau_3_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(mau_3_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(mau_3_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(mau_3_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(mau_3_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(mau_3_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(mau_3_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(mau_3_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(mau_3_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(mau_3_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(mau_3_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(mau_3_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(mau_3_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(mau_3_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(mau_3_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(mau_3_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(mau_3_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(mau_3_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(mau_3_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(mau_3_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(mau_3_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(mau_3_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(mau_3_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(mau_3_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(mau_3_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(mau_3_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(mau_3_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(mau_3_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(mau_3_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(mau_3_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(mau_3_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(mau_3_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(mau_3_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(mau_3_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(mau_3_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(mau_3_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(mau_3_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(mau_3_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(mau_3_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(mau_3_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(mau_3_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(mau_3_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(mau_3_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(mau_3_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(mau_3_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(mau_3_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(mau_3_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(mau_3_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(mau_3_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(mau_3_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(mau_3_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(mau_3_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(mau_3_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(mau_3_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(mau_3_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(mau_3_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(mau_3_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(mau_3_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(mau_3_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(mau_3_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(mau_3_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(mau_3_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(mau_3_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(mau_3_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(mau_3_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(mau_3_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(mau_3_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(mau_3_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(mau_3_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(mau_3_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(mau_3_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(mau_3_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(mau_3_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(mau_3_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(mau_3_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(mau_3_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(mau_3_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(mau_3_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(mau_3_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(mau_3_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(mau_3_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(mau_3_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(mau_3_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(mau_3_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(mau_3_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(mau_3_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(mau_3_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(mau_3_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(mau_3_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(mau_3_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(mau_3_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(mau_3_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(mau_3_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(mau_3_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(mau_3_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(mau_3_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(mau_3_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(mau_3_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(mau_3_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(mau_3_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(mau_3_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(mau_3_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(mau_3_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(mau_3_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(mau_3_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(mau_3_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(mau_3_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(mau_3_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(mau_3_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(mau_3_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(mau_3_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(mau_3_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(mau_3_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(mau_3_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(mau_3_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(mau_3_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(mau_3_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(mau_3_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(mau_3_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(mau_3_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_data_256(mau_3_io_pipe_phv_in_data_256),
    .io_pipe_phv_in_data_257(mau_3_io_pipe_phv_in_data_257),
    .io_pipe_phv_in_data_258(mau_3_io_pipe_phv_in_data_258),
    .io_pipe_phv_in_data_259(mau_3_io_pipe_phv_in_data_259),
    .io_pipe_phv_in_data_260(mau_3_io_pipe_phv_in_data_260),
    .io_pipe_phv_in_data_261(mau_3_io_pipe_phv_in_data_261),
    .io_pipe_phv_in_data_262(mau_3_io_pipe_phv_in_data_262),
    .io_pipe_phv_in_data_263(mau_3_io_pipe_phv_in_data_263),
    .io_pipe_phv_in_data_264(mau_3_io_pipe_phv_in_data_264),
    .io_pipe_phv_in_data_265(mau_3_io_pipe_phv_in_data_265),
    .io_pipe_phv_in_data_266(mau_3_io_pipe_phv_in_data_266),
    .io_pipe_phv_in_data_267(mau_3_io_pipe_phv_in_data_267),
    .io_pipe_phv_in_data_268(mau_3_io_pipe_phv_in_data_268),
    .io_pipe_phv_in_data_269(mau_3_io_pipe_phv_in_data_269),
    .io_pipe_phv_in_data_270(mau_3_io_pipe_phv_in_data_270),
    .io_pipe_phv_in_data_271(mau_3_io_pipe_phv_in_data_271),
    .io_pipe_phv_in_data_272(mau_3_io_pipe_phv_in_data_272),
    .io_pipe_phv_in_data_273(mau_3_io_pipe_phv_in_data_273),
    .io_pipe_phv_in_data_274(mau_3_io_pipe_phv_in_data_274),
    .io_pipe_phv_in_data_275(mau_3_io_pipe_phv_in_data_275),
    .io_pipe_phv_in_data_276(mau_3_io_pipe_phv_in_data_276),
    .io_pipe_phv_in_data_277(mau_3_io_pipe_phv_in_data_277),
    .io_pipe_phv_in_data_278(mau_3_io_pipe_phv_in_data_278),
    .io_pipe_phv_in_data_279(mau_3_io_pipe_phv_in_data_279),
    .io_pipe_phv_in_data_280(mau_3_io_pipe_phv_in_data_280),
    .io_pipe_phv_in_data_281(mau_3_io_pipe_phv_in_data_281),
    .io_pipe_phv_in_data_282(mau_3_io_pipe_phv_in_data_282),
    .io_pipe_phv_in_data_283(mau_3_io_pipe_phv_in_data_283),
    .io_pipe_phv_in_data_284(mau_3_io_pipe_phv_in_data_284),
    .io_pipe_phv_in_data_285(mau_3_io_pipe_phv_in_data_285),
    .io_pipe_phv_in_data_286(mau_3_io_pipe_phv_in_data_286),
    .io_pipe_phv_in_data_287(mau_3_io_pipe_phv_in_data_287),
    .io_pipe_phv_in_data_288(mau_3_io_pipe_phv_in_data_288),
    .io_pipe_phv_in_data_289(mau_3_io_pipe_phv_in_data_289),
    .io_pipe_phv_in_data_290(mau_3_io_pipe_phv_in_data_290),
    .io_pipe_phv_in_data_291(mau_3_io_pipe_phv_in_data_291),
    .io_pipe_phv_in_data_292(mau_3_io_pipe_phv_in_data_292),
    .io_pipe_phv_in_data_293(mau_3_io_pipe_phv_in_data_293),
    .io_pipe_phv_in_data_294(mau_3_io_pipe_phv_in_data_294),
    .io_pipe_phv_in_data_295(mau_3_io_pipe_phv_in_data_295),
    .io_pipe_phv_in_data_296(mau_3_io_pipe_phv_in_data_296),
    .io_pipe_phv_in_data_297(mau_3_io_pipe_phv_in_data_297),
    .io_pipe_phv_in_data_298(mau_3_io_pipe_phv_in_data_298),
    .io_pipe_phv_in_data_299(mau_3_io_pipe_phv_in_data_299),
    .io_pipe_phv_in_data_300(mau_3_io_pipe_phv_in_data_300),
    .io_pipe_phv_in_data_301(mau_3_io_pipe_phv_in_data_301),
    .io_pipe_phv_in_data_302(mau_3_io_pipe_phv_in_data_302),
    .io_pipe_phv_in_data_303(mau_3_io_pipe_phv_in_data_303),
    .io_pipe_phv_in_data_304(mau_3_io_pipe_phv_in_data_304),
    .io_pipe_phv_in_data_305(mau_3_io_pipe_phv_in_data_305),
    .io_pipe_phv_in_data_306(mau_3_io_pipe_phv_in_data_306),
    .io_pipe_phv_in_data_307(mau_3_io_pipe_phv_in_data_307),
    .io_pipe_phv_in_data_308(mau_3_io_pipe_phv_in_data_308),
    .io_pipe_phv_in_data_309(mau_3_io_pipe_phv_in_data_309),
    .io_pipe_phv_in_data_310(mau_3_io_pipe_phv_in_data_310),
    .io_pipe_phv_in_data_311(mau_3_io_pipe_phv_in_data_311),
    .io_pipe_phv_in_data_312(mau_3_io_pipe_phv_in_data_312),
    .io_pipe_phv_in_data_313(mau_3_io_pipe_phv_in_data_313),
    .io_pipe_phv_in_data_314(mau_3_io_pipe_phv_in_data_314),
    .io_pipe_phv_in_data_315(mau_3_io_pipe_phv_in_data_315),
    .io_pipe_phv_in_data_316(mau_3_io_pipe_phv_in_data_316),
    .io_pipe_phv_in_data_317(mau_3_io_pipe_phv_in_data_317),
    .io_pipe_phv_in_data_318(mau_3_io_pipe_phv_in_data_318),
    .io_pipe_phv_in_data_319(mau_3_io_pipe_phv_in_data_319),
    .io_pipe_phv_in_data_320(mau_3_io_pipe_phv_in_data_320),
    .io_pipe_phv_in_data_321(mau_3_io_pipe_phv_in_data_321),
    .io_pipe_phv_in_data_322(mau_3_io_pipe_phv_in_data_322),
    .io_pipe_phv_in_data_323(mau_3_io_pipe_phv_in_data_323),
    .io_pipe_phv_in_data_324(mau_3_io_pipe_phv_in_data_324),
    .io_pipe_phv_in_data_325(mau_3_io_pipe_phv_in_data_325),
    .io_pipe_phv_in_data_326(mau_3_io_pipe_phv_in_data_326),
    .io_pipe_phv_in_data_327(mau_3_io_pipe_phv_in_data_327),
    .io_pipe_phv_in_data_328(mau_3_io_pipe_phv_in_data_328),
    .io_pipe_phv_in_data_329(mau_3_io_pipe_phv_in_data_329),
    .io_pipe_phv_in_data_330(mau_3_io_pipe_phv_in_data_330),
    .io_pipe_phv_in_data_331(mau_3_io_pipe_phv_in_data_331),
    .io_pipe_phv_in_data_332(mau_3_io_pipe_phv_in_data_332),
    .io_pipe_phv_in_data_333(mau_3_io_pipe_phv_in_data_333),
    .io_pipe_phv_in_data_334(mau_3_io_pipe_phv_in_data_334),
    .io_pipe_phv_in_data_335(mau_3_io_pipe_phv_in_data_335),
    .io_pipe_phv_in_data_336(mau_3_io_pipe_phv_in_data_336),
    .io_pipe_phv_in_data_337(mau_3_io_pipe_phv_in_data_337),
    .io_pipe_phv_in_data_338(mau_3_io_pipe_phv_in_data_338),
    .io_pipe_phv_in_data_339(mau_3_io_pipe_phv_in_data_339),
    .io_pipe_phv_in_data_340(mau_3_io_pipe_phv_in_data_340),
    .io_pipe_phv_in_data_341(mau_3_io_pipe_phv_in_data_341),
    .io_pipe_phv_in_data_342(mau_3_io_pipe_phv_in_data_342),
    .io_pipe_phv_in_data_343(mau_3_io_pipe_phv_in_data_343),
    .io_pipe_phv_in_data_344(mau_3_io_pipe_phv_in_data_344),
    .io_pipe_phv_in_data_345(mau_3_io_pipe_phv_in_data_345),
    .io_pipe_phv_in_data_346(mau_3_io_pipe_phv_in_data_346),
    .io_pipe_phv_in_data_347(mau_3_io_pipe_phv_in_data_347),
    .io_pipe_phv_in_data_348(mau_3_io_pipe_phv_in_data_348),
    .io_pipe_phv_in_data_349(mau_3_io_pipe_phv_in_data_349),
    .io_pipe_phv_in_data_350(mau_3_io_pipe_phv_in_data_350),
    .io_pipe_phv_in_data_351(mau_3_io_pipe_phv_in_data_351),
    .io_pipe_phv_in_data_352(mau_3_io_pipe_phv_in_data_352),
    .io_pipe_phv_in_data_353(mau_3_io_pipe_phv_in_data_353),
    .io_pipe_phv_in_data_354(mau_3_io_pipe_phv_in_data_354),
    .io_pipe_phv_in_data_355(mau_3_io_pipe_phv_in_data_355),
    .io_pipe_phv_in_data_356(mau_3_io_pipe_phv_in_data_356),
    .io_pipe_phv_in_data_357(mau_3_io_pipe_phv_in_data_357),
    .io_pipe_phv_in_data_358(mau_3_io_pipe_phv_in_data_358),
    .io_pipe_phv_in_data_359(mau_3_io_pipe_phv_in_data_359),
    .io_pipe_phv_in_data_360(mau_3_io_pipe_phv_in_data_360),
    .io_pipe_phv_in_data_361(mau_3_io_pipe_phv_in_data_361),
    .io_pipe_phv_in_data_362(mau_3_io_pipe_phv_in_data_362),
    .io_pipe_phv_in_data_363(mau_3_io_pipe_phv_in_data_363),
    .io_pipe_phv_in_data_364(mau_3_io_pipe_phv_in_data_364),
    .io_pipe_phv_in_data_365(mau_3_io_pipe_phv_in_data_365),
    .io_pipe_phv_in_data_366(mau_3_io_pipe_phv_in_data_366),
    .io_pipe_phv_in_data_367(mau_3_io_pipe_phv_in_data_367),
    .io_pipe_phv_in_data_368(mau_3_io_pipe_phv_in_data_368),
    .io_pipe_phv_in_data_369(mau_3_io_pipe_phv_in_data_369),
    .io_pipe_phv_in_data_370(mau_3_io_pipe_phv_in_data_370),
    .io_pipe_phv_in_data_371(mau_3_io_pipe_phv_in_data_371),
    .io_pipe_phv_in_data_372(mau_3_io_pipe_phv_in_data_372),
    .io_pipe_phv_in_data_373(mau_3_io_pipe_phv_in_data_373),
    .io_pipe_phv_in_data_374(mau_3_io_pipe_phv_in_data_374),
    .io_pipe_phv_in_data_375(mau_3_io_pipe_phv_in_data_375),
    .io_pipe_phv_in_data_376(mau_3_io_pipe_phv_in_data_376),
    .io_pipe_phv_in_data_377(mau_3_io_pipe_phv_in_data_377),
    .io_pipe_phv_in_data_378(mau_3_io_pipe_phv_in_data_378),
    .io_pipe_phv_in_data_379(mau_3_io_pipe_phv_in_data_379),
    .io_pipe_phv_in_data_380(mau_3_io_pipe_phv_in_data_380),
    .io_pipe_phv_in_data_381(mau_3_io_pipe_phv_in_data_381),
    .io_pipe_phv_in_data_382(mau_3_io_pipe_phv_in_data_382),
    .io_pipe_phv_in_data_383(mau_3_io_pipe_phv_in_data_383),
    .io_pipe_phv_in_data_384(mau_3_io_pipe_phv_in_data_384),
    .io_pipe_phv_in_data_385(mau_3_io_pipe_phv_in_data_385),
    .io_pipe_phv_in_data_386(mau_3_io_pipe_phv_in_data_386),
    .io_pipe_phv_in_data_387(mau_3_io_pipe_phv_in_data_387),
    .io_pipe_phv_in_data_388(mau_3_io_pipe_phv_in_data_388),
    .io_pipe_phv_in_data_389(mau_3_io_pipe_phv_in_data_389),
    .io_pipe_phv_in_data_390(mau_3_io_pipe_phv_in_data_390),
    .io_pipe_phv_in_data_391(mau_3_io_pipe_phv_in_data_391),
    .io_pipe_phv_in_data_392(mau_3_io_pipe_phv_in_data_392),
    .io_pipe_phv_in_data_393(mau_3_io_pipe_phv_in_data_393),
    .io_pipe_phv_in_data_394(mau_3_io_pipe_phv_in_data_394),
    .io_pipe_phv_in_data_395(mau_3_io_pipe_phv_in_data_395),
    .io_pipe_phv_in_data_396(mau_3_io_pipe_phv_in_data_396),
    .io_pipe_phv_in_data_397(mau_3_io_pipe_phv_in_data_397),
    .io_pipe_phv_in_data_398(mau_3_io_pipe_phv_in_data_398),
    .io_pipe_phv_in_data_399(mau_3_io_pipe_phv_in_data_399),
    .io_pipe_phv_in_data_400(mau_3_io_pipe_phv_in_data_400),
    .io_pipe_phv_in_data_401(mau_3_io_pipe_phv_in_data_401),
    .io_pipe_phv_in_data_402(mau_3_io_pipe_phv_in_data_402),
    .io_pipe_phv_in_data_403(mau_3_io_pipe_phv_in_data_403),
    .io_pipe_phv_in_data_404(mau_3_io_pipe_phv_in_data_404),
    .io_pipe_phv_in_data_405(mau_3_io_pipe_phv_in_data_405),
    .io_pipe_phv_in_data_406(mau_3_io_pipe_phv_in_data_406),
    .io_pipe_phv_in_data_407(mau_3_io_pipe_phv_in_data_407),
    .io_pipe_phv_in_data_408(mau_3_io_pipe_phv_in_data_408),
    .io_pipe_phv_in_data_409(mau_3_io_pipe_phv_in_data_409),
    .io_pipe_phv_in_data_410(mau_3_io_pipe_phv_in_data_410),
    .io_pipe_phv_in_data_411(mau_3_io_pipe_phv_in_data_411),
    .io_pipe_phv_in_data_412(mau_3_io_pipe_phv_in_data_412),
    .io_pipe_phv_in_data_413(mau_3_io_pipe_phv_in_data_413),
    .io_pipe_phv_in_data_414(mau_3_io_pipe_phv_in_data_414),
    .io_pipe_phv_in_data_415(mau_3_io_pipe_phv_in_data_415),
    .io_pipe_phv_in_data_416(mau_3_io_pipe_phv_in_data_416),
    .io_pipe_phv_in_data_417(mau_3_io_pipe_phv_in_data_417),
    .io_pipe_phv_in_data_418(mau_3_io_pipe_phv_in_data_418),
    .io_pipe_phv_in_data_419(mau_3_io_pipe_phv_in_data_419),
    .io_pipe_phv_in_data_420(mau_3_io_pipe_phv_in_data_420),
    .io_pipe_phv_in_data_421(mau_3_io_pipe_phv_in_data_421),
    .io_pipe_phv_in_data_422(mau_3_io_pipe_phv_in_data_422),
    .io_pipe_phv_in_data_423(mau_3_io_pipe_phv_in_data_423),
    .io_pipe_phv_in_data_424(mau_3_io_pipe_phv_in_data_424),
    .io_pipe_phv_in_data_425(mau_3_io_pipe_phv_in_data_425),
    .io_pipe_phv_in_data_426(mau_3_io_pipe_phv_in_data_426),
    .io_pipe_phv_in_data_427(mau_3_io_pipe_phv_in_data_427),
    .io_pipe_phv_in_data_428(mau_3_io_pipe_phv_in_data_428),
    .io_pipe_phv_in_data_429(mau_3_io_pipe_phv_in_data_429),
    .io_pipe_phv_in_data_430(mau_3_io_pipe_phv_in_data_430),
    .io_pipe_phv_in_data_431(mau_3_io_pipe_phv_in_data_431),
    .io_pipe_phv_in_data_432(mau_3_io_pipe_phv_in_data_432),
    .io_pipe_phv_in_data_433(mau_3_io_pipe_phv_in_data_433),
    .io_pipe_phv_in_data_434(mau_3_io_pipe_phv_in_data_434),
    .io_pipe_phv_in_data_435(mau_3_io_pipe_phv_in_data_435),
    .io_pipe_phv_in_data_436(mau_3_io_pipe_phv_in_data_436),
    .io_pipe_phv_in_data_437(mau_3_io_pipe_phv_in_data_437),
    .io_pipe_phv_in_data_438(mau_3_io_pipe_phv_in_data_438),
    .io_pipe_phv_in_data_439(mau_3_io_pipe_phv_in_data_439),
    .io_pipe_phv_in_data_440(mau_3_io_pipe_phv_in_data_440),
    .io_pipe_phv_in_data_441(mau_3_io_pipe_phv_in_data_441),
    .io_pipe_phv_in_data_442(mau_3_io_pipe_phv_in_data_442),
    .io_pipe_phv_in_data_443(mau_3_io_pipe_phv_in_data_443),
    .io_pipe_phv_in_data_444(mau_3_io_pipe_phv_in_data_444),
    .io_pipe_phv_in_data_445(mau_3_io_pipe_phv_in_data_445),
    .io_pipe_phv_in_data_446(mau_3_io_pipe_phv_in_data_446),
    .io_pipe_phv_in_data_447(mau_3_io_pipe_phv_in_data_447),
    .io_pipe_phv_in_data_448(mau_3_io_pipe_phv_in_data_448),
    .io_pipe_phv_in_data_449(mau_3_io_pipe_phv_in_data_449),
    .io_pipe_phv_in_data_450(mau_3_io_pipe_phv_in_data_450),
    .io_pipe_phv_in_data_451(mau_3_io_pipe_phv_in_data_451),
    .io_pipe_phv_in_data_452(mau_3_io_pipe_phv_in_data_452),
    .io_pipe_phv_in_data_453(mau_3_io_pipe_phv_in_data_453),
    .io_pipe_phv_in_data_454(mau_3_io_pipe_phv_in_data_454),
    .io_pipe_phv_in_data_455(mau_3_io_pipe_phv_in_data_455),
    .io_pipe_phv_in_data_456(mau_3_io_pipe_phv_in_data_456),
    .io_pipe_phv_in_data_457(mau_3_io_pipe_phv_in_data_457),
    .io_pipe_phv_in_data_458(mau_3_io_pipe_phv_in_data_458),
    .io_pipe_phv_in_data_459(mau_3_io_pipe_phv_in_data_459),
    .io_pipe_phv_in_data_460(mau_3_io_pipe_phv_in_data_460),
    .io_pipe_phv_in_data_461(mau_3_io_pipe_phv_in_data_461),
    .io_pipe_phv_in_data_462(mau_3_io_pipe_phv_in_data_462),
    .io_pipe_phv_in_data_463(mau_3_io_pipe_phv_in_data_463),
    .io_pipe_phv_in_data_464(mau_3_io_pipe_phv_in_data_464),
    .io_pipe_phv_in_data_465(mau_3_io_pipe_phv_in_data_465),
    .io_pipe_phv_in_data_466(mau_3_io_pipe_phv_in_data_466),
    .io_pipe_phv_in_data_467(mau_3_io_pipe_phv_in_data_467),
    .io_pipe_phv_in_data_468(mau_3_io_pipe_phv_in_data_468),
    .io_pipe_phv_in_data_469(mau_3_io_pipe_phv_in_data_469),
    .io_pipe_phv_in_data_470(mau_3_io_pipe_phv_in_data_470),
    .io_pipe_phv_in_data_471(mau_3_io_pipe_phv_in_data_471),
    .io_pipe_phv_in_data_472(mau_3_io_pipe_phv_in_data_472),
    .io_pipe_phv_in_data_473(mau_3_io_pipe_phv_in_data_473),
    .io_pipe_phv_in_data_474(mau_3_io_pipe_phv_in_data_474),
    .io_pipe_phv_in_data_475(mau_3_io_pipe_phv_in_data_475),
    .io_pipe_phv_in_data_476(mau_3_io_pipe_phv_in_data_476),
    .io_pipe_phv_in_data_477(mau_3_io_pipe_phv_in_data_477),
    .io_pipe_phv_in_data_478(mau_3_io_pipe_phv_in_data_478),
    .io_pipe_phv_in_data_479(mau_3_io_pipe_phv_in_data_479),
    .io_pipe_phv_in_data_480(mau_3_io_pipe_phv_in_data_480),
    .io_pipe_phv_in_data_481(mau_3_io_pipe_phv_in_data_481),
    .io_pipe_phv_in_data_482(mau_3_io_pipe_phv_in_data_482),
    .io_pipe_phv_in_data_483(mau_3_io_pipe_phv_in_data_483),
    .io_pipe_phv_in_data_484(mau_3_io_pipe_phv_in_data_484),
    .io_pipe_phv_in_data_485(mau_3_io_pipe_phv_in_data_485),
    .io_pipe_phv_in_data_486(mau_3_io_pipe_phv_in_data_486),
    .io_pipe_phv_in_data_487(mau_3_io_pipe_phv_in_data_487),
    .io_pipe_phv_in_data_488(mau_3_io_pipe_phv_in_data_488),
    .io_pipe_phv_in_data_489(mau_3_io_pipe_phv_in_data_489),
    .io_pipe_phv_in_data_490(mau_3_io_pipe_phv_in_data_490),
    .io_pipe_phv_in_data_491(mau_3_io_pipe_phv_in_data_491),
    .io_pipe_phv_in_data_492(mau_3_io_pipe_phv_in_data_492),
    .io_pipe_phv_in_data_493(mau_3_io_pipe_phv_in_data_493),
    .io_pipe_phv_in_data_494(mau_3_io_pipe_phv_in_data_494),
    .io_pipe_phv_in_data_495(mau_3_io_pipe_phv_in_data_495),
    .io_pipe_phv_in_data_496(mau_3_io_pipe_phv_in_data_496),
    .io_pipe_phv_in_data_497(mau_3_io_pipe_phv_in_data_497),
    .io_pipe_phv_in_data_498(mau_3_io_pipe_phv_in_data_498),
    .io_pipe_phv_in_data_499(mau_3_io_pipe_phv_in_data_499),
    .io_pipe_phv_in_data_500(mau_3_io_pipe_phv_in_data_500),
    .io_pipe_phv_in_data_501(mau_3_io_pipe_phv_in_data_501),
    .io_pipe_phv_in_data_502(mau_3_io_pipe_phv_in_data_502),
    .io_pipe_phv_in_data_503(mau_3_io_pipe_phv_in_data_503),
    .io_pipe_phv_in_data_504(mau_3_io_pipe_phv_in_data_504),
    .io_pipe_phv_in_data_505(mau_3_io_pipe_phv_in_data_505),
    .io_pipe_phv_in_data_506(mau_3_io_pipe_phv_in_data_506),
    .io_pipe_phv_in_data_507(mau_3_io_pipe_phv_in_data_507),
    .io_pipe_phv_in_data_508(mau_3_io_pipe_phv_in_data_508),
    .io_pipe_phv_in_data_509(mau_3_io_pipe_phv_in_data_509),
    .io_pipe_phv_in_data_510(mau_3_io_pipe_phv_in_data_510),
    .io_pipe_phv_in_data_511(mau_3_io_pipe_phv_in_data_511),
    .io_pipe_phv_in_header_0(mau_3_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(mau_3_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(mau_3_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(mau_3_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(mau_3_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(mau_3_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(mau_3_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(mau_3_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(mau_3_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(mau_3_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(mau_3_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(mau_3_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(mau_3_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(mau_3_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(mau_3_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(mau_3_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(mau_3_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(mau_3_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(mau_3_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(mau_3_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(mau_3_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(mau_3_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(mau_3_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(mau_3_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(mau_3_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(mau_3_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(mau_3_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(mau_3_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(mau_3_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(mau_3_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(mau_3_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(mau_3_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(mau_3_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(mau_3_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(mau_3_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(mau_3_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(mau_3_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(mau_3_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(mau_3_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(mau_3_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(mau_3_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(mau_3_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(mau_3_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(mau_3_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(mau_3_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(mau_3_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(mau_3_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(mau_3_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(mau_3_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(mau_3_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(mau_3_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(mau_3_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(mau_3_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(mau_3_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(mau_3_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(mau_3_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(mau_3_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(mau_3_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(mau_3_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(mau_3_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(mau_3_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(mau_3_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(mau_3_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(mau_3_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(mau_3_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(mau_3_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(mau_3_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(mau_3_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(mau_3_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(mau_3_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(mau_3_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(mau_3_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(mau_3_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(mau_3_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(mau_3_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(mau_3_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(mau_3_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(mau_3_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(mau_3_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(mau_3_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(mau_3_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(mau_3_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(mau_3_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(mau_3_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(mau_3_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(mau_3_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(mau_3_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(mau_3_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(mau_3_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(mau_3_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(mau_3_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(mau_3_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(mau_3_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(mau_3_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(mau_3_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(mau_3_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(mau_3_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(mau_3_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(mau_3_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(mau_3_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(mau_3_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(mau_3_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(mau_3_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(mau_3_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(mau_3_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(mau_3_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(mau_3_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(mau_3_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(mau_3_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(mau_3_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(mau_3_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(mau_3_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(mau_3_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(mau_3_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(mau_3_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(mau_3_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(mau_3_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(mau_3_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(mau_3_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(mau_3_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(mau_3_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(mau_3_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(mau_3_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(mau_3_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(mau_3_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(mau_3_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(mau_3_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(mau_3_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(mau_3_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(mau_3_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(mau_3_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(mau_3_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(mau_3_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(mau_3_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(mau_3_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(mau_3_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(mau_3_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(mau_3_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(mau_3_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(mau_3_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(mau_3_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(mau_3_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(mau_3_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(mau_3_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(mau_3_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(mau_3_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(mau_3_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(mau_3_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(mau_3_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(mau_3_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(mau_3_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(mau_3_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(mau_3_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(mau_3_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(mau_3_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(mau_3_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(mau_3_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(mau_3_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(mau_3_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(mau_3_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(mau_3_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(mau_3_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(mau_3_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(mau_3_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(mau_3_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(mau_3_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(mau_3_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(mau_3_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(mau_3_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(mau_3_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(mau_3_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(mau_3_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(mau_3_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(mau_3_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(mau_3_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(mau_3_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(mau_3_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(mau_3_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(mau_3_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(mau_3_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(mau_3_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(mau_3_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(mau_3_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(mau_3_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(mau_3_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(mau_3_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(mau_3_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(mau_3_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(mau_3_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(mau_3_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(mau_3_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(mau_3_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(mau_3_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(mau_3_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(mau_3_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(mau_3_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(mau_3_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(mau_3_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(mau_3_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(mau_3_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(mau_3_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(mau_3_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(mau_3_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(mau_3_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(mau_3_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(mau_3_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(mau_3_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(mau_3_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(mau_3_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(mau_3_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(mau_3_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(mau_3_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(mau_3_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(mau_3_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(mau_3_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(mau_3_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(mau_3_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(mau_3_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(mau_3_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(mau_3_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(mau_3_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(mau_3_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(mau_3_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(mau_3_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(mau_3_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(mau_3_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(mau_3_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(mau_3_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(mau_3_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(mau_3_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(mau_3_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(mau_3_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(mau_3_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(mau_3_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(mau_3_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(mau_3_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(mau_3_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(mau_3_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(mau_3_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(mau_3_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(mau_3_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(mau_3_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(mau_3_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(mau_3_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(mau_3_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(mau_3_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(mau_3_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(mau_3_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(mau_3_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(mau_3_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(mau_3_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(mau_3_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(mau_3_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(mau_3_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(mau_3_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(mau_3_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(mau_3_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(mau_3_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(mau_3_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(mau_3_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(mau_3_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(mau_3_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(mau_3_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(mau_3_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(mau_3_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(mau_3_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(mau_3_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(mau_3_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(mau_3_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(mau_3_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(mau_3_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(mau_3_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(mau_3_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(mau_3_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(mau_3_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(mau_3_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(mau_3_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(mau_3_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_data_256(mau_3_io_pipe_phv_out_data_256),
    .io_pipe_phv_out_data_257(mau_3_io_pipe_phv_out_data_257),
    .io_pipe_phv_out_data_258(mau_3_io_pipe_phv_out_data_258),
    .io_pipe_phv_out_data_259(mau_3_io_pipe_phv_out_data_259),
    .io_pipe_phv_out_data_260(mau_3_io_pipe_phv_out_data_260),
    .io_pipe_phv_out_data_261(mau_3_io_pipe_phv_out_data_261),
    .io_pipe_phv_out_data_262(mau_3_io_pipe_phv_out_data_262),
    .io_pipe_phv_out_data_263(mau_3_io_pipe_phv_out_data_263),
    .io_pipe_phv_out_data_264(mau_3_io_pipe_phv_out_data_264),
    .io_pipe_phv_out_data_265(mau_3_io_pipe_phv_out_data_265),
    .io_pipe_phv_out_data_266(mau_3_io_pipe_phv_out_data_266),
    .io_pipe_phv_out_data_267(mau_3_io_pipe_phv_out_data_267),
    .io_pipe_phv_out_data_268(mau_3_io_pipe_phv_out_data_268),
    .io_pipe_phv_out_data_269(mau_3_io_pipe_phv_out_data_269),
    .io_pipe_phv_out_data_270(mau_3_io_pipe_phv_out_data_270),
    .io_pipe_phv_out_data_271(mau_3_io_pipe_phv_out_data_271),
    .io_pipe_phv_out_data_272(mau_3_io_pipe_phv_out_data_272),
    .io_pipe_phv_out_data_273(mau_3_io_pipe_phv_out_data_273),
    .io_pipe_phv_out_data_274(mau_3_io_pipe_phv_out_data_274),
    .io_pipe_phv_out_data_275(mau_3_io_pipe_phv_out_data_275),
    .io_pipe_phv_out_data_276(mau_3_io_pipe_phv_out_data_276),
    .io_pipe_phv_out_data_277(mau_3_io_pipe_phv_out_data_277),
    .io_pipe_phv_out_data_278(mau_3_io_pipe_phv_out_data_278),
    .io_pipe_phv_out_data_279(mau_3_io_pipe_phv_out_data_279),
    .io_pipe_phv_out_data_280(mau_3_io_pipe_phv_out_data_280),
    .io_pipe_phv_out_data_281(mau_3_io_pipe_phv_out_data_281),
    .io_pipe_phv_out_data_282(mau_3_io_pipe_phv_out_data_282),
    .io_pipe_phv_out_data_283(mau_3_io_pipe_phv_out_data_283),
    .io_pipe_phv_out_data_284(mau_3_io_pipe_phv_out_data_284),
    .io_pipe_phv_out_data_285(mau_3_io_pipe_phv_out_data_285),
    .io_pipe_phv_out_data_286(mau_3_io_pipe_phv_out_data_286),
    .io_pipe_phv_out_data_287(mau_3_io_pipe_phv_out_data_287),
    .io_pipe_phv_out_data_288(mau_3_io_pipe_phv_out_data_288),
    .io_pipe_phv_out_data_289(mau_3_io_pipe_phv_out_data_289),
    .io_pipe_phv_out_data_290(mau_3_io_pipe_phv_out_data_290),
    .io_pipe_phv_out_data_291(mau_3_io_pipe_phv_out_data_291),
    .io_pipe_phv_out_data_292(mau_3_io_pipe_phv_out_data_292),
    .io_pipe_phv_out_data_293(mau_3_io_pipe_phv_out_data_293),
    .io_pipe_phv_out_data_294(mau_3_io_pipe_phv_out_data_294),
    .io_pipe_phv_out_data_295(mau_3_io_pipe_phv_out_data_295),
    .io_pipe_phv_out_data_296(mau_3_io_pipe_phv_out_data_296),
    .io_pipe_phv_out_data_297(mau_3_io_pipe_phv_out_data_297),
    .io_pipe_phv_out_data_298(mau_3_io_pipe_phv_out_data_298),
    .io_pipe_phv_out_data_299(mau_3_io_pipe_phv_out_data_299),
    .io_pipe_phv_out_data_300(mau_3_io_pipe_phv_out_data_300),
    .io_pipe_phv_out_data_301(mau_3_io_pipe_phv_out_data_301),
    .io_pipe_phv_out_data_302(mau_3_io_pipe_phv_out_data_302),
    .io_pipe_phv_out_data_303(mau_3_io_pipe_phv_out_data_303),
    .io_pipe_phv_out_data_304(mau_3_io_pipe_phv_out_data_304),
    .io_pipe_phv_out_data_305(mau_3_io_pipe_phv_out_data_305),
    .io_pipe_phv_out_data_306(mau_3_io_pipe_phv_out_data_306),
    .io_pipe_phv_out_data_307(mau_3_io_pipe_phv_out_data_307),
    .io_pipe_phv_out_data_308(mau_3_io_pipe_phv_out_data_308),
    .io_pipe_phv_out_data_309(mau_3_io_pipe_phv_out_data_309),
    .io_pipe_phv_out_data_310(mau_3_io_pipe_phv_out_data_310),
    .io_pipe_phv_out_data_311(mau_3_io_pipe_phv_out_data_311),
    .io_pipe_phv_out_data_312(mau_3_io_pipe_phv_out_data_312),
    .io_pipe_phv_out_data_313(mau_3_io_pipe_phv_out_data_313),
    .io_pipe_phv_out_data_314(mau_3_io_pipe_phv_out_data_314),
    .io_pipe_phv_out_data_315(mau_3_io_pipe_phv_out_data_315),
    .io_pipe_phv_out_data_316(mau_3_io_pipe_phv_out_data_316),
    .io_pipe_phv_out_data_317(mau_3_io_pipe_phv_out_data_317),
    .io_pipe_phv_out_data_318(mau_3_io_pipe_phv_out_data_318),
    .io_pipe_phv_out_data_319(mau_3_io_pipe_phv_out_data_319),
    .io_pipe_phv_out_data_320(mau_3_io_pipe_phv_out_data_320),
    .io_pipe_phv_out_data_321(mau_3_io_pipe_phv_out_data_321),
    .io_pipe_phv_out_data_322(mau_3_io_pipe_phv_out_data_322),
    .io_pipe_phv_out_data_323(mau_3_io_pipe_phv_out_data_323),
    .io_pipe_phv_out_data_324(mau_3_io_pipe_phv_out_data_324),
    .io_pipe_phv_out_data_325(mau_3_io_pipe_phv_out_data_325),
    .io_pipe_phv_out_data_326(mau_3_io_pipe_phv_out_data_326),
    .io_pipe_phv_out_data_327(mau_3_io_pipe_phv_out_data_327),
    .io_pipe_phv_out_data_328(mau_3_io_pipe_phv_out_data_328),
    .io_pipe_phv_out_data_329(mau_3_io_pipe_phv_out_data_329),
    .io_pipe_phv_out_data_330(mau_3_io_pipe_phv_out_data_330),
    .io_pipe_phv_out_data_331(mau_3_io_pipe_phv_out_data_331),
    .io_pipe_phv_out_data_332(mau_3_io_pipe_phv_out_data_332),
    .io_pipe_phv_out_data_333(mau_3_io_pipe_phv_out_data_333),
    .io_pipe_phv_out_data_334(mau_3_io_pipe_phv_out_data_334),
    .io_pipe_phv_out_data_335(mau_3_io_pipe_phv_out_data_335),
    .io_pipe_phv_out_data_336(mau_3_io_pipe_phv_out_data_336),
    .io_pipe_phv_out_data_337(mau_3_io_pipe_phv_out_data_337),
    .io_pipe_phv_out_data_338(mau_3_io_pipe_phv_out_data_338),
    .io_pipe_phv_out_data_339(mau_3_io_pipe_phv_out_data_339),
    .io_pipe_phv_out_data_340(mau_3_io_pipe_phv_out_data_340),
    .io_pipe_phv_out_data_341(mau_3_io_pipe_phv_out_data_341),
    .io_pipe_phv_out_data_342(mau_3_io_pipe_phv_out_data_342),
    .io_pipe_phv_out_data_343(mau_3_io_pipe_phv_out_data_343),
    .io_pipe_phv_out_data_344(mau_3_io_pipe_phv_out_data_344),
    .io_pipe_phv_out_data_345(mau_3_io_pipe_phv_out_data_345),
    .io_pipe_phv_out_data_346(mau_3_io_pipe_phv_out_data_346),
    .io_pipe_phv_out_data_347(mau_3_io_pipe_phv_out_data_347),
    .io_pipe_phv_out_data_348(mau_3_io_pipe_phv_out_data_348),
    .io_pipe_phv_out_data_349(mau_3_io_pipe_phv_out_data_349),
    .io_pipe_phv_out_data_350(mau_3_io_pipe_phv_out_data_350),
    .io_pipe_phv_out_data_351(mau_3_io_pipe_phv_out_data_351),
    .io_pipe_phv_out_data_352(mau_3_io_pipe_phv_out_data_352),
    .io_pipe_phv_out_data_353(mau_3_io_pipe_phv_out_data_353),
    .io_pipe_phv_out_data_354(mau_3_io_pipe_phv_out_data_354),
    .io_pipe_phv_out_data_355(mau_3_io_pipe_phv_out_data_355),
    .io_pipe_phv_out_data_356(mau_3_io_pipe_phv_out_data_356),
    .io_pipe_phv_out_data_357(mau_3_io_pipe_phv_out_data_357),
    .io_pipe_phv_out_data_358(mau_3_io_pipe_phv_out_data_358),
    .io_pipe_phv_out_data_359(mau_3_io_pipe_phv_out_data_359),
    .io_pipe_phv_out_data_360(mau_3_io_pipe_phv_out_data_360),
    .io_pipe_phv_out_data_361(mau_3_io_pipe_phv_out_data_361),
    .io_pipe_phv_out_data_362(mau_3_io_pipe_phv_out_data_362),
    .io_pipe_phv_out_data_363(mau_3_io_pipe_phv_out_data_363),
    .io_pipe_phv_out_data_364(mau_3_io_pipe_phv_out_data_364),
    .io_pipe_phv_out_data_365(mau_3_io_pipe_phv_out_data_365),
    .io_pipe_phv_out_data_366(mau_3_io_pipe_phv_out_data_366),
    .io_pipe_phv_out_data_367(mau_3_io_pipe_phv_out_data_367),
    .io_pipe_phv_out_data_368(mau_3_io_pipe_phv_out_data_368),
    .io_pipe_phv_out_data_369(mau_3_io_pipe_phv_out_data_369),
    .io_pipe_phv_out_data_370(mau_3_io_pipe_phv_out_data_370),
    .io_pipe_phv_out_data_371(mau_3_io_pipe_phv_out_data_371),
    .io_pipe_phv_out_data_372(mau_3_io_pipe_phv_out_data_372),
    .io_pipe_phv_out_data_373(mau_3_io_pipe_phv_out_data_373),
    .io_pipe_phv_out_data_374(mau_3_io_pipe_phv_out_data_374),
    .io_pipe_phv_out_data_375(mau_3_io_pipe_phv_out_data_375),
    .io_pipe_phv_out_data_376(mau_3_io_pipe_phv_out_data_376),
    .io_pipe_phv_out_data_377(mau_3_io_pipe_phv_out_data_377),
    .io_pipe_phv_out_data_378(mau_3_io_pipe_phv_out_data_378),
    .io_pipe_phv_out_data_379(mau_3_io_pipe_phv_out_data_379),
    .io_pipe_phv_out_data_380(mau_3_io_pipe_phv_out_data_380),
    .io_pipe_phv_out_data_381(mau_3_io_pipe_phv_out_data_381),
    .io_pipe_phv_out_data_382(mau_3_io_pipe_phv_out_data_382),
    .io_pipe_phv_out_data_383(mau_3_io_pipe_phv_out_data_383),
    .io_pipe_phv_out_data_384(mau_3_io_pipe_phv_out_data_384),
    .io_pipe_phv_out_data_385(mau_3_io_pipe_phv_out_data_385),
    .io_pipe_phv_out_data_386(mau_3_io_pipe_phv_out_data_386),
    .io_pipe_phv_out_data_387(mau_3_io_pipe_phv_out_data_387),
    .io_pipe_phv_out_data_388(mau_3_io_pipe_phv_out_data_388),
    .io_pipe_phv_out_data_389(mau_3_io_pipe_phv_out_data_389),
    .io_pipe_phv_out_data_390(mau_3_io_pipe_phv_out_data_390),
    .io_pipe_phv_out_data_391(mau_3_io_pipe_phv_out_data_391),
    .io_pipe_phv_out_data_392(mau_3_io_pipe_phv_out_data_392),
    .io_pipe_phv_out_data_393(mau_3_io_pipe_phv_out_data_393),
    .io_pipe_phv_out_data_394(mau_3_io_pipe_phv_out_data_394),
    .io_pipe_phv_out_data_395(mau_3_io_pipe_phv_out_data_395),
    .io_pipe_phv_out_data_396(mau_3_io_pipe_phv_out_data_396),
    .io_pipe_phv_out_data_397(mau_3_io_pipe_phv_out_data_397),
    .io_pipe_phv_out_data_398(mau_3_io_pipe_phv_out_data_398),
    .io_pipe_phv_out_data_399(mau_3_io_pipe_phv_out_data_399),
    .io_pipe_phv_out_data_400(mau_3_io_pipe_phv_out_data_400),
    .io_pipe_phv_out_data_401(mau_3_io_pipe_phv_out_data_401),
    .io_pipe_phv_out_data_402(mau_3_io_pipe_phv_out_data_402),
    .io_pipe_phv_out_data_403(mau_3_io_pipe_phv_out_data_403),
    .io_pipe_phv_out_data_404(mau_3_io_pipe_phv_out_data_404),
    .io_pipe_phv_out_data_405(mau_3_io_pipe_phv_out_data_405),
    .io_pipe_phv_out_data_406(mau_3_io_pipe_phv_out_data_406),
    .io_pipe_phv_out_data_407(mau_3_io_pipe_phv_out_data_407),
    .io_pipe_phv_out_data_408(mau_3_io_pipe_phv_out_data_408),
    .io_pipe_phv_out_data_409(mau_3_io_pipe_phv_out_data_409),
    .io_pipe_phv_out_data_410(mau_3_io_pipe_phv_out_data_410),
    .io_pipe_phv_out_data_411(mau_3_io_pipe_phv_out_data_411),
    .io_pipe_phv_out_data_412(mau_3_io_pipe_phv_out_data_412),
    .io_pipe_phv_out_data_413(mau_3_io_pipe_phv_out_data_413),
    .io_pipe_phv_out_data_414(mau_3_io_pipe_phv_out_data_414),
    .io_pipe_phv_out_data_415(mau_3_io_pipe_phv_out_data_415),
    .io_pipe_phv_out_data_416(mau_3_io_pipe_phv_out_data_416),
    .io_pipe_phv_out_data_417(mau_3_io_pipe_phv_out_data_417),
    .io_pipe_phv_out_data_418(mau_3_io_pipe_phv_out_data_418),
    .io_pipe_phv_out_data_419(mau_3_io_pipe_phv_out_data_419),
    .io_pipe_phv_out_data_420(mau_3_io_pipe_phv_out_data_420),
    .io_pipe_phv_out_data_421(mau_3_io_pipe_phv_out_data_421),
    .io_pipe_phv_out_data_422(mau_3_io_pipe_phv_out_data_422),
    .io_pipe_phv_out_data_423(mau_3_io_pipe_phv_out_data_423),
    .io_pipe_phv_out_data_424(mau_3_io_pipe_phv_out_data_424),
    .io_pipe_phv_out_data_425(mau_3_io_pipe_phv_out_data_425),
    .io_pipe_phv_out_data_426(mau_3_io_pipe_phv_out_data_426),
    .io_pipe_phv_out_data_427(mau_3_io_pipe_phv_out_data_427),
    .io_pipe_phv_out_data_428(mau_3_io_pipe_phv_out_data_428),
    .io_pipe_phv_out_data_429(mau_3_io_pipe_phv_out_data_429),
    .io_pipe_phv_out_data_430(mau_3_io_pipe_phv_out_data_430),
    .io_pipe_phv_out_data_431(mau_3_io_pipe_phv_out_data_431),
    .io_pipe_phv_out_data_432(mau_3_io_pipe_phv_out_data_432),
    .io_pipe_phv_out_data_433(mau_3_io_pipe_phv_out_data_433),
    .io_pipe_phv_out_data_434(mau_3_io_pipe_phv_out_data_434),
    .io_pipe_phv_out_data_435(mau_3_io_pipe_phv_out_data_435),
    .io_pipe_phv_out_data_436(mau_3_io_pipe_phv_out_data_436),
    .io_pipe_phv_out_data_437(mau_3_io_pipe_phv_out_data_437),
    .io_pipe_phv_out_data_438(mau_3_io_pipe_phv_out_data_438),
    .io_pipe_phv_out_data_439(mau_3_io_pipe_phv_out_data_439),
    .io_pipe_phv_out_data_440(mau_3_io_pipe_phv_out_data_440),
    .io_pipe_phv_out_data_441(mau_3_io_pipe_phv_out_data_441),
    .io_pipe_phv_out_data_442(mau_3_io_pipe_phv_out_data_442),
    .io_pipe_phv_out_data_443(mau_3_io_pipe_phv_out_data_443),
    .io_pipe_phv_out_data_444(mau_3_io_pipe_phv_out_data_444),
    .io_pipe_phv_out_data_445(mau_3_io_pipe_phv_out_data_445),
    .io_pipe_phv_out_data_446(mau_3_io_pipe_phv_out_data_446),
    .io_pipe_phv_out_data_447(mau_3_io_pipe_phv_out_data_447),
    .io_pipe_phv_out_data_448(mau_3_io_pipe_phv_out_data_448),
    .io_pipe_phv_out_data_449(mau_3_io_pipe_phv_out_data_449),
    .io_pipe_phv_out_data_450(mau_3_io_pipe_phv_out_data_450),
    .io_pipe_phv_out_data_451(mau_3_io_pipe_phv_out_data_451),
    .io_pipe_phv_out_data_452(mau_3_io_pipe_phv_out_data_452),
    .io_pipe_phv_out_data_453(mau_3_io_pipe_phv_out_data_453),
    .io_pipe_phv_out_data_454(mau_3_io_pipe_phv_out_data_454),
    .io_pipe_phv_out_data_455(mau_3_io_pipe_phv_out_data_455),
    .io_pipe_phv_out_data_456(mau_3_io_pipe_phv_out_data_456),
    .io_pipe_phv_out_data_457(mau_3_io_pipe_phv_out_data_457),
    .io_pipe_phv_out_data_458(mau_3_io_pipe_phv_out_data_458),
    .io_pipe_phv_out_data_459(mau_3_io_pipe_phv_out_data_459),
    .io_pipe_phv_out_data_460(mau_3_io_pipe_phv_out_data_460),
    .io_pipe_phv_out_data_461(mau_3_io_pipe_phv_out_data_461),
    .io_pipe_phv_out_data_462(mau_3_io_pipe_phv_out_data_462),
    .io_pipe_phv_out_data_463(mau_3_io_pipe_phv_out_data_463),
    .io_pipe_phv_out_data_464(mau_3_io_pipe_phv_out_data_464),
    .io_pipe_phv_out_data_465(mau_3_io_pipe_phv_out_data_465),
    .io_pipe_phv_out_data_466(mau_3_io_pipe_phv_out_data_466),
    .io_pipe_phv_out_data_467(mau_3_io_pipe_phv_out_data_467),
    .io_pipe_phv_out_data_468(mau_3_io_pipe_phv_out_data_468),
    .io_pipe_phv_out_data_469(mau_3_io_pipe_phv_out_data_469),
    .io_pipe_phv_out_data_470(mau_3_io_pipe_phv_out_data_470),
    .io_pipe_phv_out_data_471(mau_3_io_pipe_phv_out_data_471),
    .io_pipe_phv_out_data_472(mau_3_io_pipe_phv_out_data_472),
    .io_pipe_phv_out_data_473(mau_3_io_pipe_phv_out_data_473),
    .io_pipe_phv_out_data_474(mau_3_io_pipe_phv_out_data_474),
    .io_pipe_phv_out_data_475(mau_3_io_pipe_phv_out_data_475),
    .io_pipe_phv_out_data_476(mau_3_io_pipe_phv_out_data_476),
    .io_pipe_phv_out_data_477(mau_3_io_pipe_phv_out_data_477),
    .io_pipe_phv_out_data_478(mau_3_io_pipe_phv_out_data_478),
    .io_pipe_phv_out_data_479(mau_3_io_pipe_phv_out_data_479),
    .io_pipe_phv_out_data_480(mau_3_io_pipe_phv_out_data_480),
    .io_pipe_phv_out_data_481(mau_3_io_pipe_phv_out_data_481),
    .io_pipe_phv_out_data_482(mau_3_io_pipe_phv_out_data_482),
    .io_pipe_phv_out_data_483(mau_3_io_pipe_phv_out_data_483),
    .io_pipe_phv_out_data_484(mau_3_io_pipe_phv_out_data_484),
    .io_pipe_phv_out_data_485(mau_3_io_pipe_phv_out_data_485),
    .io_pipe_phv_out_data_486(mau_3_io_pipe_phv_out_data_486),
    .io_pipe_phv_out_data_487(mau_3_io_pipe_phv_out_data_487),
    .io_pipe_phv_out_data_488(mau_3_io_pipe_phv_out_data_488),
    .io_pipe_phv_out_data_489(mau_3_io_pipe_phv_out_data_489),
    .io_pipe_phv_out_data_490(mau_3_io_pipe_phv_out_data_490),
    .io_pipe_phv_out_data_491(mau_3_io_pipe_phv_out_data_491),
    .io_pipe_phv_out_data_492(mau_3_io_pipe_phv_out_data_492),
    .io_pipe_phv_out_data_493(mau_3_io_pipe_phv_out_data_493),
    .io_pipe_phv_out_data_494(mau_3_io_pipe_phv_out_data_494),
    .io_pipe_phv_out_data_495(mau_3_io_pipe_phv_out_data_495),
    .io_pipe_phv_out_data_496(mau_3_io_pipe_phv_out_data_496),
    .io_pipe_phv_out_data_497(mau_3_io_pipe_phv_out_data_497),
    .io_pipe_phv_out_data_498(mau_3_io_pipe_phv_out_data_498),
    .io_pipe_phv_out_data_499(mau_3_io_pipe_phv_out_data_499),
    .io_pipe_phv_out_data_500(mau_3_io_pipe_phv_out_data_500),
    .io_pipe_phv_out_data_501(mau_3_io_pipe_phv_out_data_501),
    .io_pipe_phv_out_data_502(mau_3_io_pipe_phv_out_data_502),
    .io_pipe_phv_out_data_503(mau_3_io_pipe_phv_out_data_503),
    .io_pipe_phv_out_data_504(mau_3_io_pipe_phv_out_data_504),
    .io_pipe_phv_out_data_505(mau_3_io_pipe_phv_out_data_505),
    .io_pipe_phv_out_data_506(mau_3_io_pipe_phv_out_data_506),
    .io_pipe_phv_out_data_507(mau_3_io_pipe_phv_out_data_507),
    .io_pipe_phv_out_data_508(mau_3_io_pipe_phv_out_data_508),
    .io_pipe_phv_out_data_509(mau_3_io_pipe_phv_out_data_509),
    .io_pipe_phv_out_data_510(mau_3_io_pipe_phv_out_data_510),
    .io_pipe_phv_out_data_511(mau_3_io_pipe_phv_out_data_511),
    .io_pipe_phv_out_header_0(mau_3_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(mau_3_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(mau_3_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(mau_3_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(mau_3_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(mau_3_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(mau_3_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(mau_3_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(mau_3_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(mau_3_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(mau_3_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(mau_3_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(mau_3_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(mau_3_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(mau_3_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(mau_3_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(mau_3_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(mau_3_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(mau_3_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(mau_3_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(mau_3_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(mau_3_io_pipe_phv_out_is_valid_processor),
    .io_mod_state_id_mod(mau_3_io_mod_state_id_mod),
    .io_mod_state_id(mau_3_io_mod_state_id),
    .io_mod_sram_w_cs(mau_3_io_mod_sram_w_cs),
    .io_mod_sram_w_en(mau_3_io_mod_sram_w_en),
    .io_mod_sram_w_addr(mau_3_io_mod_sram_w_addr),
    .io_mod_sram_w_data(mau_3_io_mod_sram_w_data)
  );
  ParseModule mau_4 ( // @[parser_pisa.scala 31:25]
    .clock(mau_4_clock),
    .io_pipe_phv_in_data_0(mau_4_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(mau_4_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(mau_4_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(mau_4_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(mau_4_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(mau_4_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(mau_4_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(mau_4_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(mau_4_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(mau_4_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(mau_4_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(mau_4_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(mau_4_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(mau_4_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(mau_4_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(mau_4_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(mau_4_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(mau_4_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(mau_4_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(mau_4_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(mau_4_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(mau_4_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(mau_4_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(mau_4_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(mau_4_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(mau_4_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(mau_4_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(mau_4_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(mau_4_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(mau_4_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(mau_4_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(mau_4_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(mau_4_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(mau_4_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(mau_4_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(mau_4_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(mau_4_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(mau_4_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(mau_4_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(mau_4_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(mau_4_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(mau_4_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(mau_4_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(mau_4_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(mau_4_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(mau_4_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(mau_4_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(mau_4_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(mau_4_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(mau_4_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(mau_4_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(mau_4_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(mau_4_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(mau_4_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(mau_4_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(mau_4_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(mau_4_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(mau_4_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(mau_4_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(mau_4_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(mau_4_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(mau_4_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(mau_4_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(mau_4_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(mau_4_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(mau_4_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(mau_4_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(mau_4_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(mau_4_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(mau_4_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(mau_4_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(mau_4_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(mau_4_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(mau_4_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(mau_4_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(mau_4_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(mau_4_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(mau_4_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(mau_4_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(mau_4_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(mau_4_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(mau_4_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(mau_4_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(mau_4_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(mau_4_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(mau_4_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(mau_4_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(mau_4_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(mau_4_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(mau_4_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(mau_4_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(mau_4_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(mau_4_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(mau_4_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(mau_4_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(mau_4_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(mau_4_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(mau_4_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(mau_4_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(mau_4_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(mau_4_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(mau_4_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(mau_4_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(mau_4_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(mau_4_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(mau_4_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(mau_4_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(mau_4_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(mau_4_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(mau_4_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(mau_4_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(mau_4_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(mau_4_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(mau_4_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(mau_4_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(mau_4_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(mau_4_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(mau_4_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(mau_4_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(mau_4_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(mau_4_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(mau_4_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(mau_4_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(mau_4_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(mau_4_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(mau_4_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(mau_4_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(mau_4_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(mau_4_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(mau_4_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(mau_4_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(mau_4_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(mau_4_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(mau_4_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(mau_4_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(mau_4_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(mau_4_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(mau_4_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(mau_4_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(mau_4_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(mau_4_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(mau_4_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(mau_4_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(mau_4_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(mau_4_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(mau_4_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(mau_4_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(mau_4_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(mau_4_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(mau_4_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(mau_4_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(mau_4_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(mau_4_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(mau_4_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(mau_4_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(mau_4_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(mau_4_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(mau_4_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(mau_4_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(mau_4_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(mau_4_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(mau_4_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(mau_4_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(mau_4_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(mau_4_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(mau_4_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(mau_4_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(mau_4_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(mau_4_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(mau_4_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(mau_4_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(mau_4_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(mau_4_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(mau_4_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(mau_4_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(mau_4_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(mau_4_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(mau_4_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(mau_4_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(mau_4_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(mau_4_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(mau_4_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(mau_4_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(mau_4_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(mau_4_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(mau_4_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(mau_4_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(mau_4_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(mau_4_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(mau_4_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(mau_4_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(mau_4_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(mau_4_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(mau_4_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(mau_4_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(mau_4_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(mau_4_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(mau_4_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(mau_4_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(mau_4_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(mau_4_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(mau_4_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(mau_4_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(mau_4_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(mau_4_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(mau_4_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(mau_4_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(mau_4_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(mau_4_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(mau_4_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(mau_4_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(mau_4_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(mau_4_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(mau_4_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(mau_4_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(mau_4_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(mau_4_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(mau_4_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(mau_4_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(mau_4_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(mau_4_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(mau_4_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(mau_4_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(mau_4_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(mau_4_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(mau_4_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(mau_4_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(mau_4_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(mau_4_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(mau_4_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(mau_4_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(mau_4_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(mau_4_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(mau_4_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(mau_4_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(mau_4_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(mau_4_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(mau_4_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(mau_4_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(mau_4_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(mau_4_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(mau_4_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(mau_4_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(mau_4_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(mau_4_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(mau_4_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(mau_4_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(mau_4_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(mau_4_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(mau_4_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(mau_4_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(mau_4_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(mau_4_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(mau_4_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(mau_4_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(mau_4_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_data_256(mau_4_io_pipe_phv_in_data_256),
    .io_pipe_phv_in_data_257(mau_4_io_pipe_phv_in_data_257),
    .io_pipe_phv_in_data_258(mau_4_io_pipe_phv_in_data_258),
    .io_pipe_phv_in_data_259(mau_4_io_pipe_phv_in_data_259),
    .io_pipe_phv_in_data_260(mau_4_io_pipe_phv_in_data_260),
    .io_pipe_phv_in_data_261(mau_4_io_pipe_phv_in_data_261),
    .io_pipe_phv_in_data_262(mau_4_io_pipe_phv_in_data_262),
    .io_pipe_phv_in_data_263(mau_4_io_pipe_phv_in_data_263),
    .io_pipe_phv_in_data_264(mau_4_io_pipe_phv_in_data_264),
    .io_pipe_phv_in_data_265(mau_4_io_pipe_phv_in_data_265),
    .io_pipe_phv_in_data_266(mau_4_io_pipe_phv_in_data_266),
    .io_pipe_phv_in_data_267(mau_4_io_pipe_phv_in_data_267),
    .io_pipe_phv_in_data_268(mau_4_io_pipe_phv_in_data_268),
    .io_pipe_phv_in_data_269(mau_4_io_pipe_phv_in_data_269),
    .io_pipe_phv_in_data_270(mau_4_io_pipe_phv_in_data_270),
    .io_pipe_phv_in_data_271(mau_4_io_pipe_phv_in_data_271),
    .io_pipe_phv_in_data_272(mau_4_io_pipe_phv_in_data_272),
    .io_pipe_phv_in_data_273(mau_4_io_pipe_phv_in_data_273),
    .io_pipe_phv_in_data_274(mau_4_io_pipe_phv_in_data_274),
    .io_pipe_phv_in_data_275(mau_4_io_pipe_phv_in_data_275),
    .io_pipe_phv_in_data_276(mau_4_io_pipe_phv_in_data_276),
    .io_pipe_phv_in_data_277(mau_4_io_pipe_phv_in_data_277),
    .io_pipe_phv_in_data_278(mau_4_io_pipe_phv_in_data_278),
    .io_pipe_phv_in_data_279(mau_4_io_pipe_phv_in_data_279),
    .io_pipe_phv_in_data_280(mau_4_io_pipe_phv_in_data_280),
    .io_pipe_phv_in_data_281(mau_4_io_pipe_phv_in_data_281),
    .io_pipe_phv_in_data_282(mau_4_io_pipe_phv_in_data_282),
    .io_pipe_phv_in_data_283(mau_4_io_pipe_phv_in_data_283),
    .io_pipe_phv_in_data_284(mau_4_io_pipe_phv_in_data_284),
    .io_pipe_phv_in_data_285(mau_4_io_pipe_phv_in_data_285),
    .io_pipe_phv_in_data_286(mau_4_io_pipe_phv_in_data_286),
    .io_pipe_phv_in_data_287(mau_4_io_pipe_phv_in_data_287),
    .io_pipe_phv_in_data_288(mau_4_io_pipe_phv_in_data_288),
    .io_pipe_phv_in_data_289(mau_4_io_pipe_phv_in_data_289),
    .io_pipe_phv_in_data_290(mau_4_io_pipe_phv_in_data_290),
    .io_pipe_phv_in_data_291(mau_4_io_pipe_phv_in_data_291),
    .io_pipe_phv_in_data_292(mau_4_io_pipe_phv_in_data_292),
    .io_pipe_phv_in_data_293(mau_4_io_pipe_phv_in_data_293),
    .io_pipe_phv_in_data_294(mau_4_io_pipe_phv_in_data_294),
    .io_pipe_phv_in_data_295(mau_4_io_pipe_phv_in_data_295),
    .io_pipe_phv_in_data_296(mau_4_io_pipe_phv_in_data_296),
    .io_pipe_phv_in_data_297(mau_4_io_pipe_phv_in_data_297),
    .io_pipe_phv_in_data_298(mau_4_io_pipe_phv_in_data_298),
    .io_pipe_phv_in_data_299(mau_4_io_pipe_phv_in_data_299),
    .io_pipe_phv_in_data_300(mau_4_io_pipe_phv_in_data_300),
    .io_pipe_phv_in_data_301(mau_4_io_pipe_phv_in_data_301),
    .io_pipe_phv_in_data_302(mau_4_io_pipe_phv_in_data_302),
    .io_pipe_phv_in_data_303(mau_4_io_pipe_phv_in_data_303),
    .io_pipe_phv_in_data_304(mau_4_io_pipe_phv_in_data_304),
    .io_pipe_phv_in_data_305(mau_4_io_pipe_phv_in_data_305),
    .io_pipe_phv_in_data_306(mau_4_io_pipe_phv_in_data_306),
    .io_pipe_phv_in_data_307(mau_4_io_pipe_phv_in_data_307),
    .io_pipe_phv_in_data_308(mau_4_io_pipe_phv_in_data_308),
    .io_pipe_phv_in_data_309(mau_4_io_pipe_phv_in_data_309),
    .io_pipe_phv_in_data_310(mau_4_io_pipe_phv_in_data_310),
    .io_pipe_phv_in_data_311(mau_4_io_pipe_phv_in_data_311),
    .io_pipe_phv_in_data_312(mau_4_io_pipe_phv_in_data_312),
    .io_pipe_phv_in_data_313(mau_4_io_pipe_phv_in_data_313),
    .io_pipe_phv_in_data_314(mau_4_io_pipe_phv_in_data_314),
    .io_pipe_phv_in_data_315(mau_4_io_pipe_phv_in_data_315),
    .io_pipe_phv_in_data_316(mau_4_io_pipe_phv_in_data_316),
    .io_pipe_phv_in_data_317(mau_4_io_pipe_phv_in_data_317),
    .io_pipe_phv_in_data_318(mau_4_io_pipe_phv_in_data_318),
    .io_pipe_phv_in_data_319(mau_4_io_pipe_phv_in_data_319),
    .io_pipe_phv_in_data_320(mau_4_io_pipe_phv_in_data_320),
    .io_pipe_phv_in_data_321(mau_4_io_pipe_phv_in_data_321),
    .io_pipe_phv_in_data_322(mau_4_io_pipe_phv_in_data_322),
    .io_pipe_phv_in_data_323(mau_4_io_pipe_phv_in_data_323),
    .io_pipe_phv_in_data_324(mau_4_io_pipe_phv_in_data_324),
    .io_pipe_phv_in_data_325(mau_4_io_pipe_phv_in_data_325),
    .io_pipe_phv_in_data_326(mau_4_io_pipe_phv_in_data_326),
    .io_pipe_phv_in_data_327(mau_4_io_pipe_phv_in_data_327),
    .io_pipe_phv_in_data_328(mau_4_io_pipe_phv_in_data_328),
    .io_pipe_phv_in_data_329(mau_4_io_pipe_phv_in_data_329),
    .io_pipe_phv_in_data_330(mau_4_io_pipe_phv_in_data_330),
    .io_pipe_phv_in_data_331(mau_4_io_pipe_phv_in_data_331),
    .io_pipe_phv_in_data_332(mau_4_io_pipe_phv_in_data_332),
    .io_pipe_phv_in_data_333(mau_4_io_pipe_phv_in_data_333),
    .io_pipe_phv_in_data_334(mau_4_io_pipe_phv_in_data_334),
    .io_pipe_phv_in_data_335(mau_4_io_pipe_phv_in_data_335),
    .io_pipe_phv_in_data_336(mau_4_io_pipe_phv_in_data_336),
    .io_pipe_phv_in_data_337(mau_4_io_pipe_phv_in_data_337),
    .io_pipe_phv_in_data_338(mau_4_io_pipe_phv_in_data_338),
    .io_pipe_phv_in_data_339(mau_4_io_pipe_phv_in_data_339),
    .io_pipe_phv_in_data_340(mau_4_io_pipe_phv_in_data_340),
    .io_pipe_phv_in_data_341(mau_4_io_pipe_phv_in_data_341),
    .io_pipe_phv_in_data_342(mau_4_io_pipe_phv_in_data_342),
    .io_pipe_phv_in_data_343(mau_4_io_pipe_phv_in_data_343),
    .io_pipe_phv_in_data_344(mau_4_io_pipe_phv_in_data_344),
    .io_pipe_phv_in_data_345(mau_4_io_pipe_phv_in_data_345),
    .io_pipe_phv_in_data_346(mau_4_io_pipe_phv_in_data_346),
    .io_pipe_phv_in_data_347(mau_4_io_pipe_phv_in_data_347),
    .io_pipe_phv_in_data_348(mau_4_io_pipe_phv_in_data_348),
    .io_pipe_phv_in_data_349(mau_4_io_pipe_phv_in_data_349),
    .io_pipe_phv_in_data_350(mau_4_io_pipe_phv_in_data_350),
    .io_pipe_phv_in_data_351(mau_4_io_pipe_phv_in_data_351),
    .io_pipe_phv_in_data_352(mau_4_io_pipe_phv_in_data_352),
    .io_pipe_phv_in_data_353(mau_4_io_pipe_phv_in_data_353),
    .io_pipe_phv_in_data_354(mau_4_io_pipe_phv_in_data_354),
    .io_pipe_phv_in_data_355(mau_4_io_pipe_phv_in_data_355),
    .io_pipe_phv_in_data_356(mau_4_io_pipe_phv_in_data_356),
    .io_pipe_phv_in_data_357(mau_4_io_pipe_phv_in_data_357),
    .io_pipe_phv_in_data_358(mau_4_io_pipe_phv_in_data_358),
    .io_pipe_phv_in_data_359(mau_4_io_pipe_phv_in_data_359),
    .io_pipe_phv_in_data_360(mau_4_io_pipe_phv_in_data_360),
    .io_pipe_phv_in_data_361(mau_4_io_pipe_phv_in_data_361),
    .io_pipe_phv_in_data_362(mau_4_io_pipe_phv_in_data_362),
    .io_pipe_phv_in_data_363(mau_4_io_pipe_phv_in_data_363),
    .io_pipe_phv_in_data_364(mau_4_io_pipe_phv_in_data_364),
    .io_pipe_phv_in_data_365(mau_4_io_pipe_phv_in_data_365),
    .io_pipe_phv_in_data_366(mau_4_io_pipe_phv_in_data_366),
    .io_pipe_phv_in_data_367(mau_4_io_pipe_phv_in_data_367),
    .io_pipe_phv_in_data_368(mau_4_io_pipe_phv_in_data_368),
    .io_pipe_phv_in_data_369(mau_4_io_pipe_phv_in_data_369),
    .io_pipe_phv_in_data_370(mau_4_io_pipe_phv_in_data_370),
    .io_pipe_phv_in_data_371(mau_4_io_pipe_phv_in_data_371),
    .io_pipe_phv_in_data_372(mau_4_io_pipe_phv_in_data_372),
    .io_pipe_phv_in_data_373(mau_4_io_pipe_phv_in_data_373),
    .io_pipe_phv_in_data_374(mau_4_io_pipe_phv_in_data_374),
    .io_pipe_phv_in_data_375(mau_4_io_pipe_phv_in_data_375),
    .io_pipe_phv_in_data_376(mau_4_io_pipe_phv_in_data_376),
    .io_pipe_phv_in_data_377(mau_4_io_pipe_phv_in_data_377),
    .io_pipe_phv_in_data_378(mau_4_io_pipe_phv_in_data_378),
    .io_pipe_phv_in_data_379(mau_4_io_pipe_phv_in_data_379),
    .io_pipe_phv_in_data_380(mau_4_io_pipe_phv_in_data_380),
    .io_pipe_phv_in_data_381(mau_4_io_pipe_phv_in_data_381),
    .io_pipe_phv_in_data_382(mau_4_io_pipe_phv_in_data_382),
    .io_pipe_phv_in_data_383(mau_4_io_pipe_phv_in_data_383),
    .io_pipe_phv_in_data_384(mau_4_io_pipe_phv_in_data_384),
    .io_pipe_phv_in_data_385(mau_4_io_pipe_phv_in_data_385),
    .io_pipe_phv_in_data_386(mau_4_io_pipe_phv_in_data_386),
    .io_pipe_phv_in_data_387(mau_4_io_pipe_phv_in_data_387),
    .io_pipe_phv_in_data_388(mau_4_io_pipe_phv_in_data_388),
    .io_pipe_phv_in_data_389(mau_4_io_pipe_phv_in_data_389),
    .io_pipe_phv_in_data_390(mau_4_io_pipe_phv_in_data_390),
    .io_pipe_phv_in_data_391(mau_4_io_pipe_phv_in_data_391),
    .io_pipe_phv_in_data_392(mau_4_io_pipe_phv_in_data_392),
    .io_pipe_phv_in_data_393(mau_4_io_pipe_phv_in_data_393),
    .io_pipe_phv_in_data_394(mau_4_io_pipe_phv_in_data_394),
    .io_pipe_phv_in_data_395(mau_4_io_pipe_phv_in_data_395),
    .io_pipe_phv_in_data_396(mau_4_io_pipe_phv_in_data_396),
    .io_pipe_phv_in_data_397(mau_4_io_pipe_phv_in_data_397),
    .io_pipe_phv_in_data_398(mau_4_io_pipe_phv_in_data_398),
    .io_pipe_phv_in_data_399(mau_4_io_pipe_phv_in_data_399),
    .io_pipe_phv_in_data_400(mau_4_io_pipe_phv_in_data_400),
    .io_pipe_phv_in_data_401(mau_4_io_pipe_phv_in_data_401),
    .io_pipe_phv_in_data_402(mau_4_io_pipe_phv_in_data_402),
    .io_pipe_phv_in_data_403(mau_4_io_pipe_phv_in_data_403),
    .io_pipe_phv_in_data_404(mau_4_io_pipe_phv_in_data_404),
    .io_pipe_phv_in_data_405(mau_4_io_pipe_phv_in_data_405),
    .io_pipe_phv_in_data_406(mau_4_io_pipe_phv_in_data_406),
    .io_pipe_phv_in_data_407(mau_4_io_pipe_phv_in_data_407),
    .io_pipe_phv_in_data_408(mau_4_io_pipe_phv_in_data_408),
    .io_pipe_phv_in_data_409(mau_4_io_pipe_phv_in_data_409),
    .io_pipe_phv_in_data_410(mau_4_io_pipe_phv_in_data_410),
    .io_pipe_phv_in_data_411(mau_4_io_pipe_phv_in_data_411),
    .io_pipe_phv_in_data_412(mau_4_io_pipe_phv_in_data_412),
    .io_pipe_phv_in_data_413(mau_4_io_pipe_phv_in_data_413),
    .io_pipe_phv_in_data_414(mau_4_io_pipe_phv_in_data_414),
    .io_pipe_phv_in_data_415(mau_4_io_pipe_phv_in_data_415),
    .io_pipe_phv_in_data_416(mau_4_io_pipe_phv_in_data_416),
    .io_pipe_phv_in_data_417(mau_4_io_pipe_phv_in_data_417),
    .io_pipe_phv_in_data_418(mau_4_io_pipe_phv_in_data_418),
    .io_pipe_phv_in_data_419(mau_4_io_pipe_phv_in_data_419),
    .io_pipe_phv_in_data_420(mau_4_io_pipe_phv_in_data_420),
    .io_pipe_phv_in_data_421(mau_4_io_pipe_phv_in_data_421),
    .io_pipe_phv_in_data_422(mau_4_io_pipe_phv_in_data_422),
    .io_pipe_phv_in_data_423(mau_4_io_pipe_phv_in_data_423),
    .io_pipe_phv_in_data_424(mau_4_io_pipe_phv_in_data_424),
    .io_pipe_phv_in_data_425(mau_4_io_pipe_phv_in_data_425),
    .io_pipe_phv_in_data_426(mau_4_io_pipe_phv_in_data_426),
    .io_pipe_phv_in_data_427(mau_4_io_pipe_phv_in_data_427),
    .io_pipe_phv_in_data_428(mau_4_io_pipe_phv_in_data_428),
    .io_pipe_phv_in_data_429(mau_4_io_pipe_phv_in_data_429),
    .io_pipe_phv_in_data_430(mau_4_io_pipe_phv_in_data_430),
    .io_pipe_phv_in_data_431(mau_4_io_pipe_phv_in_data_431),
    .io_pipe_phv_in_data_432(mau_4_io_pipe_phv_in_data_432),
    .io_pipe_phv_in_data_433(mau_4_io_pipe_phv_in_data_433),
    .io_pipe_phv_in_data_434(mau_4_io_pipe_phv_in_data_434),
    .io_pipe_phv_in_data_435(mau_4_io_pipe_phv_in_data_435),
    .io_pipe_phv_in_data_436(mau_4_io_pipe_phv_in_data_436),
    .io_pipe_phv_in_data_437(mau_4_io_pipe_phv_in_data_437),
    .io_pipe_phv_in_data_438(mau_4_io_pipe_phv_in_data_438),
    .io_pipe_phv_in_data_439(mau_4_io_pipe_phv_in_data_439),
    .io_pipe_phv_in_data_440(mau_4_io_pipe_phv_in_data_440),
    .io_pipe_phv_in_data_441(mau_4_io_pipe_phv_in_data_441),
    .io_pipe_phv_in_data_442(mau_4_io_pipe_phv_in_data_442),
    .io_pipe_phv_in_data_443(mau_4_io_pipe_phv_in_data_443),
    .io_pipe_phv_in_data_444(mau_4_io_pipe_phv_in_data_444),
    .io_pipe_phv_in_data_445(mau_4_io_pipe_phv_in_data_445),
    .io_pipe_phv_in_data_446(mau_4_io_pipe_phv_in_data_446),
    .io_pipe_phv_in_data_447(mau_4_io_pipe_phv_in_data_447),
    .io_pipe_phv_in_data_448(mau_4_io_pipe_phv_in_data_448),
    .io_pipe_phv_in_data_449(mau_4_io_pipe_phv_in_data_449),
    .io_pipe_phv_in_data_450(mau_4_io_pipe_phv_in_data_450),
    .io_pipe_phv_in_data_451(mau_4_io_pipe_phv_in_data_451),
    .io_pipe_phv_in_data_452(mau_4_io_pipe_phv_in_data_452),
    .io_pipe_phv_in_data_453(mau_4_io_pipe_phv_in_data_453),
    .io_pipe_phv_in_data_454(mau_4_io_pipe_phv_in_data_454),
    .io_pipe_phv_in_data_455(mau_4_io_pipe_phv_in_data_455),
    .io_pipe_phv_in_data_456(mau_4_io_pipe_phv_in_data_456),
    .io_pipe_phv_in_data_457(mau_4_io_pipe_phv_in_data_457),
    .io_pipe_phv_in_data_458(mau_4_io_pipe_phv_in_data_458),
    .io_pipe_phv_in_data_459(mau_4_io_pipe_phv_in_data_459),
    .io_pipe_phv_in_data_460(mau_4_io_pipe_phv_in_data_460),
    .io_pipe_phv_in_data_461(mau_4_io_pipe_phv_in_data_461),
    .io_pipe_phv_in_data_462(mau_4_io_pipe_phv_in_data_462),
    .io_pipe_phv_in_data_463(mau_4_io_pipe_phv_in_data_463),
    .io_pipe_phv_in_data_464(mau_4_io_pipe_phv_in_data_464),
    .io_pipe_phv_in_data_465(mau_4_io_pipe_phv_in_data_465),
    .io_pipe_phv_in_data_466(mau_4_io_pipe_phv_in_data_466),
    .io_pipe_phv_in_data_467(mau_4_io_pipe_phv_in_data_467),
    .io_pipe_phv_in_data_468(mau_4_io_pipe_phv_in_data_468),
    .io_pipe_phv_in_data_469(mau_4_io_pipe_phv_in_data_469),
    .io_pipe_phv_in_data_470(mau_4_io_pipe_phv_in_data_470),
    .io_pipe_phv_in_data_471(mau_4_io_pipe_phv_in_data_471),
    .io_pipe_phv_in_data_472(mau_4_io_pipe_phv_in_data_472),
    .io_pipe_phv_in_data_473(mau_4_io_pipe_phv_in_data_473),
    .io_pipe_phv_in_data_474(mau_4_io_pipe_phv_in_data_474),
    .io_pipe_phv_in_data_475(mau_4_io_pipe_phv_in_data_475),
    .io_pipe_phv_in_data_476(mau_4_io_pipe_phv_in_data_476),
    .io_pipe_phv_in_data_477(mau_4_io_pipe_phv_in_data_477),
    .io_pipe_phv_in_data_478(mau_4_io_pipe_phv_in_data_478),
    .io_pipe_phv_in_data_479(mau_4_io_pipe_phv_in_data_479),
    .io_pipe_phv_in_data_480(mau_4_io_pipe_phv_in_data_480),
    .io_pipe_phv_in_data_481(mau_4_io_pipe_phv_in_data_481),
    .io_pipe_phv_in_data_482(mau_4_io_pipe_phv_in_data_482),
    .io_pipe_phv_in_data_483(mau_4_io_pipe_phv_in_data_483),
    .io_pipe_phv_in_data_484(mau_4_io_pipe_phv_in_data_484),
    .io_pipe_phv_in_data_485(mau_4_io_pipe_phv_in_data_485),
    .io_pipe_phv_in_data_486(mau_4_io_pipe_phv_in_data_486),
    .io_pipe_phv_in_data_487(mau_4_io_pipe_phv_in_data_487),
    .io_pipe_phv_in_data_488(mau_4_io_pipe_phv_in_data_488),
    .io_pipe_phv_in_data_489(mau_4_io_pipe_phv_in_data_489),
    .io_pipe_phv_in_data_490(mau_4_io_pipe_phv_in_data_490),
    .io_pipe_phv_in_data_491(mau_4_io_pipe_phv_in_data_491),
    .io_pipe_phv_in_data_492(mau_4_io_pipe_phv_in_data_492),
    .io_pipe_phv_in_data_493(mau_4_io_pipe_phv_in_data_493),
    .io_pipe_phv_in_data_494(mau_4_io_pipe_phv_in_data_494),
    .io_pipe_phv_in_data_495(mau_4_io_pipe_phv_in_data_495),
    .io_pipe_phv_in_data_496(mau_4_io_pipe_phv_in_data_496),
    .io_pipe_phv_in_data_497(mau_4_io_pipe_phv_in_data_497),
    .io_pipe_phv_in_data_498(mau_4_io_pipe_phv_in_data_498),
    .io_pipe_phv_in_data_499(mau_4_io_pipe_phv_in_data_499),
    .io_pipe_phv_in_data_500(mau_4_io_pipe_phv_in_data_500),
    .io_pipe_phv_in_data_501(mau_4_io_pipe_phv_in_data_501),
    .io_pipe_phv_in_data_502(mau_4_io_pipe_phv_in_data_502),
    .io_pipe_phv_in_data_503(mau_4_io_pipe_phv_in_data_503),
    .io_pipe_phv_in_data_504(mau_4_io_pipe_phv_in_data_504),
    .io_pipe_phv_in_data_505(mau_4_io_pipe_phv_in_data_505),
    .io_pipe_phv_in_data_506(mau_4_io_pipe_phv_in_data_506),
    .io_pipe_phv_in_data_507(mau_4_io_pipe_phv_in_data_507),
    .io_pipe_phv_in_data_508(mau_4_io_pipe_phv_in_data_508),
    .io_pipe_phv_in_data_509(mau_4_io_pipe_phv_in_data_509),
    .io_pipe_phv_in_data_510(mau_4_io_pipe_phv_in_data_510),
    .io_pipe_phv_in_data_511(mau_4_io_pipe_phv_in_data_511),
    .io_pipe_phv_in_header_0(mau_4_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(mau_4_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(mau_4_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(mau_4_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(mau_4_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(mau_4_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(mau_4_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(mau_4_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(mau_4_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(mau_4_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(mau_4_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(mau_4_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(mau_4_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(mau_4_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(mau_4_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(mau_4_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(mau_4_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(mau_4_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(mau_4_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(mau_4_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(mau_4_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(mau_4_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(mau_4_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(mau_4_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(mau_4_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(mau_4_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(mau_4_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(mau_4_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(mau_4_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(mau_4_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(mau_4_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(mau_4_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(mau_4_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(mau_4_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(mau_4_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(mau_4_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(mau_4_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(mau_4_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(mau_4_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(mau_4_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(mau_4_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(mau_4_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(mau_4_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(mau_4_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(mau_4_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(mau_4_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(mau_4_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(mau_4_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(mau_4_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(mau_4_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(mau_4_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(mau_4_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(mau_4_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(mau_4_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(mau_4_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(mau_4_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(mau_4_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(mau_4_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(mau_4_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(mau_4_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(mau_4_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(mau_4_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(mau_4_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(mau_4_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(mau_4_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(mau_4_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(mau_4_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(mau_4_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(mau_4_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(mau_4_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(mau_4_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(mau_4_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(mau_4_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(mau_4_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(mau_4_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(mau_4_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(mau_4_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(mau_4_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(mau_4_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(mau_4_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(mau_4_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(mau_4_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(mau_4_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(mau_4_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(mau_4_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(mau_4_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(mau_4_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(mau_4_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(mau_4_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(mau_4_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(mau_4_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(mau_4_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(mau_4_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(mau_4_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(mau_4_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(mau_4_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(mau_4_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(mau_4_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(mau_4_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(mau_4_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(mau_4_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(mau_4_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(mau_4_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(mau_4_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(mau_4_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(mau_4_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(mau_4_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(mau_4_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(mau_4_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(mau_4_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(mau_4_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(mau_4_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(mau_4_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(mau_4_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(mau_4_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(mau_4_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(mau_4_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(mau_4_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(mau_4_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(mau_4_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(mau_4_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(mau_4_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(mau_4_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(mau_4_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(mau_4_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(mau_4_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(mau_4_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(mau_4_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(mau_4_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(mau_4_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(mau_4_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(mau_4_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(mau_4_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(mau_4_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(mau_4_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(mau_4_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(mau_4_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(mau_4_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(mau_4_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(mau_4_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(mau_4_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(mau_4_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(mau_4_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(mau_4_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(mau_4_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(mau_4_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(mau_4_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(mau_4_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(mau_4_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(mau_4_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(mau_4_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(mau_4_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(mau_4_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(mau_4_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(mau_4_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(mau_4_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(mau_4_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(mau_4_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(mau_4_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(mau_4_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(mau_4_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(mau_4_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(mau_4_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(mau_4_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(mau_4_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(mau_4_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(mau_4_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(mau_4_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(mau_4_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(mau_4_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(mau_4_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(mau_4_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(mau_4_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(mau_4_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(mau_4_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(mau_4_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(mau_4_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(mau_4_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(mau_4_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(mau_4_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(mau_4_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(mau_4_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(mau_4_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(mau_4_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(mau_4_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(mau_4_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(mau_4_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(mau_4_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(mau_4_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(mau_4_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(mau_4_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(mau_4_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(mau_4_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(mau_4_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(mau_4_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(mau_4_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(mau_4_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(mau_4_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(mau_4_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(mau_4_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(mau_4_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(mau_4_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(mau_4_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(mau_4_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(mau_4_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(mau_4_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(mau_4_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(mau_4_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(mau_4_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(mau_4_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(mau_4_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(mau_4_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(mau_4_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(mau_4_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(mau_4_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(mau_4_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(mau_4_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(mau_4_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(mau_4_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(mau_4_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(mau_4_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(mau_4_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(mau_4_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(mau_4_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(mau_4_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(mau_4_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(mau_4_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(mau_4_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(mau_4_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(mau_4_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(mau_4_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(mau_4_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(mau_4_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(mau_4_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(mau_4_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(mau_4_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(mau_4_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(mau_4_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(mau_4_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(mau_4_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(mau_4_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(mau_4_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(mau_4_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(mau_4_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(mau_4_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(mau_4_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(mau_4_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(mau_4_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(mau_4_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(mau_4_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(mau_4_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(mau_4_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(mau_4_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(mau_4_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(mau_4_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(mau_4_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(mau_4_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(mau_4_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(mau_4_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(mau_4_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(mau_4_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(mau_4_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(mau_4_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(mau_4_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(mau_4_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(mau_4_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(mau_4_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(mau_4_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(mau_4_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(mau_4_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(mau_4_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(mau_4_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(mau_4_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(mau_4_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(mau_4_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(mau_4_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(mau_4_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(mau_4_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_data_256(mau_4_io_pipe_phv_out_data_256),
    .io_pipe_phv_out_data_257(mau_4_io_pipe_phv_out_data_257),
    .io_pipe_phv_out_data_258(mau_4_io_pipe_phv_out_data_258),
    .io_pipe_phv_out_data_259(mau_4_io_pipe_phv_out_data_259),
    .io_pipe_phv_out_data_260(mau_4_io_pipe_phv_out_data_260),
    .io_pipe_phv_out_data_261(mau_4_io_pipe_phv_out_data_261),
    .io_pipe_phv_out_data_262(mau_4_io_pipe_phv_out_data_262),
    .io_pipe_phv_out_data_263(mau_4_io_pipe_phv_out_data_263),
    .io_pipe_phv_out_data_264(mau_4_io_pipe_phv_out_data_264),
    .io_pipe_phv_out_data_265(mau_4_io_pipe_phv_out_data_265),
    .io_pipe_phv_out_data_266(mau_4_io_pipe_phv_out_data_266),
    .io_pipe_phv_out_data_267(mau_4_io_pipe_phv_out_data_267),
    .io_pipe_phv_out_data_268(mau_4_io_pipe_phv_out_data_268),
    .io_pipe_phv_out_data_269(mau_4_io_pipe_phv_out_data_269),
    .io_pipe_phv_out_data_270(mau_4_io_pipe_phv_out_data_270),
    .io_pipe_phv_out_data_271(mau_4_io_pipe_phv_out_data_271),
    .io_pipe_phv_out_data_272(mau_4_io_pipe_phv_out_data_272),
    .io_pipe_phv_out_data_273(mau_4_io_pipe_phv_out_data_273),
    .io_pipe_phv_out_data_274(mau_4_io_pipe_phv_out_data_274),
    .io_pipe_phv_out_data_275(mau_4_io_pipe_phv_out_data_275),
    .io_pipe_phv_out_data_276(mau_4_io_pipe_phv_out_data_276),
    .io_pipe_phv_out_data_277(mau_4_io_pipe_phv_out_data_277),
    .io_pipe_phv_out_data_278(mau_4_io_pipe_phv_out_data_278),
    .io_pipe_phv_out_data_279(mau_4_io_pipe_phv_out_data_279),
    .io_pipe_phv_out_data_280(mau_4_io_pipe_phv_out_data_280),
    .io_pipe_phv_out_data_281(mau_4_io_pipe_phv_out_data_281),
    .io_pipe_phv_out_data_282(mau_4_io_pipe_phv_out_data_282),
    .io_pipe_phv_out_data_283(mau_4_io_pipe_phv_out_data_283),
    .io_pipe_phv_out_data_284(mau_4_io_pipe_phv_out_data_284),
    .io_pipe_phv_out_data_285(mau_4_io_pipe_phv_out_data_285),
    .io_pipe_phv_out_data_286(mau_4_io_pipe_phv_out_data_286),
    .io_pipe_phv_out_data_287(mau_4_io_pipe_phv_out_data_287),
    .io_pipe_phv_out_data_288(mau_4_io_pipe_phv_out_data_288),
    .io_pipe_phv_out_data_289(mau_4_io_pipe_phv_out_data_289),
    .io_pipe_phv_out_data_290(mau_4_io_pipe_phv_out_data_290),
    .io_pipe_phv_out_data_291(mau_4_io_pipe_phv_out_data_291),
    .io_pipe_phv_out_data_292(mau_4_io_pipe_phv_out_data_292),
    .io_pipe_phv_out_data_293(mau_4_io_pipe_phv_out_data_293),
    .io_pipe_phv_out_data_294(mau_4_io_pipe_phv_out_data_294),
    .io_pipe_phv_out_data_295(mau_4_io_pipe_phv_out_data_295),
    .io_pipe_phv_out_data_296(mau_4_io_pipe_phv_out_data_296),
    .io_pipe_phv_out_data_297(mau_4_io_pipe_phv_out_data_297),
    .io_pipe_phv_out_data_298(mau_4_io_pipe_phv_out_data_298),
    .io_pipe_phv_out_data_299(mau_4_io_pipe_phv_out_data_299),
    .io_pipe_phv_out_data_300(mau_4_io_pipe_phv_out_data_300),
    .io_pipe_phv_out_data_301(mau_4_io_pipe_phv_out_data_301),
    .io_pipe_phv_out_data_302(mau_4_io_pipe_phv_out_data_302),
    .io_pipe_phv_out_data_303(mau_4_io_pipe_phv_out_data_303),
    .io_pipe_phv_out_data_304(mau_4_io_pipe_phv_out_data_304),
    .io_pipe_phv_out_data_305(mau_4_io_pipe_phv_out_data_305),
    .io_pipe_phv_out_data_306(mau_4_io_pipe_phv_out_data_306),
    .io_pipe_phv_out_data_307(mau_4_io_pipe_phv_out_data_307),
    .io_pipe_phv_out_data_308(mau_4_io_pipe_phv_out_data_308),
    .io_pipe_phv_out_data_309(mau_4_io_pipe_phv_out_data_309),
    .io_pipe_phv_out_data_310(mau_4_io_pipe_phv_out_data_310),
    .io_pipe_phv_out_data_311(mau_4_io_pipe_phv_out_data_311),
    .io_pipe_phv_out_data_312(mau_4_io_pipe_phv_out_data_312),
    .io_pipe_phv_out_data_313(mau_4_io_pipe_phv_out_data_313),
    .io_pipe_phv_out_data_314(mau_4_io_pipe_phv_out_data_314),
    .io_pipe_phv_out_data_315(mau_4_io_pipe_phv_out_data_315),
    .io_pipe_phv_out_data_316(mau_4_io_pipe_phv_out_data_316),
    .io_pipe_phv_out_data_317(mau_4_io_pipe_phv_out_data_317),
    .io_pipe_phv_out_data_318(mau_4_io_pipe_phv_out_data_318),
    .io_pipe_phv_out_data_319(mau_4_io_pipe_phv_out_data_319),
    .io_pipe_phv_out_data_320(mau_4_io_pipe_phv_out_data_320),
    .io_pipe_phv_out_data_321(mau_4_io_pipe_phv_out_data_321),
    .io_pipe_phv_out_data_322(mau_4_io_pipe_phv_out_data_322),
    .io_pipe_phv_out_data_323(mau_4_io_pipe_phv_out_data_323),
    .io_pipe_phv_out_data_324(mau_4_io_pipe_phv_out_data_324),
    .io_pipe_phv_out_data_325(mau_4_io_pipe_phv_out_data_325),
    .io_pipe_phv_out_data_326(mau_4_io_pipe_phv_out_data_326),
    .io_pipe_phv_out_data_327(mau_4_io_pipe_phv_out_data_327),
    .io_pipe_phv_out_data_328(mau_4_io_pipe_phv_out_data_328),
    .io_pipe_phv_out_data_329(mau_4_io_pipe_phv_out_data_329),
    .io_pipe_phv_out_data_330(mau_4_io_pipe_phv_out_data_330),
    .io_pipe_phv_out_data_331(mau_4_io_pipe_phv_out_data_331),
    .io_pipe_phv_out_data_332(mau_4_io_pipe_phv_out_data_332),
    .io_pipe_phv_out_data_333(mau_4_io_pipe_phv_out_data_333),
    .io_pipe_phv_out_data_334(mau_4_io_pipe_phv_out_data_334),
    .io_pipe_phv_out_data_335(mau_4_io_pipe_phv_out_data_335),
    .io_pipe_phv_out_data_336(mau_4_io_pipe_phv_out_data_336),
    .io_pipe_phv_out_data_337(mau_4_io_pipe_phv_out_data_337),
    .io_pipe_phv_out_data_338(mau_4_io_pipe_phv_out_data_338),
    .io_pipe_phv_out_data_339(mau_4_io_pipe_phv_out_data_339),
    .io_pipe_phv_out_data_340(mau_4_io_pipe_phv_out_data_340),
    .io_pipe_phv_out_data_341(mau_4_io_pipe_phv_out_data_341),
    .io_pipe_phv_out_data_342(mau_4_io_pipe_phv_out_data_342),
    .io_pipe_phv_out_data_343(mau_4_io_pipe_phv_out_data_343),
    .io_pipe_phv_out_data_344(mau_4_io_pipe_phv_out_data_344),
    .io_pipe_phv_out_data_345(mau_4_io_pipe_phv_out_data_345),
    .io_pipe_phv_out_data_346(mau_4_io_pipe_phv_out_data_346),
    .io_pipe_phv_out_data_347(mau_4_io_pipe_phv_out_data_347),
    .io_pipe_phv_out_data_348(mau_4_io_pipe_phv_out_data_348),
    .io_pipe_phv_out_data_349(mau_4_io_pipe_phv_out_data_349),
    .io_pipe_phv_out_data_350(mau_4_io_pipe_phv_out_data_350),
    .io_pipe_phv_out_data_351(mau_4_io_pipe_phv_out_data_351),
    .io_pipe_phv_out_data_352(mau_4_io_pipe_phv_out_data_352),
    .io_pipe_phv_out_data_353(mau_4_io_pipe_phv_out_data_353),
    .io_pipe_phv_out_data_354(mau_4_io_pipe_phv_out_data_354),
    .io_pipe_phv_out_data_355(mau_4_io_pipe_phv_out_data_355),
    .io_pipe_phv_out_data_356(mau_4_io_pipe_phv_out_data_356),
    .io_pipe_phv_out_data_357(mau_4_io_pipe_phv_out_data_357),
    .io_pipe_phv_out_data_358(mau_4_io_pipe_phv_out_data_358),
    .io_pipe_phv_out_data_359(mau_4_io_pipe_phv_out_data_359),
    .io_pipe_phv_out_data_360(mau_4_io_pipe_phv_out_data_360),
    .io_pipe_phv_out_data_361(mau_4_io_pipe_phv_out_data_361),
    .io_pipe_phv_out_data_362(mau_4_io_pipe_phv_out_data_362),
    .io_pipe_phv_out_data_363(mau_4_io_pipe_phv_out_data_363),
    .io_pipe_phv_out_data_364(mau_4_io_pipe_phv_out_data_364),
    .io_pipe_phv_out_data_365(mau_4_io_pipe_phv_out_data_365),
    .io_pipe_phv_out_data_366(mau_4_io_pipe_phv_out_data_366),
    .io_pipe_phv_out_data_367(mau_4_io_pipe_phv_out_data_367),
    .io_pipe_phv_out_data_368(mau_4_io_pipe_phv_out_data_368),
    .io_pipe_phv_out_data_369(mau_4_io_pipe_phv_out_data_369),
    .io_pipe_phv_out_data_370(mau_4_io_pipe_phv_out_data_370),
    .io_pipe_phv_out_data_371(mau_4_io_pipe_phv_out_data_371),
    .io_pipe_phv_out_data_372(mau_4_io_pipe_phv_out_data_372),
    .io_pipe_phv_out_data_373(mau_4_io_pipe_phv_out_data_373),
    .io_pipe_phv_out_data_374(mau_4_io_pipe_phv_out_data_374),
    .io_pipe_phv_out_data_375(mau_4_io_pipe_phv_out_data_375),
    .io_pipe_phv_out_data_376(mau_4_io_pipe_phv_out_data_376),
    .io_pipe_phv_out_data_377(mau_4_io_pipe_phv_out_data_377),
    .io_pipe_phv_out_data_378(mau_4_io_pipe_phv_out_data_378),
    .io_pipe_phv_out_data_379(mau_4_io_pipe_phv_out_data_379),
    .io_pipe_phv_out_data_380(mau_4_io_pipe_phv_out_data_380),
    .io_pipe_phv_out_data_381(mau_4_io_pipe_phv_out_data_381),
    .io_pipe_phv_out_data_382(mau_4_io_pipe_phv_out_data_382),
    .io_pipe_phv_out_data_383(mau_4_io_pipe_phv_out_data_383),
    .io_pipe_phv_out_data_384(mau_4_io_pipe_phv_out_data_384),
    .io_pipe_phv_out_data_385(mau_4_io_pipe_phv_out_data_385),
    .io_pipe_phv_out_data_386(mau_4_io_pipe_phv_out_data_386),
    .io_pipe_phv_out_data_387(mau_4_io_pipe_phv_out_data_387),
    .io_pipe_phv_out_data_388(mau_4_io_pipe_phv_out_data_388),
    .io_pipe_phv_out_data_389(mau_4_io_pipe_phv_out_data_389),
    .io_pipe_phv_out_data_390(mau_4_io_pipe_phv_out_data_390),
    .io_pipe_phv_out_data_391(mau_4_io_pipe_phv_out_data_391),
    .io_pipe_phv_out_data_392(mau_4_io_pipe_phv_out_data_392),
    .io_pipe_phv_out_data_393(mau_4_io_pipe_phv_out_data_393),
    .io_pipe_phv_out_data_394(mau_4_io_pipe_phv_out_data_394),
    .io_pipe_phv_out_data_395(mau_4_io_pipe_phv_out_data_395),
    .io_pipe_phv_out_data_396(mau_4_io_pipe_phv_out_data_396),
    .io_pipe_phv_out_data_397(mau_4_io_pipe_phv_out_data_397),
    .io_pipe_phv_out_data_398(mau_4_io_pipe_phv_out_data_398),
    .io_pipe_phv_out_data_399(mau_4_io_pipe_phv_out_data_399),
    .io_pipe_phv_out_data_400(mau_4_io_pipe_phv_out_data_400),
    .io_pipe_phv_out_data_401(mau_4_io_pipe_phv_out_data_401),
    .io_pipe_phv_out_data_402(mau_4_io_pipe_phv_out_data_402),
    .io_pipe_phv_out_data_403(mau_4_io_pipe_phv_out_data_403),
    .io_pipe_phv_out_data_404(mau_4_io_pipe_phv_out_data_404),
    .io_pipe_phv_out_data_405(mau_4_io_pipe_phv_out_data_405),
    .io_pipe_phv_out_data_406(mau_4_io_pipe_phv_out_data_406),
    .io_pipe_phv_out_data_407(mau_4_io_pipe_phv_out_data_407),
    .io_pipe_phv_out_data_408(mau_4_io_pipe_phv_out_data_408),
    .io_pipe_phv_out_data_409(mau_4_io_pipe_phv_out_data_409),
    .io_pipe_phv_out_data_410(mau_4_io_pipe_phv_out_data_410),
    .io_pipe_phv_out_data_411(mau_4_io_pipe_phv_out_data_411),
    .io_pipe_phv_out_data_412(mau_4_io_pipe_phv_out_data_412),
    .io_pipe_phv_out_data_413(mau_4_io_pipe_phv_out_data_413),
    .io_pipe_phv_out_data_414(mau_4_io_pipe_phv_out_data_414),
    .io_pipe_phv_out_data_415(mau_4_io_pipe_phv_out_data_415),
    .io_pipe_phv_out_data_416(mau_4_io_pipe_phv_out_data_416),
    .io_pipe_phv_out_data_417(mau_4_io_pipe_phv_out_data_417),
    .io_pipe_phv_out_data_418(mau_4_io_pipe_phv_out_data_418),
    .io_pipe_phv_out_data_419(mau_4_io_pipe_phv_out_data_419),
    .io_pipe_phv_out_data_420(mau_4_io_pipe_phv_out_data_420),
    .io_pipe_phv_out_data_421(mau_4_io_pipe_phv_out_data_421),
    .io_pipe_phv_out_data_422(mau_4_io_pipe_phv_out_data_422),
    .io_pipe_phv_out_data_423(mau_4_io_pipe_phv_out_data_423),
    .io_pipe_phv_out_data_424(mau_4_io_pipe_phv_out_data_424),
    .io_pipe_phv_out_data_425(mau_4_io_pipe_phv_out_data_425),
    .io_pipe_phv_out_data_426(mau_4_io_pipe_phv_out_data_426),
    .io_pipe_phv_out_data_427(mau_4_io_pipe_phv_out_data_427),
    .io_pipe_phv_out_data_428(mau_4_io_pipe_phv_out_data_428),
    .io_pipe_phv_out_data_429(mau_4_io_pipe_phv_out_data_429),
    .io_pipe_phv_out_data_430(mau_4_io_pipe_phv_out_data_430),
    .io_pipe_phv_out_data_431(mau_4_io_pipe_phv_out_data_431),
    .io_pipe_phv_out_data_432(mau_4_io_pipe_phv_out_data_432),
    .io_pipe_phv_out_data_433(mau_4_io_pipe_phv_out_data_433),
    .io_pipe_phv_out_data_434(mau_4_io_pipe_phv_out_data_434),
    .io_pipe_phv_out_data_435(mau_4_io_pipe_phv_out_data_435),
    .io_pipe_phv_out_data_436(mau_4_io_pipe_phv_out_data_436),
    .io_pipe_phv_out_data_437(mau_4_io_pipe_phv_out_data_437),
    .io_pipe_phv_out_data_438(mau_4_io_pipe_phv_out_data_438),
    .io_pipe_phv_out_data_439(mau_4_io_pipe_phv_out_data_439),
    .io_pipe_phv_out_data_440(mau_4_io_pipe_phv_out_data_440),
    .io_pipe_phv_out_data_441(mau_4_io_pipe_phv_out_data_441),
    .io_pipe_phv_out_data_442(mau_4_io_pipe_phv_out_data_442),
    .io_pipe_phv_out_data_443(mau_4_io_pipe_phv_out_data_443),
    .io_pipe_phv_out_data_444(mau_4_io_pipe_phv_out_data_444),
    .io_pipe_phv_out_data_445(mau_4_io_pipe_phv_out_data_445),
    .io_pipe_phv_out_data_446(mau_4_io_pipe_phv_out_data_446),
    .io_pipe_phv_out_data_447(mau_4_io_pipe_phv_out_data_447),
    .io_pipe_phv_out_data_448(mau_4_io_pipe_phv_out_data_448),
    .io_pipe_phv_out_data_449(mau_4_io_pipe_phv_out_data_449),
    .io_pipe_phv_out_data_450(mau_4_io_pipe_phv_out_data_450),
    .io_pipe_phv_out_data_451(mau_4_io_pipe_phv_out_data_451),
    .io_pipe_phv_out_data_452(mau_4_io_pipe_phv_out_data_452),
    .io_pipe_phv_out_data_453(mau_4_io_pipe_phv_out_data_453),
    .io_pipe_phv_out_data_454(mau_4_io_pipe_phv_out_data_454),
    .io_pipe_phv_out_data_455(mau_4_io_pipe_phv_out_data_455),
    .io_pipe_phv_out_data_456(mau_4_io_pipe_phv_out_data_456),
    .io_pipe_phv_out_data_457(mau_4_io_pipe_phv_out_data_457),
    .io_pipe_phv_out_data_458(mau_4_io_pipe_phv_out_data_458),
    .io_pipe_phv_out_data_459(mau_4_io_pipe_phv_out_data_459),
    .io_pipe_phv_out_data_460(mau_4_io_pipe_phv_out_data_460),
    .io_pipe_phv_out_data_461(mau_4_io_pipe_phv_out_data_461),
    .io_pipe_phv_out_data_462(mau_4_io_pipe_phv_out_data_462),
    .io_pipe_phv_out_data_463(mau_4_io_pipe_phv_out_data_463),
    .io_pipe_phv_out_data_464(mau_4_io_pipe_phv_out_data_464),
    .io_pipe_phv_out_data_465(mau_4_io_pipe_phv_out_data_465),
    .io_pipe_phv_out_data_466(mau_4_io_pipe_phv_out_data_466),
    .io_pipe_phv_out_data_467(mau_4_io_pipe_phv_out_data_467),
    .io_pipe_phv_out_data_468(mau_4_io_pipe_phv_out_data_468),
    .io_pipe_phv_out_data_469(mau_4_io_pipe_phv_out_data_469),
    .io_pipe_phv_out_data_470(mau_4_io_pipe_phv_out_data_470),
    .io_pipe_phv_out_data_471(mau_4_io_pipe_phv_out_data_471),
    .io_pipe_phv_out_data_472(mau_4_io_pipe_phv_out_data_472),
    .io_pipe_phv_out_data_473(mau_4_io_pipe_phv_out_data_473),
    .io_pipe_phv_out_data_474(mau_4_io_pipe_phv_out_data_474),
    .io_pipe_phv_out_data_475(mau_4_io_pipe_phv_out_data_475),
    .io_pipe_phv_out_data_476(mau_4_io_pipe_phv_out_data_476),
    .io_pipe_phv_out_data_477(mau_4_io_pipe_phv_out_data_477),
    .io_pipe_phv_out_data_478(mau_4_io_pipe_phv_out_data_478),
    .io_pipe_phv_out_data_479(mau_4_io_pipe_phv_out_data_479),
    .io_pipe_phv_out_data_480(mau_4_io_pipe_phv_out_data_480),
    .io_pipe_phv_out_data_481(mau_4_io_pipe_phv_out_data_481),
    .io_pipe_phv_out_data_482(mau_4_io_pipe_phv_out_data_482),
    .io_pipe_phv_out_data_483(mau_4_io_pipe_phv_out_data_483),
    .io_pipe_phv_out_data_484(mau_4_io_pipe_phv_out_data_484),
    .io_pipe_phv_out_data_485(mau_4_io_pipe_phv_out_data_485),
    .io_pipe_phv_out_data_486(mau_4_io_pipe_phv_out_data_486),
    .io_pipe_phv_out_data_487(mau_4_io_pipe_phv_out_data_487),
    .io_pipe_phv_out_data_488(mau_4_io_pipe_phv_out_data_488),
    .io_pipe_phv_out_data_489(mau_4_io_pipe_phv_out_data_489),
    .io_pipe_phv_out_data_490(mau_4_io_pipe_phv_out_data_490),
    .io_pipe_phv_out_data_491(mau_4_io_pipe_phv_out_data_491),
    .io_pipe_phv_out_data_492(mau_4_io_pipe_phv_out_data_492),
    .io_pipe_phv_out_data_493(mau_4_io_pipe_phv_out_data_493),
    .io_pipe_phv_out_data_494(mau_4_io_pipe_phv_out_data_494),
    .io_pipe_phv_out_data_495(mau_4_io_pipe_phv_out_data_495),
    .io_pipe_phv_out_data_496(mau_4_io_pipe_phv_out_data_496),
    .io_pipe_phv_out_data_497(mau_4_io_pipe_phv_out_data_497),
    .io_pipe_phv_out_data_498(mau_4_io_pipe_phv_out_data_498),
    .io_pipe_phv_out_data_499(mau_4_io_pipe_phv_out_data_499),
    .io_pipe_phv_out_data_500(mau_4_io_pipe_phv_out_data_500),
    .io_pipe_phv_out_data_501(mau_4_io_pipe_phv_out_data_501),
    .io_pipe_phv_out_data_502(mau_4_io_pipe_phv_out_data_502),
    .io_pipe_phv_out_data_503(mau_4_io_pipe_phv_out_data_503),
    .io_pipe_phv_out_data_504(mau_4_io_pipe_phv_out_data_504),
    .io_pipe_phv_out_data_505(mau_4_io_pipe_phv_out_data_505),
    .io_pipe_phv_out_data_506(mau_4_io_pipe_phv_out_data_506),
    .io_pipe_phv_out_data_507(mau_4_io_pipe_phv_out_data_507),
    .io_pipe_phv_out_data_508(mau_4_io_pipe_phv_out_data_508),
    .io_pipe_phv_out_data_509(mau_4_io_pipe_phv_out_data_509),
    .io_pipe_phv_out_data_510(mau_4_io_pipe_phv_out_data_510),
    .io_pipe_phv_out_data_511(mau_4_io_pipe_phv_out_data_511),
    .io_pipe_phv_out_header_0(mau_4_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(mau_4_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(mau_4_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(mau_4_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(mau_4_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(mau_4_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(mau_4_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(mau_4_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(mau_4_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(mau_4_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(mau_4_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(mau_4_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(mau_4_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(mau_4_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(mau_4_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(mau_4_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(mau_4_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(mau_4_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(mau_4_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(mau_4_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(mau_4_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(mau_4_io_pipe_phv_out_is_valid_processor),
    .io_mod_state_id_mod(mau_4_io_mod_state_id_mod),
    .io_mod_state_id(mau_4_io_mod_state_id),
    .io_mod_sram_w_cs(mau_4_io_mod_sram_w_cs),
    .io_mod_sram_w_en(mau_4_io_mod_sram_w_en),
    .io_mod_sram_w_addr(mau_4_io_mod_sram_w_addr),
    .io_mod_sram_w_data(mau_4_io_mod_sram_w_data)
  );
  ParseModule mau_5 ( // @[parser_pisa.scala 31:25]
    .clock(mau_5_clock),
    .io_pipe_phv_in_data_0(mau_5_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(mau_5_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(mau_5_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(mau_5_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(mau_5_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(mau_5_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(mau_5_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(mau_5_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(mau_5_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(mau_5_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(mau_5_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(mau_5_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(mau_5_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(mau_5_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(mau_5_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(mau_5_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(mau_5_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(mau_5_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(mau_5_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(mau_5_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(mau_5_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(mau_5_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(mau_5_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(mau_5_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(mau_5_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(mau_5_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(mau_5_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(mau_5_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(mau_5_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(mau_5_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(mau_5_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(mau_5_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(mau_5_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(mau_5_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(mau_5_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(mau_5_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(mau_5_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(mau_5_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(mau_5_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(mau_5_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(mau_5_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(mau_5_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(mau_5_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(mau_5_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(mau_5_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(mau_5_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(mau_5_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(mau_5_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(mau_5_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(mau_5_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(mau_5_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(mau_5_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(mau_5_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(mau_5_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(mau_5_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(mau_5_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(mau_5_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(mau_5_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(mau_5_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(mau_5_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(mau_5_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(mau_5_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(mau_5_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(mau_5_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(mau_5_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(mau_5_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(mau_5_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(mau_5_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(mau_5_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(mau_5_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(mau_5_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(mau_5_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(mau_5_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(mau_5_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(mau_5_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(mau_5_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(mau_5_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(mau_5_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(mau_5_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(mau_5_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(mau_5_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(mau_5_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(mau_5_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(mau_5_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(mau_5_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(mau_5_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(mau_5_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(mau_5_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(mau_5_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(mau_5_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(mau_5_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(mau_5_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(mau_5_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(mau_5_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(mau_5_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(mau_5_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(mau_5_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(mau_5_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(mau_5_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(mau_5_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(mau_5_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(mau_5_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(mau_5_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(mau_5_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(mau_5_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(mau_5_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(mau_5_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(mau_5_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(mau_5_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(mau_5_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(mau_5_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(mau_5_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(mau_5_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(mau_5_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(mau_5_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(mau_5_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(mau_5_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(mau_5_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(mau_5_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(mau_5_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(mau_5_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(mau_5_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(mau_5_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(mau_5_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(mau_5_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(mau_5_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(mau_5_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(mau_5_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(mau_5_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(mau_5_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(mau_5_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(mau_5_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(mau_5_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(mau_5_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(mau_5_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(mau_5_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(mau_5_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(mau_5_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(mau_5_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(mau_5_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(mau_5_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(mau_5_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(mau_5_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(mau_5_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(mau_5_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(mau_5_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(mau_5_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(mau_5_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(mau_5_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(mau_5_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(mau_5_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(mau_5_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(mau_5_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(mau_5_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(mau_5_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(mau_5_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(mau_5_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(mau_5_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(mau_5_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(mau_5_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(mau_5_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(mau_5_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(mau_5_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(mau_5_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(mau_5_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(mau_5_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(mau_5_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(mau_5_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(mau_5_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(mau_5_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(mau_5_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(mau_5_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(mau_5_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(mau_5_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(mau_5_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(mau_5_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(mau_5_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(mau_5_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(mau_5_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(mau_5_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(mau_5_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(mau_5_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(mau_5_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(mau_5_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(mau_5_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(mau_5_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(mau_5_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(mau_5_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(mau_5_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(mau_5_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(mau_5_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(mau_5_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(mau_5_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(mau_5_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(mau_5_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(mau_5_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(mau_5_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(mau_5_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(mau_5_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(mau_5_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(mau_5_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(mau_5_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(mau_5_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(mau_5_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(mau_5_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(mau_5_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(mau_5_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(mau_5_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(mau_5_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(mau_5_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(mau_5_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(mau_5_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(mau_5_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(mau_5_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(mau_5_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(mau_5_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(mau_5_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(mau_5_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(mau_5_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(mau_5_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(mau_5_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(mau_5_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(mau_5_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(mau_5_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(mau_5_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(mau_5_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(mau_5_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(mau_5_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(mau_5_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(mau_5_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(mau_5_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(mau_5_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(mau_5_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(mau_5_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(mau_5_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(mau_5_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(mau_5_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(mau_5_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(mau_5_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(mau_5_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(mau_5_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(mau_5_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(mau_5_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(mau_5_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(mau_5_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(mau_5_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(mau_5_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(mau_5_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(mau_5_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(mau_5_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(mau_5_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(mau_5_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(mau_5_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(mau_5_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(mau_5_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(mau_5_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_data_256(mau_5_io_pipe_phv_in_data_256),
    .io_pipe_phv_in_data_257(mau_5_io_pipe_phv_in_data_257),
    .io_pipe_phv_in_data_258(mau_5_io_pipe_phv_in_data_258),
    .io_pipe_phv_in_data_259(mau_5_io_pipe_phv_in_data_259),
    .io_pipe_phv_in_data_260(mau_5_io_pipe_phv_in_data_260),
    .io_pipe_phv_in_data_261(mau_5_io_pipe_phv_in_data_261),
    .io_pipe_phv_in_data_262(mau_5_io_pipe_phv_in_data_262),
    .io_pipe_phv_in_data_263(mau_5_io_pipe_phv_in_data_263),
    .io_pipe_phv_in_data_264(mau_5_io_pipe_phv_in_data_264),
    .io_pipe_phv_in_data_265(mau_5_io_pipe_phv_in_data_265),
    .io_pipe_phv_in_data_266(mau_5_io_pipe_phv_in_data_266),
    .io_pipe_phv_in_data_267(mau_5_io_pipe_phv_in_data_267),
    .io_pipe_phv_in_data_268(mau_5_io_pipe_phv_in_data_268),
    .io_pipe_phv_in_data_269(mau_5_io_pipe_phv_in_data_269),
    .io_pipe_phv_in_data_270(mau_5_io_pipe_phv_in_data_270),
    .io_pipe_phv_in_data_271(mau_5_io_pipe_phv_in_data_271),
    .io_pipe_phv_in_data_272(mau_5_io_pipe_phv_in_data_272),
    .io_pipe_phv_in_data_273(mau_5_io_pipe_phv_in_data_273),
    .io_pipe_phv_in_data_274(mau_5_io_pipe_phv_in_data_274),
    .io_pipe_phv_in_data_275(mau_5_io_pipe_phv_in_data_275),
    .io_pipe_phv_in_data_276(mau_5_io_pipe_phv_in_data_276),
    .io_pipe_phv_in_data_277(mau_5_io_pipe_phv_in_data_277),
    .io_pipe_phv_in_data_278(mau_5_io_pipe_phv_in_data_278),
    .io_pipe_phv_in_data_279(mau_5_io_pipe_phv_in_data_279),
    .io_pipe_phv_in_data_280(mau_5_io_pipe_phv_in_data_280),
    .io_pipe_phv_in_data_281(mau_5_io_pipe_phv_in_data_281),
    .io_pipe_phv_in_data_282(mau_5_io_pipe_phv_in_data_282),
    .io_pipe_phv_in_data_283(mau_5_io_pipe_phv_in_data_283),
    .io_pipe_phv_in_data_284(mau_5_io_pipe_phv_in_data_284),
    .io_pipe_phv_in_data_285(mau_5_io_pipe_phv_in_data_285),
    .io_pipe_phv_in_data_286(mau_5_io_pipe_phv_in_data_286),
    .io_pipe_phv_in_data_287(mau_5_io_pipe_phv_in_data_287),
    .io_pipe_phv_in_data_288(mau_5_io_pipe_phv_in_data_288),
    .io_pipe_phv_in_data_289(mau_5_io_pipe_phv_in_data_289),
    .io_pipe_phv_in_data_290(mau_5_io_pipe_phv_in_data_290),
    .io_pipe_phv_in_data_291(mau_5_io_pipe_phv_in_data_291),
    .io_pipe_phv_in_data_292(mau_5_io_pipe_phv_in_data_292),
    .io_pipe_phv_in_data_293(mau_5_io_pipe_phv_in_data_293),
    .io_pipe_phv_in_data_294(mau_5_io_pipe_phv_in_data_294),
    .io_pipe_phv_in_data_295(mau_5_io_pipe_phv_in_data_295),
    .io_pipe_phv_in_data_296(mau_5_io_pipe_phv_in_data_296),
    .io_pipe_phv_in_data_297(mau_5_io_pipe_phv_in_data_297),
    .io_pipe_phv_in_data_298(mau_5_io_pipe_phv_in_data_298),
    .io_pipe_phv_in_data_299(mau_5_io_pipe_phv_in_data_299),
    .io_pipe_phv_in_data_300(mau_5_io_pipe_phv_in_data_300),
    .io_pipe_phv_in_data_301(mau_5_io_pipe_phv_in_data_301),
    .io_pipe_phv_in_data_302(mau_5_io_pipe_phv_in_data_302),
    .io_pipe_phv_in_data_303(mau_5_io_pipe_phv_in_data_303),
    .io_pipe_phv_in_data_304(mau_5_io_pipe_phv_in_data_304),
    .io_pipe_phv_in_data_305(mau_5_io_pipe_phv_in_data_305),
    .io_pipe_phv_in_data_306(mau_5_io_pipe_phv_in_data_306),
    .io_pipe_phv_in_data_307(mau_5_io_pipe_phv_in_data_307),
    .io_pipe_phv_in_data_308(mau_5_io_pipe_phv_in_data_308),
    .io_pipe_phv_in_data_309(mau_5_io_pipe_phv_in_data_309),
    .io_pipe_phv_in_data_310(mau_5_io_pipe_phv_in_data_310),
    .io_pipe_phv_in_data_311(mau_5_io_pipe_phv_in_data_311),
    .io_pipe_phv_in_data_312(mau_5_io_pipe_phv_in_data_312),
    .io_pipe_phv_in_data_313(mau_5_io_pipe_phv_in_data_313),
    .io_pipe_phv_in_data_314(mau_5_io_pipe_phv_in_data_314),
    .io_pipe_phv_in_data_315(mau_5_io_pipe_phv_in_data_315),
    .io_pipe_phv_in_data_316(mau_5_io_pipe_phv_in_data_316),
    .io_pipe_phv_in_data_317(mau_5_io_pipe_phv_in_data_317),
    .io_pipe_phv_in_data_318(mau_5_io_pipe_phv_in_data_318),
    .io_pipe_phv_in_data_319(mau_5_io_pipe_phv_in_data_319),
    .io_pipe_phv_in_data_320(mau_5_io_pipe_phv_in_data_320),
    .io_pipe_phv_in_data_321(mau_5_io_pipe_phv_in_data_321),
    .io_pipe_phv_in_data_322(mau_5_io_pipe_phv_in_data_322),
    .io_pipe_phv_in_data_323(mau_5_io_pipe_phv_in_data_323),
    .io_pipe_phv_in_data_324(mau_5_io_pipe_phv_in_data_324),
    .io_pipe_phv_in_data_325(mau_5_io_pipe_phv_in_data_325),
    .io_pipe_phv_in_data_326(mau_5_io_pipe_phv_in_data_326),
    .io_pipe_phv_in_data_327(mau_5_io_pipe_phv_in_data_327),
    .io_pipe_phv_in_data_328(mau_5_io_pipe_phv_in_data_328),
    .io_pipe_phv_in_data_329(mau_5_io_pipe_phv_in_data_329),
    .io_pipe_phv_in_data_330(mau_5_io_pipe_phv_in_data_330),
    .io_pipe_phv_in_data_331(mau_5_io_pipe_phv_in_data_331),
    .io_pipe_phv_in_data_332(mau_5_io_pipe_phv_in_data_332),
    .io_pipe_phv_in_data_333(mau_5_io_pipe_phv_in_data_333),
    .io_pipe_phv_in_data_334(mau_5_io_pipe_phv_in_data_334),
    .io_pipe_phv_in_data_335(mau_5_io_pipe_phv_in_data_335),
    .io_pipe_phv_in_data_336(mau_5_io_pipe_phv_in_data_336),
    .io_pipe_phv_in_data_337(mau_5_io_pipe_phv_in_data_337),
    .io_pipe_phv_in_data_338(mau_5_io_pipe_phv_in_data_338),
    .io_pipe_phv_in_data_339(mau_5_io_pipe_phv_in_data_339),
    .io_pipe_phv_in_data_340(mau_5_io_pipe_phv_in_data_340),
    .io_pipe_phv_in_data_341(mau_5_io_pipe_phv_in_data_341),
    .io_pipe_phv_in_data_342(mau_5_io_pipe_phv_in_data_342),
    .io_pipe_phv_in_data_343(mau_5_io_pipe_phv_in_data_343),
    .io_pipe_phv_in_data_344(mau_5_io_pipe_phv_in_data_344),
    .io_pipe_phv_in_data_345(mau_5_io_pipe_phv_in_data_345),
    .io_pipe_phv_in_data_346(mau_5_io_pipe_phv_in_data_346),
    .io_pipe_phv_in_data_347(mau_5_io_pipe_phv_in_data_347),
    .io_pipe_phv_in_data_348(mau_5_io_pipe_phv_in_data_348),
    .io_pipe_phv_in_data_349(mau_5_io_pipe_phv_in_data_349),
    .io_pipe_phv_in_data_350(mau_5_io_pipe_phv_in_data_350),
    .io_pipe_phv_in_data_351(mau_5_io_pipe_phv_in_data_351),
    .io_pipe_phv_in_data_352(mau_5_io_pipe_phv_in_data_352),
    .io_pipe_phv_in_data_353(mau_5_io_pipe_phv_in_data_353),
    .io_pipe_phv_in_data_354(mau_5_io_pipe_phv_in_data_354),
    .io_pipe_phv_in_data_355(mau_5_io_pipe_phv_in_data_355),
    .io_pipe_phv_in_data_356(mau_5_io_pipe_phv_in_data_356),
    .io_pipe_phv_in_data_357(mau_5_io_pipe_phv_in_data_357),
    .io_pipe_phv_in_data_358(mau_5_io_pipe_phv_in_data_358),
    .io_pipe_phv_in_data_359(mau_5_io_pipe_phv_in_data_359),
    .io_pipe_phv_in_data_360(mau_5_io_pipe_phv_in_data_360),
    .io_pipe_phv_in_data_361(mau_5_io_pipe_phv_in_data_361),
    .io_pipe_phv_in_data_362(mau_5_io_pipe_phv_in_data_362),
    .io_pipe_phv_in_data_363(mau_5_io_pipe_phv_in_data_363),
    .io_pipe_phv_in_data_364(mau_5_io_pipe_phv_in_data_364),
    .io_pipe_phv_in_data_365(mau_5_io_pipe_phv_in_data_365),
    .io_pipe_phv_in_data_366(mau_5_io_pipe_phv_in_data_366),
    .io_pipe_phv_in_data_367(mau_5_io_pipe_phv_in_data_367),
    .io_pipe_phv_in_data_368(mau_5_io_pipe_phv_in_data_368),
    .io_pipe_phv_in_data_369(mau_5_io_pipe_phv_in_data_369),
    .io_pipe_phv_in_data_370(mau_5_io_pipe_phv_in_data_370),
    .io_pipe_phv_in_data_371(mau_5_io_pipe_phv_in_data_371),
    .io_pipe_phv_in_data_372(mau_5_io_pipe_phv_in_data_372),
    .io_pipe_phv_in_data_373(mau_5_io_pipe_phv_in_data_373),
    .io_pipe_phv_in_data_374(mau_5_io_pipe_phv_in_data_374),
    .io_pipe_phv_in_data_375(mau_5_io_pipe_phv_in_data_375),
    .io_pipe_phv_in_data_376(mau_5_io_pipe_phv_in_data_376),
    .io_pipe_phv_in_data_377(mau_5_io_pipe_phv_in_data_377),
    .io_pipe_phv_in_data_378(mau_5_io_pipe_phv_in_data_378),
    .io_pipe_phv_in_data_379(mau_5_io_pipe_phv_in_data_379),
    .io_pipe_phv_in_data_380(mau_5_io_pipe_phv_in_data_380),
    .io_pipe_phv_in_data_381(mau_5_io_pipe_phv_in_data_381),
    .io_pipe_phv_in_data_382(mau_5_io_pipe_phv_in_data_382),
    .io_pipe_phv_in_data_383(mau_5_io_pipe_phv_in_data_383),
    .io_pipe_phv_in_data_384(mau_5_io_pipe_phv_in_data_384),
    .io_pipe_phv_in_data_385(mau_5_io_pipe_phv_in_data_385),
    .io_pipe_phv_in_data_386(mau_5_io_pipe_phv_in_data_386),
    .io_pipe_phv_in_data_387(mau_5_io_pipe_phv_in_data_387),
    .io_pipe_phv_in_data_388(mau_5_io_pipe_phv_in_data_388),
    .io_pipe_phv_in_data_389(mau_5_io_pipe_phv_in_data_389),
    .io_pipe_phv_in_data_390(mau_5_io_pipe_phv_in_data_390),
    .io_pipe_phv_in_data_391(mau_5_io_pipe_phv_in_data_391),
    .io_pipe_phv_in_data_392(mau_5_io_pipe_phv_in_data_392),
    .io_pipe_phv_in_data_393(mau_5_io_pipe_phv_in_data_393),
    .io_pipe_phv_in_data_394(mau_5_io_pipe_phv_in_data_394),
    .io_pipe_phv_in_data_395(mau_5_io_pipe_phv_in_data_395),
    .io_pipe_phv_in_data_396(mau_5_io_pipe_phv_in_data_396),
    .io_pipe_phv_in_data_397(mau_5_io_pipe_phv_in_data_397),
    .io_pipe_phv_in_data_398(mau_5_io_pipe_phv_in_data_398),
    .io_pipe_phv_in_data_399(mau_5_io_pipe_phv_in_data_399),
    .io_pipe_phv_in_data_400(mau_5_io_pipe_phv_in_data_400),
    .io_pipe_phv_in_data_401(mau_5_io_pipe_phv_in_data_401),
    .io_pipe_phv_in_data_402(mau_5_io_pipe_phv_in_data_402),
    .io_pipe_phv_in_data_403(mau_5_io_pipe_phv_in_data_403),
    .io_pipe_phv_in_data_404(mau_5_io_pipe_phv_in_data_404),
    .io_pipe_phv_in_data_405(mau_5_io_pipe_phv_in_data_405),
    .io_pipe_phv_in_data_406(mau_5_io_pipe_phv_in_data_406),
    .io_pipe_phv_in_data_407(mau_5_io_pipe_phv_in_data_407),
    .io_pipe_phv_in_data_408(mau_5_io_pipe_phv_in_data_408),
    .io_pipe_phv_in_data_409(mau_5_io_pipe_phv_in_data_409),
    .io_pipe_phv_in_data_410(mau_5_io_pipe_phv_in_data_410),
    .io_pipe_phv_in_data_411(mau_5_io_pipe_phv_in_data_411),
    .io_pipe_phv_in_data_412(mau_5_io_pipe_phv_in_data_412),
    .io_pipe_phv_in_data_413(mau_5_io_pipe_phv_in_data_413),
    .io_pipe_phv_in_data_414(mau_5_io_pipe_phv_in_data_414),
    .io_pipe_phv_in_data_415(mau_5_io_pipe_phv_in_data_415),
    .io_pipe_phv_in_data_416(mau_5_io_pipe_phv_in_data_416),
    .io_pipe_phv_in_data_417(mau_5_io_pipe_phv_in_data_417),
    .io_pipe_phv_in_data_418(mau_5_io_pipe_phv_in_data_418),
    .io_pipe_phv_in_data_419(mau_5_io_pipe_phv_in_data_419),
    .io_pipe_phv_in_data_420(mau_5_io_pipe_phv_in_data_420),
    .io_pipe_phv_in_data_421(mau_5_io_pipe_phv_in_data_421),
    .io_pipe_phv_in_data_422(mau_5_io_pipe_phv_in_data_422),
    .io_pipe_phv_in_data_423(mau_5_io_pipe_phv_in_data_423),
    .io_pipe_phv_in_data_424(mau_5_io_pipe_phv_in_data_424),
    .io_pipe_phv_in_data_425(mau_5_io_pipe_phv_in_data_425),
    .io_pipe_phv_in_data_426(mau_5_io_pipe_phv_in_data_426),
    .io_pipe_phv_in_data_427(mau_5_io_pipe_phv_in_data_427),
    .io_pipe_phv_in_data_428(mau_5_io_pipe_phv_in_data_428),
    .io_pipe_phv_in_data_429(mau_5_io_pipe_phv_in_data_429),
    .io_pipe_phv_in_data_430(mau_5_io_pipe_phv_in_data_430),
    .io_pipe_phv_in_data_431(mau_5_io_pipe_phv_in_data_431),
    .io_pipe_phv_in_data_432(mau_5_io_pipe_phv_in_data_432),
    .io_pipe_phv_in_data_433(mau_5_io_pipe_phv_in_data_433),
    .io_pipe_phv_in_data_434(mau_5_io_pipe_phv_in_data_434),
    .io_pipe_phv_in_data_435(mau_5_io_pipe_phv_in_data_435),
    .io_pipe_phv_in_data_436(mau_5_io_pipe_phv_in_data_436),
    .io_pipe_phv_in_data_437(mau_5_io_pipe_phv_in_data_437),
    .io_pipe_phv_in_data_438(mau_5_io_pipe_phv_in_data_438),
    .io_pipe_phv_in_data_439(mau_5_io_pipe_phv_in_data_439),
    .io_pipe_phv_in_data_440(mau_5_io_pipe_phv_in_data_440),
    .io_pipe_phv_in_data_441(mau_5_io_pipe_phv_in_data_441),
    .io_pipe_phv_in_data_442(mau_5_io_pipe_phv_in_data_442),
    .io_pipe_phv_in_data_443(mau_5_io_pipe_phv_in_data_443),
    .io_pipe_phv_in_data_444(mau_5_io_pipe_phv_in_data_444),
    .io_pipe_phv_in_data_445(mau_5_io_pipe_phv_in_data_445),
    .io_pipe_phv_in_data_446(mau_5_io_pipe_phv_in_data_446),
    .io_pipe_phv_in_data_447(mau_5_io_pipe_phv_in_data_447),
    .io_pipe_phv_in_data_448(mau_5_io_pipe_phv_in_data_448),
    .io_pipe_phv_in_data_449(mau_5_io_pipe_phv_in_data_449),
    .io_pipe_phv_in_data_450(mau_5_io_pipe_phv_in_data_450),
    .io_pipe_phv_in_data_451(mau_5_io_pipe_phv_in_data_451),
    .io_pipe_phv_in_data_452(mau_5_io_pipe_phv_in_data_452),
    .io_pipe_phv_in_data_453(mau_5_io_pipe_phv_in_data_453),
    .io_pipe_phv_in_data_454(mau_5_io_pipe_phv_in_data_454),
    .io_pipe_phv_in_data_455(mau_5_io_pipe_phv_in_data_455),
    .io_pipe_phv_in_data_456(mau_5_io_pipe_phv_in_data_456),
    .io_pipe_phv_in_data_457(mau_5_io_pipe_phv_in_data_457),
    .io_pipe_phv_in_data_458(mau_5_io_pipe_phv_in_data_458),
    .io_pipe_phv_in_data_459(mau_5_io_pipe_phv_in_data_459),
    .io_pipe_phv_in_data_460(mau_5_io_pipe_phv_in_data_460),
    .io_pipe_phv_in_data_461(mau_5_io_pipe_phv_in_data_461),
    .io_pipe_phv_in_data_462(mau_5_io_pipe_phv_in_data_462),
    .io_pipe_phv_in_data_463(mau_5_io_pipe_phv_in_data_463),
    .io_pipe_phv_in_data_464(mau_5_io_pipe_phv_in_data_464),
    .io_pipe_phv_in_data_465(mau_5_io_pipe_phv_in_data_465),
    .io_pipe_phv_in_data_466(mau_5_io_pipe_phv_in_data_466),
    .io_pipe_phv_in_data_467(mau_5_io_pipe_phv_in_data_467),
    .io_pipe_phv_in_data_468(mau_5_io_pipe_phv_in_data_468),
    .io_pipe_phv_in_data_469(mau_5_io_pipe_phv_in_data_469),
    .io_pipe_phv_in_data_470(mau_5_io_pipe_phv_in_data_470),
    .io_pipe_phv_in_data_471(mau_5_io_pipe_phv_in_data_471),
    .io_pipe_phv_in_data_472(mau_5_io_pipe_phv_in_data_472),
    .io_pipe_phv_in_data_473(mau_5_io_pipe_phv_in_data_473),
    .io_pipe_phv_in_data_474(mau_5_io_pipe_phv_in_data_474),
    .io_pipe_phv_in_data_475(mau_5_io_pipe_phv_in_data_475),
    .io_pipe_phv_in_data_476(mau_5_io_pipe_phv_in_data_476),
    .io_pipe_phv_in_data_477(mau_5_io_pipe_phv_in_data_477),
    .io_pipe_phv_in_data_478(mau_5_io_pipe_phv_in_data_478),
    .io_pipe_phv_in_data_479(mau_5_io_pipe_phv_in_data_479),
    .io_pipe_phv_in_data_480(mau_5_io_pipe_phv_in_data_480),
    .io_pipe_phv_in_data_481(mau_5_io_pipe_phv_in_data_481),
    .io_pipe_phv_in_data_482(mau_5_io_pipe_phv_in_data_482),
    .io_pipe_phv_in_data_483(mau_5_io_pipe_phv_in_data_483),
    .io_pipe_phv_in_data_484(mau_5_io_pipe_phv_in_data_484),
    .io_pipe_phv_in_data_485(mau_5_io_pipe_phv_in_data_485),
    .io_pipe_phv_in_data_486(mau_5_io_pipe_phv_in_data_486),
    .io_pipe_phv_in_data_487(mau_5_io_pipe_phv_in_data_487),
    .io_pipe_phv_in_data_488(mau_5_io_pipe_phv_in_data_488),
    .io_pipe_phv_in_data_489(mau_5_io_pipe_phv_in_data_489),
    .io_pipe_phv_in_data_490(mau_5_io_pipe_phv_in_data_490),
    .io_pipe_phv_in_data_491(mau_5_io_pipe_phv_in_data_491),
    .io_pipe_phv_in_data_492(mau_5_io_pipe_phv_in_data_492),
    .io_pipe_phv_in_data_493(mau_5_io_pipe_phv_in_data_493),
    .io_pipe_phv_in_data_494(mau_5_io_pipe_phv_in_data_494),
    .io_pipe_phv_in_data_495(mau_5_io_pipe_phv_in_data_495),
    .io_pipe_phv_in_data_496(mau_5_io_pipe_phv_in_data_496),
    .io_pipe_phv_in_data_497(mau_5_io_pipe_phv_in_data_497),
    .io_pipe_phv_in_data_498(mau_5_io_pipe_phv_in_data_498),
    .io_pipe_phv_in_data_499(mau_5_io_pipe_phv_in_data_499),
    .io_pipe_phv_in_data_500(mau_5_io_pipe_phv_in_data_500),
    .io_pipe_phv_in_data_501(mau_5_io_pipe_phv_in_data_501),
    .io_pipe_phv_in_data_502(mau_5_io_pipe_phv_in_data_502),
    .io_pipe_phv_in_data_503(mau_5_io_pipe_phv_in_data_503),
    .io_pipe_phv_in_data_504(mau_5_io_pipe_phv_in_data_504),
    .io_pipe_phv_in_data_505(mau_5_io_pipe_phv_in_data_505),
    .io_pipe_phv_in_data_506(mau_5_io_pipe_phv_in_data_506),
    .io_pipe_phv_in_data_507(mau_5_io_pipe_phv_in_data_507),
    .io_pipe_phv_in_data_508(mau_5_io_pipe_phv_in_data_508),
    .io_pipe_phv_in_data_509(mau_5_io_pipe_phv_in_data_509),
    .io_pipe_phv_in_data_510(mau_5_io_pipe_phv_in_data_510),
    .io_pipe_phv_in_data_511(mau_5_io_pipe_phv_in_data_511),
    .io_pipe_phv_in_header_0(mau_5_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(mau_5_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(mau_5_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(mau_5_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(mau_5_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(mau_5_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(mau_5_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(mau_5_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(mau_5_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(mau_5_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(mau_5_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(mau_5_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(mau_5_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(mau_5_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(mau_5_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(mau_5_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(mau_5_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(mau_5_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(mau_5_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(mau_5_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(mau_5_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(mau_5_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(mau_5_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(mau_5_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(mau_5_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(mau_5_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(mau_5_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(mau_5_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(mau_5_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(mau_5_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(mau_5_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(mau_5_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(mau_5_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(mau_5_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(mau_5_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(mau_5_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(mau_5_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(mau_5_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(mau_5_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(mau_5_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(mau_5_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(mau_5_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(mau_5_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(mau_5_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(mau_5_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(mau_5_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(mau_5_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(mau_5_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(mau_5_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(mau_5_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(mau_5_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(mau_5_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(mau_5_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(mau_5_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(mau_5_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(mau_5_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(mau_5_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(mau_5_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(mau_5_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(mau_5_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(mau_5_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(mau_5_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(mau_5_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(mau_5_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(mau_5_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(mau_5_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(mau_5_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(mau_5_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(mau_5_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(mau_5_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(mau_5_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(mau_5_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(mau_5_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(mau_5_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(mau_5_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(mau_5_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(mau_5_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(mau_5_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(mau_5_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(mau_5_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(mau_5_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(mau_5_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(mau_5_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(mau_5_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(mau_5_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(mau_5_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(mau_5_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(mau_5_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(mau_5_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(mau_5_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(mau_5_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(mau_5_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(mau_5_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(mau_5_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(mau_5_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(mau_5_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(mau_5_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(mau_5_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(mau_5_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(mau_5_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(mau_5_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(mau_5_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(mau_5_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(mau_5_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(mau_5_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(mau_5_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(mau_5_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(mau_5_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(mau_5_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(mau_5_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(mau_5_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(mau_5_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(mau_5_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(mau_5_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(mau_5_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(mau_5_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(mau_5_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(mau_5_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(mau_5_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(mau_5_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(mau_5_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(mau_5_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(mau_5_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(mau_5_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(mau_5_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(mau_5_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(mau_5_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(mau_5_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(mau_5_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(mau_5_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(mau_5_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(mau_5_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(mau_5_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(mau_5_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(mau_5_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(mau_5_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(mau_5_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(mau_5_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(mau_5_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(mau_5_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(mau_5_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(mau_5_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(mau_5_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(mau_5_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(mau_5_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(mau_5_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(mau_5_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(mau_5_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(mau_5_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(mau_5_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(mau_5_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(mau_5_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(mau_5_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(mau_5_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(mau_5_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(mau_5_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(mau_5_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(mau_5_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(mau_5_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(mau_5_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(mau_5_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(mau_5_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(mau_5_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(mau_5_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(mau_5_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(mau_5_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(mau_5_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(mau_5_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(mau_5_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(mau_5_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(mau_5_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(mau_5_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(mau_5_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(mau_5_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(mau_5_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(mau_5_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(mau_5_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(mau_5_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(mau_5_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(mau_5_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(mau_5_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(mau_5_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(mau_5_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(mau_5_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(mau_5_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(mau_5_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(mau_5_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(mau_5_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(mau_5_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(mau_5_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(mau_5_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(mau_5_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(mau_5_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(mau_5_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(mau_5_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(mau_5_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(mau_5_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(mau_5_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(mau_5_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(mau_5_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(mau_5_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(mau_5_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(mau_5_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(mau_5_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(mau_5_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(mau_5_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(mau_5_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(mau_5_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(mau_5_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(mau_5_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(mau_5_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(mau_5_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(mau_5_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(mau_5_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(mau_5_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(mau_5_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(mau_5_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(mau_5_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(mau_5_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(mau_5_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(mau_5_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(mau_5_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(mau_5_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(mau_5_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(mau_5_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(mau_5_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(mau_5_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(mau_5_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(mau_5_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(mau_5_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(mau_5_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(mau_5_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(mau_5_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(mau_5_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(mau_5_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(mau_5_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(mau_5_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(mau_5_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(mau_5_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(mau_5_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(mau_5_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(mau_5_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(mau_5_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(mau_5_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(mau_5_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(mau_5_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(mau_5_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(mau_5_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(mau_5_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(mau_5_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(mau_5_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(mau_5_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(mau_5_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(mau_5_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(mau_5_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(mau_5_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(mau_5_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(mau_5_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(mau_5_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(mau_5_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(mau_5_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(mau_5_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(mau_5_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(mau_5_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(mau_5_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(mau_5_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(mau_5_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(mau_5_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(mau_5_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(mau_5_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(mau_5_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(mau_5_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(mau_5_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(mau_5_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(mau_5_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(mau_5_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(mau_5_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(mau_5_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_data_256(mau_5_io_pipe_phv_out_data_256),
    .io_pipe_phv_out_data_257(mau_5_io_pipe_phv_out_data_257),
    .io_pipe_phv_out_data_258(mau_5_io_pipe_phv_out_data_258),
    .io_pipe_phv_out_data_259(mau_5_io_pipe_phv_out_data_259),
    .io_pipe_phv_out_data_260(mau_5_io_pipe_phv_out_data_260),
    .io_pipe_phv_out_data_261(mau_5_io_pipe_phv_out_data_261),
    .io_pipe_phv_out_data_262(mau_5_io_pipe_phv_out_data_262),
    .io_pipe_phv_out_data_263(mau_5_io_pipe_phv_out_data_263),
    .io_pipe_phv_out_data_264(mau_5_io_pipe_phv_out_data_264),
    .io_pipe_phv_out_data_265(mau_5_io_pipe_phv_out_data_265),
    .io_pipe_phv_out_data_266(mau_5_io_pipe_phv_out_data_266),
    .io_pipe_phv_out_data_267(mau_5_io_pipe_phv_out_data_267),
    .io_pipe_phv_out_data_268(mau_5_io_pipe_phv_out_data_268),
    .io_pipe_phv_out_data_269(mau_5_io_pipe_phv_out_data_269),
    .io_pipe_phv_out_data_270(mau_5_io_pipe_phv_out_data_270),
    .io_pipe_phv_out_data_271(mau_5_io_pipe_phv_out_data_271),
    .io_pipe_phv_out_data_272(mau_5_io_pipe_phv_out_data_272),
    .io_pipe_phv_out_data_273(mau_5_io_pipe_phv_out_data_273),
    .io_pipe_phv_out_data_274(mau_5_io_pipe_phv_out_data_274),
    .io_pipe_phv_out_data_275(mau_5_io_pipe_phv_out_data_275),
    .io_pipe_phv_out_data_276(mau_5_io_pipe_phv_out_data_276),
    .io_pipe_phv_out_data_277(mau_5_io_pipe_phv_out_data_277),
    .io_pipe_phv_out_data_278(mau_5_io_pipe_phv_out_data_278),
    .io_pipe_phv_out_data_279(mau_5_io_pipe_phv_out_data_279),
    .io_pipe_phv_out_data_280(mau_5_io_pipe_phv_out_data_280),
    .io_pipe_phv_out_data_281(mau_5_io_pipe_phv_out_data_281),
    .io_pipe_phv_out_data_282(mau_5_io_pipe_phv_out_data_282),
    .io_pipe_phv_out_data_283(mau_5_io_pipe_phv_out_data_283),
    .io_pipe_phv_out_data_284(mau_5_io_pipe_phv_out_data_284),
    .io_pipe_phv_out_data_285(mau_5_io_pipe_phv_out_data_285),
    .io_pipe_phv_out_data_286(mau_5_io_pipe_phv_out_data_286),
    .io_pipe_phv_out_data_287(mau_5_io_pipe_phv_out_data_287),
    .io_pipe_phv_out_data_288(mau_5_io_pipe_phv_out_data_288),
    .io_pipe_phv_out_data_289(mau_5_io_pipe_phv_out_data_289),
    .io_pipe_phv_out_data_290(mau_5_io_pipe_phv_out_data_290),
    .io_pipe_phv_out_data_291(mau_5_io_pipe_phv_out_data_291),
    .io_pipe_phv_out_data_292(mau_5_io_pipe_phv_out_data_292),
    .io_pipe_phv_out_data_293(mau_5_io_pipe_phv_out_data_293),
    .io_pipe_phv_out_data_294(mau_5_io_pipe_phv_out_data_294),
    .io_pipe_phv_out_data_295(mau_5_io_pipe_phv_out_data_295),
    .io_pipe_phv_out_data_296(mau_5_io_pipe_phv_out_data_296),
    .io_pipe_phv_out_data_297(mau_5_io_pipe_phv_out_data_297),
    .io_pipe_phv_out_data_298(mau_5_io_pipe_phv_out_data_298),
    .io_pipe_phv_out_data_299(mau_5_io_pipe_phv_out_data_299),
    .io_pipe_phv_out_data_300(mau_5_io_pipe_phv_out_data_300),
    .io_pipe_phv_out_data_301(mau_5_io_pipe_phv_out_data_301),
    .io_pipe_phv_out_data_302(mau_5_io_pipe_phv_out_data_302),
    .io_pipe_phv_out_data_303(mau_5_io_pipe_phv_out_data_303),
    .io_pipe_phv_out_data_304(mau_5_io_pipe_phv_out_data_304),
    .io_pipe_phv_out_data_305(mau_5_io_pipe_phv_out_data_305),
    .io_pipe_phv_out_data_306(mau_5_io_pipe_phv_out_data_306),
    .io_pipe_phv_out_data_307(mau_5_io_pipe_phv_out_data_307),
    .io_pipe_phv_out_data_308(mau_5_io_pipe_phv_out_data_308),
    .io_pipe_phv_out_data_309(mau_5_io_pipe_phv_out_data_309),
    .io_pipe_phv_out_data_310(mau_5_io_pipe_phv_out_data_310),
    .io_pipe_phv_out_data_311(mau_5_io_pipe_phv_out_data_311),
    .io_pipe_phv_out_data_312(mau_5_io_pipe_phv_out_data_312),
    .io_pipe_phv_out_data_313(mau_5_io_pipe_phv_out_data_313),
    .io_pipe_phv_out_data_314(mau_5_io_pipe_phv_out_data_314),
    .io_pipe_phv_out_data_315(mau_5_io_pipe_phv_out_data_315),
    .io_pipe_phv_out_data_316(mau_5_io_pipe_phv_out_data_316),
    .io_pipe_phv_out_data_317(mau_5_io_pipe_phv_out_data_317),
    .io_pipe_phv_out_data_318(mau_5_io_pipe_phv_out_data_318),
    .io_pipe_phv_out_data_319(mau_5_io_pipe_phv_out_data_319),
    .io_pipe_phv_out_data_320(mau_5_io_pipe_phv_out_data_320),
    .io_pipe_phv_out_data_321(mau_5_io_pipe_phv_out_data_321),
    .io_pipe_phv_out_data_322(mau_5_io_pipe_phv_out_data_322),
    .io_pipe_phv_out_data_323(mau_5_io_pipe_phv_out_data_323),
    .io_pipe_phv_out_data_324(mau_5_io_pipe_phv_out_data_324),
    .io_pipe_phv_out_data_325(mau_5_io_pipe_phv_out_data_325),
    .io_pipe_phv_out_data_326(mau_5_io_pipe_phv_out_data_326),
    .io_pipe_phv_out_data_327(mau_5_io_pipe_phv_out_data_327),
    .io_pipe_phv_out_data_328(mau_5_io_pipe_phv_out_data_328),
    .io_pipe_phv_out_data_329(mau_5_io_pipe_phv_out_data_329),
    .io_pipe_phv_out_data_330(mau_5_io_pipe_phv_out_data_330),
    .io_pipe_phv_out_data_331(mau_5_io_pipe_phv_out_data_331),
    .io_pipe_phv_out_data_332(mau_5_io_pipe_phv_out_data_332),
    .io_pipe_phv_out_data_333(mau_5_io_pipe_phv_out_data_333),
    .io_pipe_phv_out_data_334(mau_5_io_pipe_phv_out_data_334),
    .io_pipe_phv_out_data_335(mau_5_io_pipe_phv_out_data_335),
    .io_pipe_phv_out_data_336(mau_5_io_pipe_phv_out_data_336),
    .io_pipe_phv_out_data_337(mau_5_io_pipe_phv_out_data_337),
    .io_pipe_phv_out_data_338(mau_5_io_pipe_phv_out_data_338),
    .io_pipe_phv_out_data_339(mau_5_io_pipe_phv_out_data_339),
    .io_pipe_phv_out_data_340(mau_5_io_pipe_phv_out_data_340),
    .io_pipe_phv_out_data_341(mau_5_io_pipe_phv_out_data_341),
    .io_pipe_phv_out_data_342(mau_5_io_pipe_phv_out_data_342),
    .io_pipe_phv_out_data_343(mau_5_io_pipe_phv_out_data_343),
    .io_pipe_phv_out_data_344(mau_5_io_pipe_phv_out_data_344),
    .io_pipe_phv_out_data_345(mau_5_io_pipe_phv_out_data_345),
    .io_pipe_phv_out_data_346(mau_5_io_pipe_phv_out_data_346),
    .io_pipe_phv_out_data_347(mau_5_io_pipe_phv_out_data_347),
    .io_pipe_phv_out_data_348(mau_5_io_pipe_phv_out_data_348),
    .io_pipe_phv_out_data_349(mau_5_io_pipe_phv_out_data_349),
    .io_pipe_phv_out_data_350(mau_5_io_pipe_phv_out_data_350),
    .io_pipe_phv_out_data_351(mau_5_io_pipe_phv_out_data_351),
    .io_pipe_phv_out_data_352(mau_5_io_pipe_phv_out_data_352),
    .io_pipe_phv_out_data_353(mau_5_io_pipe_phv_out_data_353),
    .io_pipe_phv_out_data_354(mau_5_io_pipe_phv_out_data_354),
    .io_pipe_phv_out_data_355(mau_5_io_pipe_phv_out_data_355),
    .io_pipe_phv_out_data_356(mau_5_io_pipe_phv_out_data_356),
    .io_pipe_phv_out_data_357(mau_5_io_pipe_phv_out_data_357),
    .io_pipe_phv_out_data_358(mau_5_io_pipe_phv_out_data_358),
    .io_pipe_phv_out_data_359(mau_5_io_pipe_phv_out_data_359),
    .io_pipe_phv_out_data_360(mau_5_io_pipe_phv_out_data_360),
    .io_pipe_phv_out_data_361(mau_5_io_pipe_phv_out_data_361),
    .io_pipe_phv_out_data_362(mau_5_io_pipe_phv_out_data_362),
    .io_pipe_phv_out_data_363(mau_5_io_pipe_phv_out_data_363),
    .io_pipe_phv_out_data_364(mau_5_io_pipe_phv_out_data_364),
    .io_pipe_phv_out_data_365(mau_5_io_pipe_phv_out_data_365),
    .io_pipe_phv_out_data_366(mau_5_io_pipe_phv_out_data_366),
    .io_pipe_phv_out_data_367(mau_5_io_pipe_phv_out_data_367),
    .io_pipe_phv_out_data_368(mau_5_io_pipe_phv_out_data_368),
    .io_pipe_phv_out_data_369(mau_5_io_pipe_phv_out_data_369),
    .io_pipe_phv_out_data_370(mau_5_io_pipe_phv_out_data_370),
    .io_pipe_phv_out_data_371(mau_5_io_pipe_phv_out_data_371),
    .io_pipe_phv_out_data_372(mau_5_io_pipe_phv_out_data_372),
    .io_pipe_phv_out_data_373(mau_5_io_pipe_phv_out_data_373),
    .io_pipe_phv_out_data_374(mau_5_io_pipe_phv_out_data_374),
    .io_pipe_phv_out_data_375(mau_5_io_pipe_phv_out_data_375),
    .io_pipe_phv_out_data_376(mau_5_io_pipe_phv_out_data_376),
    .io_pipe_phv_out_data_377(mau_5_io_pipe_phv_out_data_377),
    .io_pipe_phv_out_data_378(mau_5_io_pipe_phv_out_data_378),
    .io_pipe_phv_out_data_379(mau_5_io_pipe_phv_out_data_379),
    .io_pipe_phv_out_data_380(mau_5_io_pipe_phv_out_data_380),
    .io_pipe_phv_out_data_381(mau_5_io_pipe_phv_out_data_381),
    .io_pipe_phv_out_data_382(mau_5_io_pipe_phv_out_data_382),
    .io_pipe_phv_out_data_383(mau_5_io_pipe_phv_out_data_383),
    .io_pipe_phv_out_data_384(mau_5_io_pipe_phv_out_data_384),
    .io_pipe_phv_out_data_385(mau_5_io_pipe_phv_out_data_385),
    .io_pipe_phv_out_data_386(mau_5_io_pipe_phv_out_data_386),
    .io_pipe_phv_out_data_387(mau_5_io_pipe_phv_out_data_387),
    .io_pipe_phv_out_data_388(mau_5_io_pipe_phv_out_data_388),
    .io_pipe_phv_out_data_389(mau_5_io_pipe_phv_out_data_389),
    .io_pipe_phv_out_data_390(mau_5_io_pipe_phv_out_data_390),
    .io_pipe_phv_out_data_391(mau_5_io_pipe_phv_out_data_391),
    .io_pipe_phv_out_data_392(mau_5_io_pipe_phv_out_data_392),
    .io_pipe_phv_out_data_393(mau_5_io_pipe_phv_out_data_393),
    .io_pipe_phv_out_data_394(mau_5_io_pipe_phv_out_data_394),
    .io_pipe_phv_out_data_395(mau_5_io_pipe_phv_out_data_395),
    .io_pipe_phv_out_data_396(mau_5_io_pipe_phv_out_data_396),
    .io_pipe_phv_out_data_397(mau_5_io_pipe_phv_out_data_397),
    .io_pipe_phv_out_data_398(mau_5_io_pipe_phv_out_data_398),
    .io_pipe_phv_out_data_399(mau_5_io_pipe_phv_out_data_399),
    .io_pipe_phv_out_data_400(mau_5_io_pipe_phv_out_data_400),
    .io_pipe_phv_out_data_401(mau_5_io_pipe_phv_out_data_401),
    .io_pipe_phv_out_data_402(mau_5_io_pipe_phv_out_data_402),
    .io_pipe_phv_out_data_403(mau_5_io_pipe_phv_out_data_403),
    .io_pipe_phv_out_data_404(mau_5_io_pipe_phv_out_data_404),
    .io_pipe_phv_out_data_405(mau_5_io_pipe_phv_out_data_405),
    .io_pipe_phv_out_data_406(mau_5_io_pipe_phv_out_data_406),
    .io_pipe_phv_out_data_407(mau_5_io_pipe_phv_out_data_407),
    .io_pipe_phv_out_data_408(mau_5_io_pipe_phv_out_data_408),
    .io_pipe_phv_out_data_409(mau_5_io_pipe_phv_out_data_409),
    .io_pipe_phv_out_data_410(mau_5_io_pipe_phv_out_data_410),
    .io_pipe_phv_out_data_411(mau_5_io_pipe_phv_out_data_411),
    .io_pipe_phv_out_data_412(mau_5_io_pipe_phv_out_data_412),
    .io_pipe_phv_out_data_413(mau_5_io_pipe_phv_out_data_413),
    .io_pipe_phv_out_data_414(mau_5_io_pipe_phv_out_data_414),
    .io_pipe_phv_out_data_415(mau_5_io_pipe_phv_out_data_415),
    .io_pipe_phv_out_data_416(mau_5_io_pipe_phv_out_data_416),
    .io_pipe_phv_out_data_417(mau_5_io_pipe_phv_out_data_417),
    .io_pipe_phv_out_data_418(mau_5_io_pipe_phv_out_data_418),
    .io_pipe_phv_out_data_419(mau_5_io_pipe_phv_out_data_419),
    .io_pipe_phv_out_data_420(mau_5_io_pipe_phv_out_data_420),
    .io_pipe_phv_out_data_421(mau_5_io_pipe_phv_out_data_421),
    .io_pipe_phv_out_data_422(mau_5_io_pipe_phv_out_data_422),
    .io_pipe_phv_out_data_423(mau_5_io_pipe_phv_out_data_423),
    .io_pipe_phv_out_data_424(mau_5_io_pipe_phv_out_data_424),
    .io_pipe_phv_out_data_425(mau_5_io_pipe_phv_out_data_425),
    .io_pipe_phv_out_data_426(mau_5_io_pipe_phv_out_data_426),
    .io_pipe_phv_out_data_427(mau_5_io_pipe_phv_out_data_427),
    .io_pipe_phv_out_data_428(mau_5_io_pipe_phv_out_data_428),
    .io_pipe_phv_out_data_429(mau_5_io_pipe_phv_out_data_429),
    .io_pipe_phv_out_data_430(mau_5_io_pipe_phv_out_data_430),
    .io_pipe_phv_out_data_431(mau_5_io_pipe_phv_out_data_431),
    .io_pipe_phv_out_data_432(mau_5_io_pipe_phv_out_data_432),
    .io_pipe_phv_out_data_433(mau_5_io_pipe_phv_out_data_433),
    .io_pipe_phv_out_data_434(mau_5_io_pipe_phv_out_data_434),
    .io_pipe_phv_out_data_435(mau_5_io_pipe_phv_out_data_435),
    .io_pipe_phv_out_data_436(mau_5_io_pipe_phv_out_data_436),
    .io_pipe_phv_out_data_437(mau_5_io_pipe_phv_out_data_437),
    .io_pipe_phv_out_data_438(mau_5_io_pipe_phv_out_data_438),
    .io_pipe_phv_out_data_439(mau_5_io_pipe_phv_out_data_439),
    .io_pipe_phv_out_data_440(mau_5_io_pipe_phv_out_data_440),
    .io_pipe_phv_out_data_441(mau_5_io_pipe_phv_out_data_441),
    .io_pipe_phv_out_data_442(mau_5_io_pipe_phv_out_data_442),
    .io_pipe_phv_out_data_443(mau_5_io_pipe_phv_out_data_443),
    .io_pipe_phv_out_data_444(mau_5_io_pipe_phv_out_data_444),
    .io_pipe_phv_out_data_445(mau_5_io_pipe_phv_out_data_445),
    .io_pipe_phv_out_data_446(mau_5_io_pipe_phv_out_data_446),
    .io_pipe_phv_out_data_447(mau_5_io_pipe_phv_out_data_447),
    .io_pipe_phv_out_data_448(mau_5_io_pipe_phv_out_data_448),
    .io_pipe_phv_out_data_449(mau_5_io_pipe_phv_out_data_449),
    .io_pipe_phv_out_data_450(mau_5_io_pipe_phv_out_data_450),
    .io_pipe_phv_out_data_451(mau_5_io_pipe_phv_out_data_451),
    .io_pipe_phv_out_data_452(mau_5_io_pipe_phv_out_data_452),
    .io_pipe_phv_out_data_453(mau_5_io_pipe_phv_out_data_453),
    .io_pipe_phv_out_data_454(mau_5_io_pipe_phv_out_data_454),
    .io_pipe_phv_out_data_455(mau_5_io_pipe_phv_out_data_455),
    .io_pipe_phv_out_data_456(mau_5_io_pipe_phv_out_data_456),
    .io_pipe_phv_out_data_457(mau_5_io_pipe_phv_out_data_457),
    .io_pipe_phv_out_data_458(mau_5_io_pipe_phv_out_data_458),
    .io_pipe_phv_out_data_459(mau_5_io_pipe_phv_out_data_459),
    .io_pipe_phv_out_data_460(mau_5_io_pipe_phv_out_data_460),
    .io_pipe_phv_out_data_461(mau_5_io_pipe_phv_out_data_461),
    .io_pipe_phv_out_data_462(mau_5_io_pipe_phv_out_data_462),
    .io_pipe_phv_out_data_463(mau_5_io_pipe_phv_out_data_463),
    .io_pipe_phv_out_data_464(mau_5_io_pipe_phv_out_data_464),
    .io_pipe_phv_out_data_465(mau_5_io_pipe_phv_out_data_465),
    .io_pipe_phv_out_data_466(mau_5_io_pipe_phv_out_data_466),
    .io_pipe_phv_out_data_467(mau_5_io_pipe_phv_out_data_467),
    .io_pipe_phv_out_data_468(mau_5_io_pipe_phv_out_data_468),
    .io_pipe_phv_out_data_469(mau_5_io_pipe_phv_out_data_469),
    .io_pipe_phv_out_data_470(mau_5_io_pipe_phv_out_data_470),
    .io_pipe_phv_out_data_471(mau_5_io_pipe_phv_out_data_471),
    .io_pipe_phv_out_data_472(mau_5_io_pipe_phv_out_data_472),
    .io_pipe_phv_out_data_473(mau_5_io_pipe_phv_out_data_473),
    .io_pipe_phv_out_data_474(mau_5_io_pipe_phv_out_data_474),
    .io_pipe_phv_out_data_475(mau_5_io_pipe_phv_out_data_475),
    .io_pipe_phv_out_data_476(mau_5_io_pipe_phv_out_data_476),
    .io_pipe_phv_out_data_477(mau_5_io_pipe_phv_out_data_477),
    .io_pipe_phv_out_data_478(mau_5_io_pipe_phv_out_data_478),
    .io_pipe_phv_out_data_479(mau_5_io_pipe_phv_out_data_479),
    .io_pipe_phv_out_data_480(mau_5_io_pipe_phv_out_data_480),
    .io_pipe_phv_out_data_481(mau_5_io_pipe_phv_out_data_481),
    .io_pipe_phv_out_data_482(mau_5_io_pipe_phv_out_data_482),
    .io_pipe_phv_out_data_483(mau_5_io_pipe_phv_out_data_483),
    .io_pipe_phv_out_data_484(mau_5_io_pipe_phv_out_data_484),
    .io_pipe_phv_out_data_485(mau_5_io_pipe_phv_out_data_485),
    .io_pipe_phv_out_data_486(mau_5_io_pipe_phv_out_data_486),
    .io_pipe_phv_out_data_487(mau_5_io_pipe_phv_out_data_487),
    .io_pipe_phv_out_data_488(mau_5_io_pipe_phv_out_data_488),
    .io_pipe_phv_out_data_489(mau_5_io_pipe_phv_out_data_489),
    .io_pipe_phv_out_data_490(mau_5_io_pipe_phv_out_data_490),
    .io_pipe_phv_out_data_491(mau_5_io_pipe_phv_out_data_491),
    .io_pipe_phv_out_data_492(mau_5_io_pipe_phv_out_data_492),
    .io_pipe_phv_out_data_493(mau_5_io_pipe_phv_out_data_493),
    .io_pipe_phv_out_data_494(mau_5_io_pipe_phv_out_data_494),
    .io_pipe_phv_out_data_495(mau_5_io_pipe_phv_out_data_495),
    .io_pipe_phv_out_data_496(mau_5_io_pipe_phv_out_data_496),
    .io_pipe_phv_out_data_497(mau_5_io_pipe_phv_out_data_497),
    .io_pipe_phv_out_data_498(mau_5_io_pipe_phv_out_data_498),
    .io_pipe_phv_out_data_499(mau_5_io_pipe_phv_out_data_499),
    .io_pipe_phv_out_data_500(mau_5_io_pipe_phv_out_data_500),
    .io_pipe_phv_out_data_501(mau_5_io_pipe_phv_out_data_501),
    .io_pipe_phv_out_data_502(mau_5_io_pipe_phv_out_data_502),
    .io_pipe_phv_out_data_503(mau_5_io_pipe_phv_out_data_503),
    .io_pipe_phv_out_data_504(mau_5_io_pipe_phv_out_data_504),
    .io_pipe_phv_out_data_505(mau_5_io_pipe_phv_out_data_505),
    .io_pipe_phv_out_data_506(mau_5_io_pipe_phv_out_data_506),
    .io_pipe_phv_out_data_507(mau_5_io_pipe_phv_out_data_507),
    .io_pipe_phv_out_data_508(mau_5_io_pipe_phv_out_data_508),
    .io_pipe_phv_out_data_509(mau_5_io_pipe_phv_out_data_509),
    .io_pipe_phv_out_data_510(mau_5_io_pipe_phv_out_data_510),
    .io_pipe_phv_out_data_511(mau_5_io_pipe_phv_out_data_511),
    .io_pipe_phv_out_header_0(mau_5_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(mau_5_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(mau_5_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(mau_5_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(mau_5_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(mau_5_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(mau_5_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(mau_5_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(mau_5_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(mau_5_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(mau_5_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(mau_5_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(mau_5_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(mau_5_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(mau_5_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(mau_5_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(mau_5_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(mau_5_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(mau_5_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(mau_5_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(mau_5_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(mau_5_io_pipe_phv_out_is_valid_processor),
    .io_mod_state_id_mod(mau_5_io_mod_state_id_mod),
    .io_mod_state_id(mau_5_io_mod_state_id),
    .io_mod_sram_w_cs(mau_5_io_mod_sram_w_cs),
    .io_mod_sram_w_en(mau_5_io_mod_sram_w_en),
    .io_mod_sram_w_addr(mau_5_io_mod_sram_w_addr),
    .io_mod_sram_w_data(mau_5_io_mod_sram_w_data)
  );
  ParseModule mau_6 ( // @[parser_pisa.scala 31:25]
    .clock(mau_6_clock),
    .io_pipe_phv_in_data_0(mau_6_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(mau_6_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(mau_6_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(mau_6_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(mau_6_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(mau_6_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(mau_6_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(mau_6_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(mau_6_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(mau_6_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(mau_6_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(mau_6_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(mau_6_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(mau_6_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(mau_6_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(mau_6_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(mau_6_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(mau_6_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(mau_6_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(mau_6_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(mau_6_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(mau_6_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(mau_6_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(mau_6_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(mau_6_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(mau_6_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(mau_6_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(mau_6_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(mau_6_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(mau_6_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(mau_6_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(mau_6_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(mau_6_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(mau_6_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(mau_6_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(mau_6_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(mau_6_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(mau_6_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(mau_6_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(mau_6_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(mau_6_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(mau_6_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(mau_6_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(mau_6_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(mau_6_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(mau_6_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(mau_6_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(mau_6_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(mau_6_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(mau_6_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(mau_6_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(mau_6_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(mau_6_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(mau_6_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(mau_6_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(mau_6_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(mau_6_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(mau_6_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(mau_6_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(mau_6_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(mau_6_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(mau_6_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(mau_6_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(mau_6_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(mau_6_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(mau_6_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(mau_6_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(mau_6_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(mau_6_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(mau_6_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(mau_6_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(mau_6_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(mau_6_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(mau_6_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(mau_6_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(mau_6_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(mau_6_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(mau_6_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(mau_6_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(mau_6_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(mau_6_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(mau_6_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(mau_6_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(mau_6_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(mau_6_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(mau_6_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(mau_6_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(mau_6_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(mau_6_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(mau_6_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(mau_6_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(mau_6_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(mau_6_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(mau_6_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(mau_6_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(mau_6_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(mau_6_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(mau_6_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(mau_6_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(mau_6_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(mau_6_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(mau_6_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(mau_6_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(mau_6_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(mau_6_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(mau_6_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(mau_6_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(mau_6_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(mau_6_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(mau_6_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(mau_6_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(mau_6_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(mau_6_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(mau_6_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(mau_6_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(mau_6_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(mau_6_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(mau_6_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(mau_6_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(mau_6_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(mau_6_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(mau_6_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(mau_6_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(mau_6_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(mau_6_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(mau_6_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(mau_6_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(mau_6_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(mau_6_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(mau_6_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(mau_6_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(mau_6_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(mau_6_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(mau_6_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(mau_6_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(mau_6_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(mau_6_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(mau_6_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(mau_6_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(mau_6_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(mau_6_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(mau_6_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(mau_6_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(mau_6_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(mau_6_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(mau_6_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(mau_6_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(mau_6_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(mau_6_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(mau_6_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(mau_6_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(mau_6_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(mau_6_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(mau_6_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(mau_6_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(mau_6_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(mau_6_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(mau_6_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(mau_6_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(mau_6_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(mau_6_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(mau_6_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(mau_6_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(mau_6_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(mau_6_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(mau_6_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(mau_6_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(mau_6_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(mau_6_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(mau_6_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(mau_6_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(mau_6_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(mau_6_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(mau_6_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(mau_6_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(mau_6_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(mau_6_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(mau_6_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(mau_6_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(mau_6_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(mau_6_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(mau_6_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(mau_6_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(mau_6_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(mau_6_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(mau_6_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(mau_6_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(mau_6_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(mau_6_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(mau_6_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(mau_6_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(mau_6_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(mau_6_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(mau_6_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(mau_6_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(mau_6_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(mau_6_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(mau_6_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(mau_6_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(mau_6_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(mau_6_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(mau_6_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(mau_6_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(mau_6_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(mau_6_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(mau_6_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(mau_6_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(mau_6_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(mau_6_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(mau_6_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(mau_6_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(mau_6_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(mau_6_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(mau_6_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(mau_6_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(mau_6_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(mau_6_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(mau_6_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(mau_6_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(mau_6_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(mau_6_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(mau_6_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(mau_6_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(mau_6_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(mau_6_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(mau_6_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(mau_6_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(mau_6_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(mau_6_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(mau_6_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(mau_6_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(mau_6_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(mau_6_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(mau_6_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(mau_6_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(mau_6_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(mau_6_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(mau_6_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(mau_6_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(mau_6_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(mau_6_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(mau_6_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(mau_6_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(mau_6_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(mau_6_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(mau_6_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(mau_6_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(mau_6_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(mau_6_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(mau_6_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(mau_6_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(mau_6_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(mau_6_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(mau_6_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(mau_6_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(mau_6_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_data_256(mau_6_io_pipe_phv_in_data_256),
    .io_pipe_phv_in_data_257(mau_6_io_pipe_phv_in_data_257),
    .io_pipe_phv_in_data_258(mau_6_io_pipe_phv_in_data_258),
    .io_pipe_phv_in_data_259(mau_6_io_pipe_phv_in_data_259),
    .io_pipe_phv_in_data_260(mau_6_io_pipe_phv_in_data_260),
    .io_pipe_phv_in_data_261(mau_6_io_pipe_phv_in_data_261),
    .io_pipe_phv_in_data_262(mau_6_io_pipe_phv_in_data_262),
    .io_pipe_phv_in_data_263(mau_6_io_pipe_phv_in_data_263),
    .io_pipe_phv_in_data_264(mau_6_io_pipe_phv_in_data_264),
    .io_pipe_phv_in_data_265(mau_6_io_pipe_phv_in_data_265),
    .io_pipe_phv_in_data_266(mau_6_io_pipe_phv_in_data_266),
    .io_pipe_phv_in_data_267(mau_6_io_pipe_phv_in_data_267),
    .io_pipe_phv_in_data_268(mau_6_io_pipe_phv_in_data_268),
    .io_pipe_phv_in_data_269(mau_6_io_pipe_phv_in_data_269),
    .io_pipe_phv_in_data_270(mau_6_io_pipe_phv_in_data_270),
    .io_pipe_phv_in_data_271(mau_6_io_pipe_phv_in_data_271),
    .io_pipe_phv_in_data_272(mau_6_io_pipe_phv_in_data_272),
    .io_pipe_phv_in_data_273(mau_6_io_pipe_phv_in_data_273),
    .io_pipe_phv_in_data_274(mau_6_io_pipe_phv_in_data_274),
    .io_pipe_phv_in_data_275(mau_6_io_pipe_phv_in_data_275),
    .io_pipe_phv_in_data_276(mau_6_io_pipe_phv_in_data_276),
    .io_pipe_phv_in_data_277(mau_6_io_pipe_phv_in_data_277),
    .io_pipe_phv_in_data_278(mau_6_io_pipe_phv_in_data_278),
    .io_pipe_phv_in_data_279(mau_6_io_pipe_phv_in_data_279),
    .io_pipe_phv_in_data_280(mau_6_io_pipe_phv_in_data_280),
    .io_pipe_phv_in_data_281(mau_6_io_pipe_phv_in_data_281),
    .io_pipe_phv_in_data_282(mau_6_io_pipe_phv_in_data_282),
    .io_pipe_phv_in_data_283(mau_6_io_pipe_phv_in_data_283),
    .io_pipe_phv_in_data_284(mau_6_io_pipe_phv_in_data_284),
    .io_pipe_phv_in_data_285(mau_6_io_pipe_phv_in_data_285),
    .io_pipe_phv_in_data_286(mau_6_io_pipe_phv_in_data_286),
    .io_pipe_phv_in_data_287(mau_6_io_pipe_phv_in_data_287),
    .io_pipe_phv_in_data_288(mau_6_io_pipe_phv_in_data_288),
    .io_pipe_phv_in_data_289(mau_6_io_pipe_phv_in_data_289),
    .io_pipe_phv_in_data_290(mau_6_io_pipe_phv_in_data_290),
    .io_pipe_phv_in_data_291(mau_6_io_pipe_phv_in_data_291),
    .io_pipe_phv_in_data_292(mau_6_io_pipe_phv_in_data_292),
    .io_pipe_phv_in_data_293(mau_6_io_pipe_phv_in_data_293),
    .io_pipe_phv_in_data_294(mau_6_io_pipe_phv_in_data_294),
    .io_pipe_phv_in_data_295(mau_6_io_pipe_phv_in_data_295),
    .io_pipe_phv_in_data_296(mau_6_io_pipe_phv_in_data_296),
    .io_pipe_phv_in_data_297(mau_6_io_pipe_phv_in_data_297),
    .io_pipe_phv_in_data_298(mau_6_io_pipe_phv_in_data_298),
    .io_pipe_phv_in_data_299(mau_6_io_pipe_phv_in_data_299),
    .io_pipe_phv_in_data_300(mau_6_io_pipe_phv_in_data_300),
    .io_pipe_phv_in_data_301(mau_6_io_pipe_phv_in_data_301),
    .io_pipe_phv_in_data_302(mau_6_io_pipe_phv_in_data_302),
    .io_pipe_phv_in_data_303(mau_6_io_pipe_phv_in_data_303),
    .io_pipe_phv_in_data_304(mau_6_io_pipe_phv_in_data_304),
    .io_pipe_phv_in_data_305(mau_6_io_pipe_phv_in_data_305),
    .io_pipe_phv_in_data_306(mau_6_io_pipe_phv_in_data_306),
    .io_pipe_phv_in_data_307(mau_6_io_pipe_phv_in_data_307),
    .io_pipe_phv_in_data_308(mau_6_io_pipe_phv_in_data_308),
    .io_pipe_phv_in_data_309(mau_6_io_pipe_phv_in_data_309),
    .io_pipe_phv_in_data_310(mau_6_io_pipe_phv_in_data_310),
    .io_pipe_phv_in_data_311(mau_6_io_pipe_phv_in_data_311),
    .io_pipe_phv_in_data_312(mau_6_io_pipe_phv_in_data_312),
    .io_pipe_phv_in_data_313(mau_6_io_pipe_phv_in_data_313),
    .io_pipe_phv_in_data_314(mau_6_io_pipe_phv_in_data_314),
    .io_pipe_phv_in_data_315(mau_6_io_pipe_phv_in_data_315),
    .io_pipe_phv_in_data_316(mau_6_io_pipe_phv_in_data_316),
    .io_pipe_phv_in_data_317(mau_6_io_pipe_phv_in_data_317),
    .io_pipe_phv_in_data_318(mau_6_io_pipe_phv_in_data_318),
    .io_pipe_phv_in_data_319(mau_6_io_pipe_phv_in_data_319),
    .io_pipe_phv_in_data_320(mau_6_io_pipe_phv_in_data_320),
    .io_pipe_phv_in_data_321(mau_6_io_pipe_phv_in_data_321),
    .io_pipe_phv_in_data_322(mau_6_io_pipe_phv_in_data_322),
    .io_pipe_phv_in_data_323(mau_6_io_pipe_phv_in_data_323),
    .io_pipe_phv_in_data_324(mau_6_io_pipe_phv_in_data_324),
    .io_pipe_phv_in_data_325(mau_6_io_pipe_phv_in_data_325),
    .io_pipe_phv_in_data_326(mau_6_io_pipe_phv_in_data_326),
    .io_pipe_phv_in_data_327(mau_6_io_pipe_phv_in_data_327),
    .io_pipe_phv_in_data_328(mau_6_io_pipe_phv_in_data_328),
    .io_pipe_phv_in_data_329(mau_6_io_pipe_phv_in_data_329),
    .io_pipe_phv_in_data_330(mau_6_io_pipe_phv_in_data_330),
    .io_pipe_phv_in_data_331(mau_6_io_pipe_phv_in_data_331),
    .io_pipe_phv_in_data_332(mau_6_io_pipe_phv_in_data_332),
    .io_pipe_phv_in_data_333(mau_6_io_pipe_phv_in_data_333),
    .io_pipe_phv_in_data_334(mau_6_io_pipe_phv_in_data_334),
    .io_pipe_phv_in_data_335(mau_6_io_pipe_phv_in_data_335),
    .io_pipe_phv_in_data_336(mau_6_io_pipe_phv_in_data_336),
    .io_pipe_phv_in_data_337(mau_6_io_pipe_phv_in_data_337),
    .io_pipe_phv_in_data_338(mau_6_io_pipe_phv_in_data_338),
    .io_pipe_phv_in_data_339(mau_6_io_pipe_phv_in_data_339),
    .io_pipe_phv_in_data_340(mau_6_io_pipe_phv_in_data_340),
    .io_pipe_phv_in_data_341(mau_6_io_pipe_phv_in_data_341),
    .io_pipe_phv_in_data_342(mau_6_io_pipe_phv_in_data_342),
    .io_pipe_phv_in_data_343(mau_6_io_pipe_phv_in_data_343),
    .io_pipe_phv_in_data_344(mau_6_io_pipe_phv_in_data_344),
    .io_pipe_phv_in_data_345(mau_6_io_pipe_phv_in_data_345),
    .io_pipe_phv_in_data_346(mau_6_io_pipe_phv_in_data_346),
    .io_pipe_phv_in_data_347(mau_6_io_pipe_phv_in_data_347),
    .io_pipe_phv_in_data_348(mau_6_io_pipe_phv_in_data_348),
    .io_pipe_phv_in_data_349(mau_6_io_pipe_phv_in_data_349),
    .io_pipe_phv_in_data_350(mau_6_io_pipe_phv_in_data_350),
    .io_pipe_phv_in_data_351(mau_6_io_pipe_phv_in_data_351),
    .io_pipe_phv_in_data_352(mau_6_io_pipe_phv_in_data_352),
    .io_pipe_phv_in_data_353(mau_6_io_pipe_phv_in_data_353),
    .io_pipe_phv_in_data_354(mau_6_io_pipe_phv_in_data_354),
    .io_pipe_phv_in_data_355(mau_6_io_pipe_phv_in_data_355),
    .io_pipe_phv_in_data_356(mau_6_io_pipe_phv_in_data_356),
    .io_pipe_phv_in_data_357(mau_6_io_pipe_phv_in_data_357),
    .io_pipe_phv_in_data_358(mau_6_io_pipe_phv_in_data_358),
    .io_pipe_phv_in_data_359(mau_6_io_pipe_phv_in_data_359),
    .io_pipe_phv_in_data_360(mau_6_io_pipe_phv_in_data_360),
    .io_pipe_phv_in_data_361(mau_6_io_pipe_phv_in_data_361),
    .io_pipe_phv_in_data_362(mau_6_io_pipe_phv_in_data_362),
    .io_pipe_phv_in_data_363(mau_6_io_pipe_phv_in_data_363),
    .io_pipe_phv_in_data_364(mau_6_io_pipe_phv_in_data_364),
    .io_pipe_phv_in_data_365(mau_6_io_pipe_phv_in_data_365),
    .io_pipe_phv_in_data_366(mau_6_io_pipe_phv_in_data_366),
    .io_pipe_phv_in_data_367(mau_6_io_pipe_phv_in_data_367),
    .io_pipe_phv_in_data_368(mau_6_io_pipe_phv_in_data_368),
    .io_pipe_phv_in_data_369(mau_6_io_pipe_phv_in_data_369),
    .io_pipe_phv_in_data_370(mau_6_io_pipe_phv_in_data_370),
    .io_pipe_phv_in_data_371(mau_6_io_pipe_phv_in_data_371),
    .io_pipe_phv_in_data_372(mau_6_io_pipe_phv_in_data_372),
    .io_pipe_phv_in_data_373(mau_6_io_pipe_phv_in_data_373),
    .io_pipe_phv_in_data_374(mau_6_io_pipe_phv_in_data_374),
    .io_pipe_phv_in_data_375(mau_6_io_pipe_phv_in_data_375),
    .io_pipe_phv_in_data_376(mau_6_io_pipe_phv_in_data_376),
    .io_pipe_phv_in_data_377(mau_6_io_pipe_phv_in_data_377),
    .io_pipe_phv_in_data_378(mau_6_io_pipe_phv_in_data_378),
    .io_pipe_phv_in_data_379(mau_6_io_pipe_phv_in_data_379),
    .io_pipe_phv_in_data_380(mau_6_io_pipe_phv_in_data_380),
    .io_pipe_phv_in_data_381(mau_6_io_pipe_phv_in_data_381),
    .io_pipe_phv_in_data_382(mau_6_io_pipe_phv_in_data_382),
    .io_pipe_phv_in_data_383(mau_6_io_pipe_phv_in_data_383),
    .io_pipe_phv_in_data_384(mau_6_io_pipe_phv_in_data_384),
    .io_pipe_phv_in_data_385(mau_6_io_pipe_phv_in_data_385),
    .io_pipe_phv_in_data_386(mau_6_io_pipe_phv_in_data_386),
    .io_pipe_phv_in_data_387(mau_6_io_pipe_phv_in_data_387),
    .io_pipe_phv_in_data_388(mau_6_io_pipe_phv_in_data_388),
    .io_pipe_phv_in_data_389(mau_6_io_pipe_phv_in_data_389),
    .io_pipe_phv_in_data_390(mau_6_io_pipe_phv_in_data_390),
    .io_pipe_phv_in_data_391(mau_6_io_pipe_phv_in_data_391),
    .io_pipe_phv_in_data_392(mau_6_io_pipe_phv_in_data_392),
    .io_pipe_phv_in_data_393(mau_6_io_pipe_phv_in_data_393),
    .io_pipe_phv_in_data_394(mau_6_io_pipe_phv_in_data_394),
    .io_pipe_phv_in_data_395(mau_6_io_pipe_phv_in_data_395),
    .io_pipe_phv_in_data_396(mau_6_io_pipe_phv_in_data_396),
    .io_pipe_phv_in_data_397(mau_6_io_pipe_phv_in_data_397),
    .io_pipe_phv_in_data_398(mau_6_io_pipe_phv_in_data_398),
    .io_pipe_phv_in_data_399(mau_6_io_pipe_phv_in_data_399),
    .io_pipe_phv_in_data_400(mau_6_io_pipe_phv_in_data_400),
    .io_pipe_phv_in_data_401(mau_6_io_pipe_phv_in_data_401),
    .io_pipe_phv_in_data_402(mau_6_io_pipe_phv_in_data_402),
    .io_pipe_phv_in_data_403(mau_6_io_pipe_phv_in_data_403),
    .io_pipe_phv_in_data_404(mau_6_io_pipe_phv_in_data_404),
    .io_pipe_phv_in_data_405(mau_6_io_pipe_phv_in_data_405),
    .io_pipe_phv_in_data_406(mau_6_io_pipe_phv_in_data_406),
    .io_pipe_phv_in_data_407(mau_6_io_pipe_phv_in_data_407),
    .io_pipe_phv_in_data_408(mau_6_io_pipe_phv_in_data_408),
    .io_pipe_phv_in_data_409(mau_6_io_pipe_phv_in_data_409),
    .io_pipe_phv_in_data_410(mau_6_io_pipe_phv_in_data_410),
    .io_pipe_phv_in_data_411(mau_6_io_pipe_phv_in_data_411),
    .io_pipe_phv_in_data_412(mau_6_io_pipe_phv_in_data_412),
    .io_pipe_phv_in_data_413(mau_6_io_pipe_phv_in_data_413),
    .io_pipe_phv_in_data_414(mau_6_io_pipe_phv_in_data_414),
    .io_pipe_phv_in_data_415(mau_6_io_pipe_phv_in_data_415),
    .io_pipe_phv_in_data_416(mau_6_io_pipe_phv_in_data_416),
    .io_pipe_phv_in_data_417(mau_6_io_pipe_phv_in_data_417),
    .io_pipe_phv_in_data_418(mau_6_io_pipe_phv_in_data_418),
    .io_pipe_phv_in_data_419(mau_6_io_pipe_phv_in_data_419),
    .io_pipe_phv_in_data_420(mau_6_io_pipe_phv_in_data_420),
    .io_pipe_phv_in_data_421(mau_6_io_pipe_phv_in_data_421),
    .io_pipe_phv_in_data_422(mau_6_io_pipe_phv_in_data_422),
    .io_pipe_phv_in_data_423(mau_6_io_pipe_phv_in_data_423),
    .io_pipe_phv_in_data_424(mau_6_io_pipe_phv_in_data_424),
    .io_pipe_phv_in_data_425(mau_6_io_pipe_phv_in_data_425),
    .io_pipe_phv_in_data_426(mau_6_io_pipe_phv_in_data_426),
    .io_pipe_phv_in_data_427(mau_6_io_pipe_phv_in_data_427),
    .io_pipe_phv_in_data_428(mau_6_io_pipe_phv_in_data_428),
    .io_pipe_phv_in_data_429(mau_6_io_pipe_phv_in_data_429),
    .io_pipe_phv_in_data_430(mau_6_io_pipe_phv_in_data_430),
    .io_pipe_phv_in_data_431(mau_6_io_pipe_phv_in_data_431),
    .io_pipe_phv_in_data_432(mau_6_io_pipe_phv_in_data_432),
    .io_pipe_phv_in_data_433(mau_6_io_pipe_phv_in_data_433),
    .io_pipe_phv_in_data_434(mau_6_io_pipe_phv_in_data_434),
    .io_pipe_phv_in_data_435(mau_6_io_pipe_phv_in_data_435),
    .io_pipe_phv_in_data_436(mau_6_io_pipe_phv_in_data_436),
    .io_pipe_phv_in_data_437(mau_6_io_pipe_phv_in_data_437),
    .io_pipe_phv_in_data_438(mau_6_io_pipe_phv_in_data_438),
    .io_pipe_phv_in_data_439(mau_6_io_pipe_phv_in_data_439),
    .io_pipe_phv_in_data_440(mau_6_io_pipe_phv_in_data_440),
    .io_pipe_phv_in_data_441(mau_6_io_pipe_phv_in_data_441),
    .io_pipe_phv_in_data_442(mau_6_io_pipe_phv_in_data_442),
    .io_pipe_phv_in_data_443(mau_6_io_pipe_phv_in_data_443),
    .io_pipe_phv_in_data_444(mau_6_io_pipe_phv_in_data_444),
    .io_pipe_phv_in_data_445(mau_6_io_pipe_phv_in_data_445),
    .io_pipe_phv_in_data_446(mau_6_io_pipe_phv_in_data_446),
    .io_pipe_phv_in_data_447(mau_6_io_pipe_phv_in_data_447),
    .io_pipe_phv_in_data_448(mau_6_io_pipe_phv_in_data_448),
    .io_pipe_phv_in_data_449(mau_6_io_pipe_phv_in_data_449),
    .io_pipe_phv_in_data_450(mau_6_io_pipe_phv_in_data_450),
    .io_pipe_phv_in_data_451(mau_6_io_pipe_phv_in_data_451),
    .io_pipe_phv_in_data_452(mau_6_io_pipe_phv_in_data_452),
    .io_pipe_phv_in_data_453(mau_6_io_pipe_phv_in_data_453),
    .io_pipe_phv_in_data_454(mau_6_io_pipe_phv_in_data_454),
    .io_pipe_phv_in_data_455(mau_6_io_pipe_phv_in_data_455),
    .io_pipe_phv_in_data_456(mau_6_io_pipe_phv_in_data_456),
    .io_pipe_phv_in_data_457(mau_6_io_pipe_phv_in_data_457),
    .io_pipe_phv_in_data_458(mau_6_io_pipe_phv_in_data_458),
    .io_pipe_phv_in_data_459(mau_6_io_pipe_phv_in_data_459),
    .io_pipe_phv_in_data_460(mau_6_io_pipe_phv_in_data_460),
    .io_pipe_phv_in_data_461(mau_6_io_pipe_phv_in_data_461),
    .io_pipe_phv_in_data_462(mau_6_io_pipe_phv_in_data_462),
    .io_pipe_phv_in_data_463(mau_6_io_pipe_phv_in_data_463),
    .io_pipe_phv_in_data_464(mau_6_io_pipe_phv_in_data_464),
    .io_pipe_phv_in_data_465(mau_6_io_pipe_phv_in_data_465),
    .io_pipe_phv_in_data_466(mau_6_io_pipe_phv_in_data_466),
    .io_pipe_phv_in_data_467(mau_6_io_pipe_phv_in_data_467),
    .io_pipe_phv_in_data_468(mau_6_io_pipe_phv_in_data_468),
    .io_pipe_phv_in_data_469(mau_6_io_pipe_phv_in_data_469),
    .io_pipe_phv_in_data_470(mau_6_io_pipe_phv_in_data_470),
    .io_pipe_phv_in_data_471(mau_6_io_pipe_phv_in_data_471),
    .io_pipe_phv_in_data_472(mau_6_io_pipe_phv_in_data_472),
    .io_pipe_phv_in_data_473(mau_6_io_pipe_phv_in_data_473),
    .io_pipe_phv_in_data_474(mau_6_io_pipe_phv_in_data_474),
    .io_pipe_phv_in_data_475(mau_6_io_pipe_phv_in_data_475),
    .io_pipe_phv_in_data_476(mau_6_io_pipe_phv_in_data_476),
    .io_pipe_phv_in_data_477(mau_6_io_pipe_phv_in_data_477),
    .io_pipe_phv_in_data_478(mau_6_io_pipe_phv_in_data_478),
    .io_pipe_phv_in_data_479(mau_6_io_pipe_phv_in_data_479),
    .io_pipe_phv_in_data_480(mau_6_io_pipe_phv_in_data_480),
    .io_pipe_phv_in_data_481(mau_6_io_pipe_phv_in_data_481),
    .io_pipe_phv_in_data_482(mau_6_io_pipe_phv_in_data_482),
    .io_pipe_phv_in_data_483(mau_6_io_pipe_phv_in_data_483),
    .io_pipe_phv_in_data_484(mau_6_io_pipe_phv_in_data_484),
    .io_pipe_phv_in_data_485(mau_6_io_pipe_phv_in_data_485),
    .io_pipe_phv_in_data_486(mau_6_io_pipe_phv_in_data_486),
    .io_pipe_phv_in_data_487(mau_6_io_pipe_phv_in_data_487),
    .io_pipe_phv_in_data_488(mau_6_io_pipe_phv_in_data_488),
    .io_pipe_phv_in_data_489(mau_6_io_pipe_phv_in_data_489),
    .io_pipe_phv_in_data_490(mau_6_io_pipe_phv_in_data_490),
    .io_pipe_phv_in_data_491(mau_6_io_pipe_phv_in_data_491),
    .io_pipe_phv_in_data_492(mau_6_io_pipe_phv_in_data_492),
    .io_pipe_phv_in_data_493(mau_6_io_pipe_phv_in_data_493),
    .io_pipe_phv_in_data_494(mau_6_io_pipe_phv_in_data_494),
    .io_pipe_phv_in_data_495(mau_6_io_pipe_phv_in_data_495),
    .io_pipe_phv_in_data_496(mau_6_io_pipe_phv_in_data_496),
    .io_pipe_phv_in_data_497(mau_6_io_pipe_phv_in_data_497),
    .io_pipe_phv_in_data_498(mau_6_io_pipe_phv_in_data_498),
    .io_pipe_phv_in_data_499(mau_6_io_pipe_phv_in_data_499),
    .io_pipe_phv_in_data_500(mau_6_io_pipe_phv_in_data_500),
    .io_pipe_phv_in_data_501(mau_6_io_pipe_phv_in_data_501),
    .io_pipe_phv_in_data_502(mau_6_io_pipe_phv_in_data_502),
    .io_pipe_phv_in_data_503(mau_6_io_pipe_phv_in_data_503),
    .io_pipe_phv_in_data_504(mau_6_io_pipe_phv_in_data_504),
    .io_pipe_phv_in_data_505(mau_6_io_pipe_phv_in_data_505),
    .io_pipe_phv_in_data_506(mau_6_io_pipe_phv_in_data_506),
    .io_pipe_phv_in_data_507(mau_6_io_pipe_phv_in_data_507),
    .io_pipe_phv_in_data_508(mau_6_io_pipe_phv_in_data_508),
    .io_pipe_phv_in_data_509(mau_6_io_pipe_phv_in_data_509),
    .io_pipe_phv_in_data_510(mau_6_io_pipe_phv_in_data_510),
    .io_pipe_phv_in_data_511(mau_6_io_pipe_phv_in_data_511),
    .io_pipe_phv_in_header_0(mau_6_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(mau_6_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(mau_6_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(mau_6_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(mau_6_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(mau_6_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(mau_6_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(mau_6_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(mau_6_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(mau_6_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(mau_6_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(mau_6_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(mau_6_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(mau_6_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(mau_6_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(mau_6_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(mau_6_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(mau_6_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(mau_6_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(mau_6_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(mau_6_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(mau_6_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(mau_6_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(mau_6_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(mau_6_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(mau_6_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(mau_6_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(mau_6_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(mau_6_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(mau_6_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(mau_6_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(mau_6_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(mau_6_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(mau_6_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(mau_6_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(mau_6_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(mau_6_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(mau_6_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(mau_6_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(mau_6_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(mau_6_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(mau_6_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(mau_6_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(mau_6_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(mau_6_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(mau_6_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(mau_6_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(mau_6_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(mau_6_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(mau_6_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(mau_6_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(mau_6_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(mau_6_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(mau_6_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(mau_6_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(mau_6_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(mau_6_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(mau_6_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(mau_6_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(mau_6_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(mau_6_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(mau_6_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(mau_6_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(mau_6_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(mau_6_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(mau_6_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(mau_6_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(mau_6_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(mau_6_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(mau_6_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(mau_6_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(mau_6_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(mau_6_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(mau_6_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(mau_6_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(mau_6_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(mau_6_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(mau_6_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(mau_6_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(mau_6_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(mau_6_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(mau_6_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(mau_6_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(mau_6_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(mau_6_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(mau_6_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(mau_6_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(mau_6_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(mau_6_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(mau_6_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(mau_6_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(mau_6_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(mau_6_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(mau_6_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(mau_6_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(mau_6_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(mau_6_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(mau_6_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(mau_6_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(mau_6_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(mau_6_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(mau_6_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(mau_6_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(mau_6_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(mau_6_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(mau_6_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(mau_6_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(mau_6_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(mau_6_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(mau_6_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(mau_6_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(mau_6_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(mau_6_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(mau_6_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(mau_6_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(mau_6_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(mau_6_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(mau_6_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(mau_6_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(mau_6_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(mau_6_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(mau_6_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(mau_6_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(mau_6_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(mau_6_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(mau_6_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(mau_6_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(mau_6_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(mau_6_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(mau_6_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(mau_6_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(mau_6_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(mau_6_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(mau_6_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(mau_6_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(mau_6_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(mau_6_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(mau_6_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(mau_6_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(mau_6_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(mau_6_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(mau_6_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(mau_6_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(mau_6_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(mau_6_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(mau_6_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(mau_6_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(mau_6_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(mau_6_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(mau_6_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(mau_6_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(mau_6_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(mau_6_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(mau_6_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(mau_6_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(mau_6_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(mau_6_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(mau_6_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(mau_6_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(mau_6_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(mau_6_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(mau_6_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(mau_6_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(mau_6_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(mau_6_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(mau_6_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(mau_6_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(mau_6_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(mau_6_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(mau_6_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(mau_6_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(mau_6_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(mau_6_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(mau_6_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(mau_6_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(mau_6_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(mau_6_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(mau_6_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(mau_6_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(mau_6_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(mau_6_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(mau_6_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(mau_6_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(mau_6_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(mau_6_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(mau_6_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(mau_6_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(mau_6_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(mau_6_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(mau_6_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(mau_6_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(mau_6_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(mau_6_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(mau_6_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(mau_6_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(mau_6_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(mau_6_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(mau_6_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(mau_6_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(mau_6_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(mau_6_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(mau_6_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(mau_6_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(mau_6_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(mau_6_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(mau_6_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(mau_6_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(mau_6_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(mau_6_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(mau_6_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(mau_6_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(mau_6_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(mau_6_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(mau_6_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(mau_6_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(mau_6_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(mau_6_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(mau_6_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(mau_6_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(mau_6_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(mau_6_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(mau_6_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(mau_6_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(mau_6_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(mau_6_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(mau_6_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(mau_6_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(mau_6_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(mau_6_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(mau_6_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(mau_6_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(mau_6_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(mau_6_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(mau_6_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(mau_6_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(mau_6_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(mau_6_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(mau_6_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(mau_6_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(mau_6_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(mau_6_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(mau_6_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(mau_6_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(mau_6_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(mau_6_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(mau_6_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(mau_6_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(mau_6_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(mau_6_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(mau_6_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(mau_6_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(mau_6_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(mau_6_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(mau_6_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(mau_6_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(mau_6_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(mau_6_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(mau_6_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(mau_6_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(mau_6_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(mau_6_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(mau_6_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(mau_6_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(mau_6_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(mau_6_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(mau_6_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(mau_6_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(mau_6_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(mau_6_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(mau_6_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(mau_6_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(mau_6_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(mau_6_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(mau_6_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(mau_6_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(mau_6_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(mau_6_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(mau_6_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_data_256(mau_6_io_pipe_phv_out_data_256),
    .io_pipe_phv_out_data_257(mau_6_io_pipe_phv_out_data_257),
    .io_pipe_phv_out_data_258(mau_6_io_pipe_phv_out_data_258),
    .io_pipe_phv_out_data_259(mau_6_io_pipe_phv_out_data_259),
    .io_pipe_phv_out_data_260(mau_6_io_pipe_phv_out_data_260),
    .io_pipe_phv_out_data_261(mau_6_io_pipe_phv_out_data_261),
    .io_pipe_phv_out_data_262(mau_6_io_pipe_phv_out_data_262),
    .io_pipe_phv_out_data_263(mau_6_io_pipe_phv_out_data_263),
    .io_pipe_phv_out_data_264(mau_6_io_pipe_phv_out_data_264),
    .io_pipe_phv_out_data_265(mau_6_io_pipe_phv_out_data_265),
    .io_pipe_phv_out_data_266(mau_6_io_pipe_phv_out_data_266),
    .io_pipe_phv_out_data_267(mau_6_io_pipe_phv_out_data_267),
    .io_pipe_phv_out_data_268(mau_6_io_pipe_phv_out_data_268),
    .io_pipe_phv_out_data_269(mau_6_io_pipe_phv_out_data_269),
    .io_pipe_phv_out_data_270(mau_6_io_pipe_phv_out_data_270),
    .io_pipe_phv_out_data_271(mau_6_io_pipe_phv_out_data_271),
    .io_pipe_phv_out_data_272(mau_6_io_pipe_phv_out_data_272),
    .io_pipe_phv_out_data_273(mau_6_io_pipe_phv_out_data_273),
    .io_pipe_phv_out_data_274(mau_6_io_pipe_phv_out_data_274),
    .io_pipe_phv_out_data_275(mau_6_io_pipe_phv_out_data_275),
    .io_pipe_phv_out_data_276(mau_6_io_pipe_phv_out_data_276),
    .io_pipe_phv_out_data_277(mau_6_io_pipe_phv_out_data_277),
    .io_pipe_phv_out_data_278(mau_6_io_pipe_phv_out_data_278),
    .io_pipe_phv_out_data_279(mau_6_io_pipe_phv_out_data_279),
    .io_pipe_phv_out_data_280(mau_6_io_pipe_phv_out_data_280),
    .io_pipe_phv_out_data_281(mau_6_io_pipe_phv_out_data_281),
    .io_pipe_phv_out_data_282(mau_6_io_pipe_phv_out_data_282),
    .io_pipe_phv_out_data_283(mau_6_io_pipe_phv_out_data_283),
    .io_pipe_phv_out_data_284(mau_6_io_pipe_phv_out_data_284),
    .io_pipe_phv_out_data_285(mau_6_io_pipe_phv_out_data_285),
    .io_pipe_phv_out_data_286(mau_6_io_pipe_phv_out_data_286),
    .io_pipe_phv_out_data_287(mau_6_io_pipe_phv_out_data_287),
    .io_pipe_phv_out_data_288(mau_6_io_pipe_phv_out_data_288),
    .io_pipe_phv_out_data_289(mau_6_io_pipe_phv_out_data_289),
    .io_pipe_phv_out_data_290(mau_6_io_pipe_phv_out_data_290),
    .io_pipe_phv_out_data_291(mau_6_io_pipe_phv_out_data_291),
    .io_pipe_phv_out_data_292(mau_6_io_pipe_phv_out_data_292),
    .io_pipe_phv_out_data_293(mau_6_io_pipe_phv_out_data_293),
    .io_pipe_phv_out_data_294(mau_6_io_pipe_phv_out_data_294),
    .io_pipe_phv_out_data_295(mau_6_io_pipe_phv_out_data_295),
    .io_pipe_phv_out_data_296(mau_6_io_pipe_phv_out_data_296),
    .io_pipe_phv_out_data_297(mau_6_io_pipe_phv_out_data_297),
    .io_pipe_phv_out_data_298(mau_6_io_pipe_phv_out_data_298),
    .io_pipe_phv_out_data_299(mau_6_io_pipe_phv_out_data_299),
    .io_pipe_phv_out_data_300(mau_6_io_pipe_phv_out_data_300),
    .io_pipe_phv_out_data_301(mau_6_io_pipe_phv_out_data_301),
    .io_pipe_phv_out_data_302(mau_6_io_pipe_phv_out_data_302),
    .io_pipe_phv_out_data_303(mau_6_io_pipe_phv_out_data_303),
    .io_pipe_phv_out_data_304(mau_6_io_pipe_phv_out_data_304),
    .io_pipe_phv_out_data_305(mau_6_io_pipe_phv_out_data_305),
    .io_pipe_phv_out_data_306(mau_6_io_pipe_phv_out_data_306),
    .io_pipe_phv_out_data_307(mau_6_io_pipe_phv_out_data_307),
    .io_pipe_phv_out_data_308(mau_6_io_pipe_phv_out_data_308),
    .io_pipe_phv_out_data_309(mau_6_io_pipe_phv_out_data_309),
    .io_pipe_phv_out_data_310(mau_6_io_pipe_phv_out_data_310),
    .io_pipe_phv_out_data_311(mau_6_io_pipe_phv_out_data_311),
    .io_pipe_phv_out_data_312(mau_6_io_pipe_phv_out_data_312),
    .io_pipe_phv_out_data_313(mau_6_io_pipe_phv_out_data_313),
    .io_pipe_phv_out_data_314(mau_6_io_pipe_phv_out_data_314),
    .io_pipe_phv_out_data_315(mau_6_io_pipe_phv_out_data_315),
    .io_pipe_phv_out_data_316(mau_6_io_pipe_phv_out_data_316),
    .io_pipe_phv_out_data_317(mau_6_io_pipe_phv_out_data_317),
    .io_pipe_phv_out_data_318(mau_6_io_pipe_phv_out_data_318),
    .io_pipe_phv_out_data_319(mau_6_io_pipe_phv_out_data_319),
    .io_pipe_phv_out_data_320(mau_6_io_pipe_phv_out_data_320),
    .io_pipe_phv_out_data_321(mau_6_io_pipe_phv_out_data_321),
    .io_pipe_phv_out_data_322(mau_6_io_pipe_phv_out_data_322),
    .io_pipe_phv_out_data_323(mau_6_io_pipe_phv_out_data_323),
    .io_pipe_phv_out_data_324(mau_6_io_pipe_phv_out_data_324),
    .io_pipe_phv_out_data_325(mau_6_io_pipe_phv_out_data_325),
    .io_pipe_phv_out_data_326(mau_6_io_pipe_phv_out_data_326),
    .io_pipe_phv_out_data_327(mau_6_io_pipe_phv_out_data_327),
    .io_pipe_phv_out_data_328(mau_6_io_pipe_phv_out_data_328),
    .io_pipe_phv_out_data_329(mau_6_io_pipe_phv_out_data_329),
    .io_pipe_phv_out_data_330(mau_6_io_pipe_phv_out_data_330),
    .io_pipe_phv_out_data_331(mau_6_io_pipe_phv_out_data_331),
    .io_pipe_phv_out_data_332(mau_6_io_pipe_phv_out_data_332),
    .io_pipe_phv_out_data_333(mau_6_io_pipe_phv_out_data_333),
    .io_pipe_phv_out_data_334(mau_6_io_pipe_phv_out_data_334),
    .io_pipe_phv_out_data_335(mau_6_io_pipe_phv_out_data_335),
    .io_pipe_phv_out_data_336(mau_6_io_pipe_phv_out_data_336),
    .io_pipe_phv_out_data_337(mau_6_io_pipe_phv_out_data_337),
    .io_pipe_phv_out_data_338(mau_6_io_pipe_phv_out_data_338),
    .io_pipe_phv_out_data_339(mau_6_io_pipe_phv_out_data_339),
    .io_pipe_phv_out_data_340(mau_6_io_pipe_phv_out_data_340),
    .io_pipe_phv_out_data_341(mau_6_io_pipe_phv_out_data_341),
    .io_pipe_phv_out_data_342(mau_6_io_pipe_phv_out_data_342),
    .io_pipe_phv_out_data_343(mau_6_io_pipe_phv_out_data_343),
    .io_pipe_phv_out_data_344(mau_6_io_pipe_phv_out_data_344),
    .io_pipe_phv_out_data_345(mau_6_io_pipe_phv_out_data_345),
    .io_pipe_phv_out_data_346(mau_6_io_pipe_phv_out_data_346),
    .io_pipe_phv_out_data_347(mau_6_io_pipe_phv_out_data_347),
    .io_pipe_phv_out_data_348(mau_6_io_pipe_phv_out_data_348),
    .io_pipe_phv_out_data_349(mau_6_io_pipe_phv_out_data_349),
    .io_pipe_phv_out_data_350(mau_6_io_pipe_phv_out_data_350),
    .io_pipe_phv_out_data_351(mau_6_io_pipe_phv_out_data_351),
    .io_pipe_phv_out_data_352(mau_6_io_pipe_phv_out_data_352),
    .io_pipe_phv_out_data_353(mau_6_io_pipe_phv_out_data_353),
    .io_pipe_phv_out_data_354(mau_6_io_pipe_phv_out_data_354),
    .io_pipe_phv_out_data_355(mau_6_io_pipe_phv_out_data_355),
    .io_pipe_phv_out_data_356(mau_6_io_pipe_phv_out_data_356),
    .io_pipe_phv_out_data_357(mau_6_io_pipe_phv_out_data_357),
    .io_pipe_phv_out_data_358(mau_6_io_pipe_phv_out_data_358),
    .io_pipe_phv_out_data_359(mau_6_io_pipe_phv_out_data_359),
    .io_pipe_phv_out_data_360(mau_6_io_pipe_phv_out_data_360),
    .io_pipe_phv_out_data_361(mau_6_io_pipe_phv_out_data_361),
    .io_pipe_phv_out_data_362(mau_6_io_pipe_phv_out_data_362),
    .io_pipe_phv_out_data_363(mau_6_io_pipe_phv_out_data_363),
    .io_pipe_phv_out_data_364(mau_6_io_pipe_phv_out_data_364),
    .io_pipe_phv_out_data_365(mau_6_io_pipe_phv_out_data_365),
    .io_pipe_phv_out_data_366(mau_6_io_pipe_phv_out_data_366),
    .io_pipe_phv_out_data_367(mau_6_io_pipe_phv_out_data_367),
    .io_pipe_phv_out_data_368(mau_6_io_pipe_phv_out_data_368),
    .io_pipe_phv_out_data_369(mau_6_io_pipe_phv_out_data_369),
    .io_pipe_phv_out_data_370(mau_6_io_pipe_phv_out_data_370),
    .io_pipe_phv_out_data_371(mau_6_io_pipe_phv_out_data_371),
    .io_pipe_phv_out_data_372(mau_6_io_pipe_phv_out_data_372),
    .io_pipe_phv_out_data_373(mau_6_io_pipe_phv_out_data_373),
    .io_pipe_phv_out_data_374(mau_6_io_pipe_phv_out_data_374),
    .io_pipe_phv_out_data_375(mau_6_io_pipe_phv_out_data_375),
    .io_pipe_phv_out_data_376(mau_6_io_pipe_phv_out_data_376),
    .io_pipe_phv_out_data_377(mau_6_io_pipe_phv_out_data_377),
    .io_pipe_phv_out_data_378(mau_6_io_pipe_phv_out_data_378),
    .io_pipe_phv_out_data_379(mau_6_io_pipe_phv_out_data_379),
    .io_pipe_phv_out_data_380(mau_6_io_pipe_phv_out_data_380),
    .io_pipe_phv_out_data_381(mau_6_io_pipe_phv_out_data_381),
    .io_pipe_phv_out_data_382(mau_6_io_pipe_phv_out_data_382),
    .io_pipe_phv_out_data_383(mau_6_io_pipe_phv_out_data_383),
    .io_pipe_phv_out_data_384(mau_6_io_pipe_phv_out_data_384),
    .io_pipe_phv_out_data_385(mau_6_io_pipe_phv_out_data_385),
    .io_pipe_phv_out_data_386(mau_6_io_pipe_phv_out_data_386),
    .io_pipe_phv_out_data_387(mau_6_io_pipe_phv_out_data_387),
    .io_pipe_phv_out_data_388(mau_6_io_pipe_phv_out_data_388),
    .io_pipe_phv_out_data_389(mau_6_io_pipe_phv_out_data_389),
    .io_pipe_phv_out_data_390(mau_6_io_pipe_phv_out_data_390),
    .io_pipe_phv_out_data_391(mau_6_io_pipe_phv_out_data_391),
    .io_pipe_phv_out_data_392(mau_6_io_pipe_phv_out_data_392),
    .io_pipe_phv_out_data_393(mau_6_io_pipe_phv_out_data_393),
    .io_pipe_phv_out_data_394(mau_6_io_pipe_phv_out_data_394),
    .io_pipe_phv_out_data_395(mau_6_io_pipe_phv_out_data_395),
    .io_pipe_phv_out_data_396(mau_6_io_pipe_phv_out_data_396),
    .io_pipe_phv_out_data_397(mau_6_io_pipe_phv_out_data_397),
    .io_pipe_phv_out_data_398(mau_6_io_pipe_phv_out_data_398),
    .io_pipe_phv_out_data_399(mau_6_io_pipe_phv_out_data_399),
    .io_pipe_phv_out_data_400(mau_6_io_pipe_phv_out_data_400),
    .io_pipe_phv_out_data_401(mau_6_io_pipe_phv_out_data_401),
    .io_pipe_phv_out_data_402(mau_6_io_pipe_phv_out_data_402),
    .io_pipe_phv_out_data_403(mau_6_io_pipe_phv_out_data_403),
    .io_pipe_phv_out_data_404(mau_6_io_pipe_phv_out_data_404),
    .io_pipe_phv_out_data_405(mau_6_io_pipe_phv_out_data_405),
    .io_pipe_phv_out_data_406(mau_6_io_pipe_phv_out_data_406),
    .io_pipe_phv_out_data_407(mau_6_io_pipe_phv_out_data_407),
    .io_pipe_phv_out_data_408(mau_6_io_pipe_phv_out_data_408),
    .io_pipe_phv_out_data_409(mau_6_io_pipe_phv_out_data_409),
    .io_pipe_phv_out_data_410(mau_6_io_pipe_phv_out_data_410),
    .io_pipe_phv_out_data_411(mau_6_io_pipe_phv_out_data_411),
    .io_pipe_phv_out_data_412(mau_6_io_pipe_phv_out_data_412),
    .io_pipe_phv_out_data_413(mau_6_io_pipe_phv_out_data_413),
    .io_pipe_phv_out_data_414(mau_6_io_pipe_phv_out_data_414),
    .io_pipe_phv_out_data_415(mau_6_io_pipe_phv_out_data_415),
    .io_pipe_phv_out_data_416(mau_6_io_pipe_phv_out_data_416),
    .io_pipe_phv_out_data_417(mau_6_io_pipe_phv_out_data_417),
    .io_pipe_phv_out_data_418(mau_6_io_pipe_phv_out_data_418),
    .io_pipe_phv_out_data_419(mau_6_io_pipe_phv_out_data_419),
    .io_pipe_phv_out_data_420(mau_6_io_pipe_phv_out_data_420),
    .io_pipe_phv_out_data_421(mau_6_io_pipe_phv_out_data_421),
    .io_pipe_phv_out_data_422(mau_6_io_pipe_phv_out_data_422),
    .io_pipe_phv_out_data_423(mau_6_io_pipe_phv_out_data_423),
    .io_pipe_phv_out_data_424(mau_6_io_pipe_phv_out_data_424),
    .io_pipe_phv_out_data_425(mau_6_io_pipe_phv_out_data_425),
    .io_pipe_phv_out_data_426(mau_6_io_pipe_phv_out_data_426),
    .io_pipe_phv_out_data_427(mau_6_io_pipe_phv_out_data_427),
    .io_pipe_phv_out_data_428(mau_6_io_pipe_phv_out_data_428),
    .io_pipe_phv_out_data_429(mau_6_io_pipe_phv_out_data_429),
    .io_pipe_phv_out_data_430(mau_6_io_pipe_phv_out_data_430),
    .io_pipe_phv_out_data_431(mau_6_io_pipe_phv_out_data_431),
    .io_pipe_phv_out_data_432(mau_6_io_pipe_phv_out_data_432),
    .io_pipe_phv_out_data_433(mau_6_io_pipe_phv_out_data_433),
    .io_pipe_phv_out_data_434(mau_6_io_pipe_phv_out_data_434),
    .io_pipe_phv_out_data_435(mau_6_io_pipe_phv_out_data_435),
    .io_pipe_phv_out_data_436(mau_6_io_pipe_phv_out_data_436),
    .io_pipe_phv_out_data_437(mau_6_io_pipe_phv_out_data_437),
    .io_pipe_phv_out_data_438(mau_6_io_pipe_phv_out_data_438),
    .io_pipe_phv_out_data_439(mau_6_io_pipe_phv_out_data_439),
    .io_pipe_phv_out_data_440(mau_6_io_pipe_phv_out_data_440),
    .io_pipe_phv_out_data_441(mau_6_io_pipe_phv_out_data_441),
    .io_pipe_phv_out_data_442(mau_6_io_pipe_phv_out_data_442),
    .io_pipe_phv_out_data_443(mau_6_io_pipe_phv_out_data_443),
    .io_pipe_phv_out_data_444(mau_6_io_pipe_phv_out_data_444),
    .io_pipe_phv_out_data_445(mau_6_io_pipe_phv_out_data_445),
    .io_pipe_phv_out_data_446(mau_6_io_pipe_phv_out_data_446),
    .io_pipe_phv_out_data_447(mau_6_io_pipe_phv_out_data_447),
    .io_pipe_phv_out_data_448(mau_6_io_pipe_phv_out_data_448),
    .io_pipe_phv_out_data_449(mau_6_io_pipe_phv_out_data_449),
    .io_pipe_phv_out_data_450(mau_6_io_pipe_phv_out_data_450),
    .io_pipe_phv_out_data_451(mau_6_io_pipe_phv_out_data_451),
    .io_pipe_phv_out_data_452(mau_6_io_pipe_phv_out_data_452),
    .io_pipe_phv_out_data_453(mau_6_io_pipe_phv_out_data_453),
    .io_pipe_phv_out_data_454(mau_6_io_pipe_phv_out_data_454),
    .io_pipe_phv_out_data_455(mau_6_io_pipe_phv_out_data_455),
    .io_pipe_phv_out_data_456(mau_6_io_pipe_phv_out_data_456),
    .io_pipe_phv_out_data_457(mau_6_io_pipe_phv_out_data_457),
    .io_pipe_phv_out_data_458(mau_6_io_pipe_phv_out_data_458),
    .io_pipe_phv_out_data_459(mau_6_io_pipe_phv_out_data_459),
    .io_pipe_phv_out_data_460(mau_6_io_pipe_phv_out_data_460),
    .io_pipe_phv_out_data_461(mau_6_io_pipe_phv_out_data_461),
    .io_pipe_phv_out_data_462(mau_6_io_pipe_phv_out_data_462),
    .io_pipe_phv_out_data_463(mau_6_io_pipe_phv_out_data_463),
    .io_pipe_phv_out_data_464(mau_6_io_pipe_phv_out_data_464),
    .io_pipe_phv_out_data_465(mau_6_io_pipe_phv_out_data_465),
    .io_pipe_phv_out_data_466(mau_6_io_pipe_phv_out_data_466),
    .io_pipe_phv_out_data_467(mau_6_io_pipe_phv_out_data_467),
    .io_pipe_phv_out_data_468(mau_6_io_pipe_phv_out_data_468),
    .io_pipe_phv_out_data_469(mau_6_io_pipe_phv_out_data_469),
    .io_pipe_phv_out_data_470(mau_6_io_pipe_phv_out_data_470),
    .io_pipe_phv_out_data_471(mau_6_io_pipe_phv_out_data_471),
    .io_pipe_phv_out_data_472(mau_6_io_pipe_phv_out_data_472),
    .io_pipe_phv_out_data_473(mau_6_io_pipe_phv_out_data_473),
    .io_pipe_phv_out_data_474(mau_6_io_pipe_phv_out_data_474),
    .io_pipe_phv_out_data_475(mau_6_io_pipe_phv_out_data_475),
    .io_pipe_phv_out_data_476(mau_6_io_pipe_phv_out_data_476),
    .io_pipe_phv_out_data_477(mau_6_io_pipe_phv_out_data_477),
    .io_pipe_phv_out_data_478(mau_6_io_pipe_phv_out_data_478),
    .io_pipe_phv_out_data_479(mau_6_io_pipe_phv_out_data_479),
    .io_pipe_phv_out_data_480(mau_6_io_pipe_phv_out_data_480),
    .io_pipe_phv_out_data_481(mau_6_io_pipe_phv_out_data_481),
    .io_pipe_phv_out_data_482(mau_6_io_pipe_phv_out_data_482),
    .io_pipe_phv_out_data_483(mau_6_io_pipe_phv_out_data_483),
    .io_pipe_phv_out_data_484(mau_6_io_pipe_phv_out_data_484),
    .io_pipe_phv_out_data_485(mau_6_io_pipe_phv_out_data_485),
    .io_pipe_phv_out_data_486(mau_6_io_pipe_phv_out_data_486),
    .io_pipe_phv_out_data_487(mau_6_io_pipe_phv_out_data_487),
    .io_pipe_phv_out_data_488(mau_6_io_pipe_phv_out_data_488),
    .io_pipe_phv_out_data_489(mau_6_io_pipe_phv_out_data_489),
    .io_pipe_phv_out_data_490(mau_6_io_pipe_phv_out_data_490),
    .io_pipe_phv_out_data_491(mau_6_io_pipe_phv_out_data_491),
    .io_pipe_phv_out_data_492(mau_6_io_pipe_phv_out_data_492),
    .io_pipe_phv_out_data_493(mau_6_io_pipe_phv_out_data_493),
    .io_pipe_phv_out_data_494(mau_6_io_pipe_phv_out_data_494),
    .io_pipe_phv_out_data_495(mau_6_io_pipe_phv_out_data_495),
    .io_pipe_phv_out_data_496(mau_6_io_pipe_phv_out_data_496),
    .io_pipe_phv_out_data_497(mau_6_io_pipe_phv_out_data_497),
    .io_pipe_phv_out_data_498(mau_6_io_pipe_phv_out_data_498),
    .io_pipe_phv_out_data_499(mau_6_io_pipe_phv_out_data_499),
    .io_pipe_phv_out_data_500(mau_6_io_pipe_phv_out_data_500),
    .io_pipe_phv_out_data_501(mau_6_io_pipe_phv_out_data_501),
    .io_pipe_phv_out_data_502(mau_6_io_pipe_phv_out_data_502),
    .io_pipe_phv_out_data_503(mau_6_io_pipe_phv_out_data_503),
    .io_pipe_phv_out_data_504(mau_6_io_pipe_phv_out_data_504),
    .io_pipe_phv_out_data_505(mau_6_io_pipe_phv_out_data_505),
    .io_pipe_phv_out_data_506(mau_6_io_pipe_phv_out_data_506),
    .io_pipe_phv_out_data_507(mau_6_io_pipe_phv_out_data_507),
    .io_pipe_phv_out_data_508(mau_6_io_pipe_phv_out_data_508),
    .io_pipe_phv_out_data_509(mau_6_io_pipe_phv_out_data_509),
    .io_pipe_phv_out_data_510(mau_6_io_pipe_phv_out_data_510),
    .io_pipe_phv_out_data_511(mau_6_io_pipe_phv_out_data_511),
    .io_pipe_phv_out_header_0(mau_6_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(mau_6_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(mau_6_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(mau_6_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(mau_6_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(mau_6_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(mau_6_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(mau_6_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(mau_6_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(mau_6_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(mau_6_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(mau_6_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(mau_6_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(mau_6_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(mau_6_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(mau_6_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(mau_6_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(mau_6_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(mau_6_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(mau_6_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(mau_6_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(mau_6_io_pipe_phv_out_is_valid_processor),
    .io_mod_state_id_mod(mau_6_io_mod_state_id_mod),
    .io_mod_state_id(mau_6_io_mod_state_id),
    .io_mod_sram_w_cs(mau_6_io_mod_sram_w_cs),
    .io_mod_sram_w_en(mau_6_io_mod_sram_w_en),
    .io_mod_sram_w_addr(mau_6_io_mod_sram_w_addr),
    .io_mod_sram_w_data(mau_6_io_mod_sram_w_data)
  );
  ParseModule mau_7 ( // @[parser_pisa.scala 31:25]
    .clock(mau_7_clock),
    .io_pipe_phv_in_data_0(mau_7_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(mau_7_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(mau_7_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(mau_7_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(mau_7_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(mau_7_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(mau_7_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(mau_7_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(mau_7_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(mau_7_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(mau_7_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(mau_7_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(mau_7_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(mau_7_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(mau_7_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(mau_7_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(mau_7_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(mau_7_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(mau_7_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(mau_7_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(mau_7_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(mau_7_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(mau_7_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(mau_7_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(mau_7_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(mau_7_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(mau_7_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(mau_7_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(mau_7_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(mau_7_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(mau_7_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(mau_7_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(mau_7_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(mau_7_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(mau_7_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(mau_7_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(mau_7_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(mau_7_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(mau_7_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(mau_7_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(mau_7_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(mau_7_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(mau_7_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(mau_7_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(mau_7_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(mau_7_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(mau_7_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(mau_7_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(mau_7_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(mau_7_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(mau_7_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(mau_7_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(mau_7_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(mau_7_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(mau_7_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(mau_7_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(mau_7_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(mau_7_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(mau_7_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(mau_7_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(mau_7_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(mau_7_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(mau_7_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(mau_7_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(mau_7_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(mau_7_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(mau_7_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(mau_7_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(mau_7_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(mau_7_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(mau_7_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(mau_7_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(mau_7_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(mau_7_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(mau_7_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(mau_7_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(mau_7_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(mau_7_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(mau_7_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(mau_7_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(mau_7_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(mau_7_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(mau_7_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(mau_7_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(mau_7_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(mau_7_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(mau_7_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(mau_7_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(mau_7_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(mau_7_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(mau_7_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(mau_7_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(mau_7_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(mau_7_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(mau_7_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(mau_7_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(mau_7_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(mau_7_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(mau_7_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(mau_7_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(mau_7_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(mau_7_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(mau_7_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(mau_7_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(mau_7_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(mau_7_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(mau_7_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(mau_7_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(mau_7_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(mau_7_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(mau_7_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(mau_7_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(mau_7_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(mau_7_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(mau_7_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(mau_7_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(mau_7_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(mau_7_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(mau_7_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(mau_7_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(mau_7_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(mau_7_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(mau_7_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(mau_7_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(mau_7_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(mau_7_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(mau_7_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(mau_7_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(mau_7_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(mau_7_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(mau_7_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(mau_7_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(mau_7_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(mau_7_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(mau_7_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(mau_7_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(mau_7_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(mau_7_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(mau_7_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(mau_7_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(mau_7_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(mau_7_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(mau_7_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(mau_7_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(mau_7_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(mau_7_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(mau_7_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(mau_7_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(mau_7_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(mau_7_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(mau_7_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(mau_7_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(mau_7_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(mau_7_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(mau_7_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(mau_7_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(mau_7_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(mau_7_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(mau_7_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(mau_7_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(mau_7_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(mau_7_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(mau_7_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(mau_7_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(mau_7_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(mau_7_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(mau_7_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(mau_7_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(mau_7_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(mau_7_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(mau_7_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(mau_7_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(mau_7_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(mau_7_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(mau_7_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(mau_7_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(mau_7_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(mau_7_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(mau_7_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(mau_7_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(mau_7_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(mau_7_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(mau_7_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(mau_7_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(mau_7_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(mau_7_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(mau_7_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(mau_7_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(mau_7_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(mau_7_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(mau_7_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(mau_7_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(mau_7_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(mau_7_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(mau_7_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(mau_7_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(mau_7_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(mau_7_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(mau_7_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(mau_7_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(mau_7_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(mau_7_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(mau_7_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(mau_7_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(mau_7_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(mau_7_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(mau_7_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(mau_7_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(mau_7_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(mau_7_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(mau_7_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(mau_7_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(mau_7_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(mau_7_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(mau_7_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(mau_7_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(mau_7_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(mau_7_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(mau_7_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(mau_7_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(mau_7_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(mau_7_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(mau_7_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(mau_7_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(mau_7_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(mau_7_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(mau_7_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(mau_7_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(mau_7_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(mau_7_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(mau_7_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(mau_7_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(mau_7_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(mau_7_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(mau_7_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(mau_7_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(mau_7_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(mau_7_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(mau_7_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(mau_7_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(mau_7_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(mau_7_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(mau_7_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(mau_7_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(mau_7_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(mau_7_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(mau_7_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(mau_7_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(mau_7_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(mau_7_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(mau_7_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(mau_7_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(mau_7_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(mau_7_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(mau_7_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(mau_7_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_data_256(mau_7_io_pipe_phv_in_data_256),
    .io_pipe_phv_in_data_257(mau_7_io_pipe_phv_in_data_257),
    .io_pipe_phv_in_data_258(mau_7_io_pipe_phv_in_data_258),
    .io_pipe_phv_in_data_259(mau_7_io_pipe_phv_in_data_259),
    .io_pipe_phv_in_data_260(mau_7_io_pipe_phv_in_data_260),
    .io_pipe_phv_in_data_261(mau_7_io_pipe_phv_in_data_261),
    .io_pipe_phv_in_data_262(mau_7_io_pipe_phv_in_data_262),
    .io_pipe_phv_in_data_263(mau_7_io_pipe_phv_in_data_263),
    .io_pipe_phv_in_data_264(mau_7_io_pipe_phv_in_data_264),
    .io_pipe_phv_in_data_265(mau_7_io_pipe_phv_in_data_265),
    .io_pipe_phv_in_data_266(mau_7_io_pipe_phv_in_data_266),
    .io_pipe_phv_in_data_267(mau_7_io_pipe_phv_in_data_267),
    .io_pipe_phv_in_data_268(mau_7_io_pipe_phv_in_data_268),
    .io_pipe_phv_in_data_269(mau_7_io_pipe_phv_in_data_269),
    .io_pipe_phv_in_data_270(mau_7_io_pipe_phv_in_data_270),
    .io_pipe_phv_in_data_271(mau_7_io_pipe_phv_in_data_271),
    .io_pipe_phv_in_data_272(mau_7_io_pipe_phv_in_data_272),
    .io_pipe_phv_in_data_273(mau_7_io_pipe_phv_in_data_273),
    .io_pipe_phv_in_data_274(mau_7_io_pipe_phv_in_data_274),
    .io_pipe_phv_in_data_275(mau_7_io_pipe_phv_in_data_275),
    .io_pipe_phv_in_data_276(mau_7_io_pipe_phv_in_data_276),
    .io_pipe_phv_in_data_277(mau_7_io_pipe_phv_in_data_277),
    .io_pipe_phv_in_data_278(mau_7_io_pipe_phv_in_data_278),
    .io_pipe_phv_in_data_279(mau_7_io_pipe_phv_in_data_279),
    .io_pipe_phv_in_data_280(mau_7_io_pipe_phv_in_data_280),
    .io_pipe_phv_in_data_281(mau_7_io_pipe_phv_in_data_281),
    .io_pipe_phv_in_data_282(mau_7_io_pipe_phv_in_data_282),
    .io_pipe_phv_in_data_283(mau_7_io_pipe_phv_in_data_283),
    .io_pipe_phv_in_data_284(mau_7_io_pipe_phv_in_data_284),
    .io_pipe_phv_in_data_285(mau_7_io_pipe_phv_in_data_285),
    .io_pipe_phv_in_data_286(mau_7_io_pipe_phv_in_data_286),
    .io_pipe_phv_in_data_287(mau_7_io_pipe_phv_in_data_287),
    .io_pipe_phv_in_data_288(mau_7_io_pipe_phv_in_data_288),
    .io_pipe_phv_in_data_289(mau_7_io_pipe_phv_in_data_289),
    .io_pipe_phv_in_data_290(mau_7_io_pipe_phv_in_data_290),
    .io_pipe_phv_in_data_291(mau_7_io_pipe_phv_in_data_291),
    .io_pipe_phv_in_data_292(mau_7_io_pipe_phv_in_data_292),
    .io_pipe_phv_in_data_293(mau_7_io_pipe_phv_in_data_293),
    .io_pipe_phv_in_data_294(mau_7_io_pipe_phv_in_data_294),
    .io_pipe_phv_in_data_295(mau_7_io_pipe_phv_in_data_295),
    .io_pipe_phv_in_data_296(mau_7_io_pipe_phv_in_data_296),
    .io_pipe_phv_in_data_297(mau_7_io_pipe_phv_in_data_297),
    .io_pipe_phv_in_data_298(mau_7_io_pipe_phv_in_data_298),
    .io_pipe_phv_in_data_299(mau_7_io_pipe_phv_in_data_299),
    .io_pipe_phv_in_data_300(mau_7_io_pipe_phv_in_data_300),
    .io_pipe_phv_in_data_301(mau_7_io_pipe_phv_in_data_301),
    .io_pipe_phv_in_data_302(mau_7_io_pipe_phv_in_data_302),
    .io_pipe_phv_in_data_303(mau_7_io_pipe_phv_in_data_303),
    .io_pipe_phv_in_data_304(mau_7_io_pipe_phv_in_data_304),
    .io_pipe_phv_in_data_305(mau_7_io_pipe_phv_in_data_305),
    .io_pipe_phv_in_data_306(mau_7_io_pipe_phv_in_data_306),
    .io_pipe_phv_in_data_307(mau_7_io_pipe_phv_in_data_307),
    .io_pipe_phv_in_data_308(mau_7_io_pipe_phv_in_data_308),
    .io_pipe_phv_in_data_309(mau_7_io_pipe_phv_in_data_309),
    .io_pipe_phv_in_data_310(mau_7_io_pipe_phv_in_data_310),
    .io_pipe_phv_in_data_311(mau_7_io_pipe_phv_in_data_311),
    .io_pipe_phv_in_data_312(mau_7_io_pipe_phv_in_data_312),
    .io_pipe_phv_in_data_313(mau_7_io_pipe_phv_in_data_313),
    .io_pipe_phv_in_data_314(mau_7_io_pipe_phv_in_data_314),
    .io_pipe_phv_in_data_315(mau_7_io_pipe_phv_in_data_315),
    .io_pipe_phv_in_data_316(mau_7_io_pipe_phv_in_data_316),
    .io_pipe_phv_in_data_317(mau_7_io_pipe_phv_in_data_317),
    .io_pipe_phv_in_data_318(mau_7_io_pipe_phv_in_data_318),
    .io_pipe_phv_in_data_319(mau_7_io_pipe_phv_in_data_319),
    .io_pipe_phv_in_data_320(mau_7_io_pipe_phv_in_data_320),
    .io_pipe_phv_in_data_321(mau_7_io_pipe_phv_in_data_321),
    .io_pipe_phv_in_data_322(mau_7_io_pipe_phv_in_data_322),
    .io_pipe_phv_in_data_323(mau_7_io_pipe_phv_in_data_323),
    .io_pipe_phv_in_data_324(mau_7_io_pipe_phv_in_data_324),
    .io_pipe_phv_in_data_325(mau_7_io_pipe_phv_in_data_325),
    .io_pipe_phv_in_data_326(mau_7_io_pipe_phv_in_data_326),
    .io_pipe_phv_in_data_327(mau_7_io_pipe_phv_in_data_327),
    .io_pipe_phv_in_data_328(mau_7_io_pipe_phv_in_data_328),
    .io_pipe_phv_in_data_329(mau_7_io_pipe_phv_in_data_329),
    .io_pipe_phv_in_data_330(mau_7_io_pipe_phv_in_data_330),
    .io_pipe_phv_in_data_331(mau_7_io_pipe_phv_in_data_331),
    .io_pipe_phv_in_data_332(mau_7_io_pipe_phv_in_data_332),
    .io_pipe_phv_in_data_333(mau_7_io_pipe_phv_in_data_333),
    .io_pipe_phv_in_data_334(mau_7_io_pipe_phv_in_data_334),
    .io_pipe_phv_in_data_335(mau_7_io_pipe_phv_in_data_335),
    .io_pipe_phv_in_data_336(mau_7_io_pipe_phv_in_data_336),
    .io_pipe_phv_in_data_337(mau_7_io_pipe_phv_in_data_337),
    .io_pipe_phv_in_data_338(mau_7_io_pipe_phv_in_data_338),
    .io_pipe_phv_in_data_339(mau_7_io_pipe_phv_in_data_339),
    .io_pipe_phv_in_data_340(mau_7_io_pipe_phv_in_data_340),
    .io_pipe_phv_in_data_341(mau_7_io_pipe_phv_in_data_341),
    .io_pipe_phv_in_data_342(mau_7_io_pipe_phv_in_data_342),
    .io_pipe_phv_in_data_343(mau_7_io_pipe_phv_in_data_343),
    .io_pipe_phv_in_data_344(mau_7_io_pipe_phv_in_data_344),
    .io_pipe_phv_in_data_345(mau_7_io_pipe_phv_in_data_345),
    .io_pipe_phv_in_data_346(mau_7_io_pipe_phv_in_data_346),
    .io_pipe_phv_in_data_347(mau_7_io_pipe_phv_in_data_347),
    .io_pipe_phv_in_data_348(mau_7_io_pipe_phv_in_data_348),
    .io_pipe_phv_in_data_349(mau_7_io_pipe_phv_in_data_349),
    .io_pipe_phv_in_data_350(mau_7_io_pipe_phv_in_data_350),
    .io_pipe_phv_in_data_351(mau_7_io_pipe_phv_in_data_351),
    .io_pipe_phv_in_data_352(mau_7_io_pipe_phv_in_data_352),
    .io_pipe_phv_in_data_353(mau_7_io_pipe_phv_in_data_353),
    .io_pipe_phv_in_data_354(mau_7_io_pipe_phv_in_data_354),
    .io_pipe_phv_in_data_355(mau_7_io_pipe_phv_in_data_355),
    .io_pipe_phv_in_data_356(mau_7_io_pipe_phv_in_data_356),
    .io_pipe_phv_in_data_357(mau_7_io_pipe_phv_in_data_357),
    .io_pipe_phv_in_data_358(mau_7_io_pipe_phv_in_data_358),
    .io_pipe_phv_in_data_359(mau_7_io_pipe_phv_in_data_359),
    .io_pipe_phv_in_data_360(mau_7_io_pipe_phv_in_data_360),
    .io_pipe_phv_in_data_361(mau_7_io_pipe_phv_in_data_361),
    .io_pipe_phv_in_data_362(mau_7_io_pipe_phv_in_data_362),
    .io_pipe_phv_in_data_363(mau_7_io_pipe_phv_in_data_363),
    .io_pipe_phv_in_data_364(mau_7_io_pipe_phv_in_data_364),
    .io_pipe_phv_in_data_365(mau_7_io_pipe_phv_in_data_365),
    .io_pipe_phv_in_data_366(mau_7_io_pipe_phv_in_data_366),
    .io_pipe_phv_in_data_367(mau_7_io_pipe_phv_in_data_367),
    .io_pipe_phv_in_data_368(mau_7_io_pipe_phv_in_data_368),
    .io_pipe_phv_in_data_369(mau_7_io_pipe_phv_in_data_369),
    .io_pipe_phv_in_data_370(mau_7_io_pipe_phv_in_data_370),
    .io_pipe_phv_in_data_371(mau_7_io_pipe_phv_in_data_371),
    .io_pipe_phv_in_data_372(mau_7_io_pipe_phv_in_data_372),
    .io_pipe_phv_in_data_373(mau_7_io_pipe_phv_in_data_373),
    .io_pipe_phv_in_data_374(mau_7_io_pipe_phv_in_data_374),
    .io_pipe_phv_in_data_375(mau_7_io_pipe_phv_in_data_375),
    .io_pipe_phv_in_data_376(mau_7_io_pipe_phv_in_data_376),
    .io_pipe_phv_in_data_377(mau_7_io_pipe_phv_in_data_377),
    .io_pipe_phv_in_data_378(mau_7_io_pipe_phv_in_data_378),
    .io_pipe_phv_in_data_379(mau_7_io_pipe_phv_in_data_379),
    .io_pipe_phv_in_data_380(mau_7_io_pipe_phv_in_data_380),
    .io_pipe_phv_in_data_381(mau_7_io_pipe_phv_in_data_381),
    .io_pipe_phv_in_data_382(mau_7_io_pipe_phv_in_data_382),
    .io_pipe_phv_in_data_383(mau_7_io_pipe_phv_in_data_383),
    .io_pipe_phv_in_data_384(mau_7_io_pipe_phv_in_data_384),
    .io_pipe_phv_in_data_385(mau_7_io_pipe_phv_in_data_385),
    .io_pipe_phv_in_data_386(mau_7_io_pipe_phv_in_data_386),
    .io_pipe_phv_in_data_387(mau_7_io_pipe_phv_in_data_387),
    .io_pipe_phv_in_data_388(mau_7_io_pipe_phv_in_data_388),
    .io_pipe_phv_in_data_389(mau_7_io_pipe_phv_in_data_389),
    .io_pipe_phv_in_data_390(mau_7_io_pipe_phv_in_data_390),
    .io_pipe_phv_in_data_391(mau_7_io_pipe_phv_in_data_391),
    .io_pipe_phv_in_data_392(mau_7_io_pipe_phv_in_data_392),
    .io_pipe_phv_in_data_393(mau_7_io_pipe_phv_in_data_393),
    .io_pipe_phv_in_data_394(mau_7_io_pipe_phv_in_data_394),
    .io_pipe_phv_in_data_395(mau_7_io_pipe_phv_in_data_395),
    .io_pipe_phv_in_data_396(mau_7_io_pipe_phv_in_data_396),
    .io_pipe_phv_in_data_397(mau_7_io_pipe_phv_in_data_397),
    .io_pipe_phv_in_data_398(mau_7_io_pipe_phv_in_data_398),
    .io_pipe_phv_in_data_399(mau_7_io_pipe_phv_in_data_399),
    .io_pipe_phv_in_data_400(mau_7_io_pipe_phv_in_data_400),
    .io_pipe_phv_in_data_401(mau_7_io_pipe_phv_in_data_401),
    .io_pipe_phv_in_data_402(mau_7_io_pipe_phv_in_data_402),
    .io_pipe_phv_in_data_403(mau_7_io_pipe_phv_in_data_403),
    .io_pipe_phv_in_data_404(mau_7_io_pipe_phv_in_data_404),
    .io_pipe_phv_in_data_405(mau_7_io_pipe_phv_in_data_405),
    .io_pipe_phv_in_data_406(mau_7_io_pipe_phv_in_data_406),
    .io_pipe_phv_in_data_407(mau_7_io_pipe_phv_in_data_407),
    .io_pipe_phv_in_data_408(mau_7_io_pipe_phv_in_data_408),
    .io_pipe_phv_in_data_409(mau_7_io_pipe_phv_in_data_409),
    .io_pipe_phv_in_data_410(mau_7_io_pipe_phv_in_data_410),
    .io_pipe_phv_in_data_411(mau_7_io_pipe_phv_in_data_411),
    .io_pipe_phv_in_data_412(mau_7_io_pipe_phv_in_data_412),
    .io_pipe_phv_in_data_413(mau_7_io_pipe_phv_in_data_413),
    .io_pipe_phv_in_data_414(mau_7_io_pipe_phv_in_data_414),
    .io_pipe_phv_in_data_415(mau_7_io_pipe_phv_in_data_415),
    .io_pipe_phv_in_data_416(mau_7_io_pipe_phv_in_data_416),
    .io_pipe_phv_in_data_417(mau_7_io_pipe_phv_in_data_417),
    .io_pipe_phv_in_data_418(mau_7_io_pipe_phv_in_data_418),
    .io_pipe_phv_in_data_419(mau_7_io_pipe_phv_in_data_419),
    .io_pipe_phv_in_data_420(mau_7_io_pipe_phv_in_data_420),
    .io_pipe_phv_in_data_421(mau_7_io_pipe_phv_in_data_421),
    .io_pipe_phv_in_data_422(mau_7_io_pipe_phv_in_data_422),
    .io_pipe_phv_in_data_423(mau_7_io_pipe_phv_in_data_423),
    .io_pipe_phv_in_data_424(mau_7_io_pipe_phv_in_data_424),
    .io_pipe_phv_in_data_425(mau_7_io_pipe_phv_in_data_425),
    .io_pipe_phv_in_data_426(mau_7_io_pipe_phv_in_data_426),
    .io_pipe_phv_in_data_427(mau_7_io_pipe_phv_in_data_427),
    .io_pipe_phv_in_data_428(mau_7_io_pipe_phv_in_data_428),
    .io_pipe_phv_in_data_429(mau_7_io_pipe_phv_in_data_429),
    .io_pipe_phv_in_data_430(mau_7_io_pipe_phv_in_data_430),
    .io_pipe_phv_in_data_431(mau_7_io_pipe_phv_in_data_431),
    .io_pipe_phv_in_data_432(mau_7_io_pipe_phv_in_data_432),
    .io_pipe_phv_in_data_433(mau_7_io_pipe_phv_in_data_433),
    .io_pipe_phv_in_data_434(mau_7_io_pipe_phv_in_data_434),
    .io_pipe_phv_in_data_435(mau_7_io_pipe_phv_in_data_435),
    .io_pipe_phv_in_data_436(mau_7_io_pipe_phv_in_data_436),
    .io_pipe_phv_in_data_437(mau_7_io_pipe_phv_in_data_437),
    .io_pipe_phv_in_data_438(mau_7_io_pipe_phv_in_data_438),
    .io_pipe_phv_in_data_439(mau_7_io_pipe_phv_in_data_439),
    .io_pipe_phv_in_data_440(mau_7_io_pipe_phv_in_data_440),
    .io_pipe_phv_in_data_441(mau_7_io_pipe_phv_in_data_441),
    .io_pipe_phv_in_data_442(mau_7_io_pipe_phv_in_data_442),
    .io_pipe_phv_in_data_443(mau_7_io_pipe_phv_in_data_443),
    .io_pipe_phv_in_data_444(mau_7_io_pipe_phv_in_data_444),
    .io_pipe_phv_in_data_445(mau_7_io_pipe_phv_in_data_445),
    .io_pipe_phv_in_data_446(mau_7_io_pipe_phv_in_data_446),
    .io_pipe_phv_in_data_447(mau_7_io_pipe_phv_in_data_447),
    .io_pipe_phv_in_data_448(mau_7_io_pipe_phv_in_data_448),
    .io_pipe_phv_in_data_449(mau_7_io_pipe_phv_in_data_449),
    .io_pipe_phv_in_data_450(mau_7_io_pipe_phv_in_data_450),
    .io_pipe_phv_in_data_451(mau_7_io_pipe_phv_in_data_451),
    .io_pipe_phv_in_data_452(mau_7_io_pipe_phv_in_data_452),
    .io_pipe_phv_in_data_453(mau_7_io_pipe_phv_in_data_453),
    .io_pipe_phv_in_data_454(mau_7_io_pipe_phv_in_data_454),
    .io_pipe_phv_in_data_455(mau_7_io_pipe_phv_in_data_455),
    .io_pipe_phv_in_data_456(mau_7_io_pipe_phv_in_data_456),
    .io_pipe_phv_in_data_457(mau_7_io_pipe_phv_in_data_457),
    .io_pipe_phv_in_data_458(mau_7_io_pipe_phv_in_data_458),
    .io_pipe_phv_in_data_459(mau_7_io_pipe_phv_in_data_459),
    .io_pipe_phv_in_data_460(mau_7_io_pipe_phv_in_data_460),
    .io_pipe_phv_in_data_461(mau_7_io_pipe_phv_in_data_461),
    .io_pipe_phv_in_data_462(mau_7_io_pipe_phv_in_data_462),
    .io_pipe_phv_in_data_463(mau_7_io_pipe_phv_in_data_463),
    .io_pipe_phv_in_data_464(mau_7_io_pipe_phv_in_data_464),
    .io_pipe_phv_in_data_465(mau_7_io_pipe_phv_in_data_465),
    .io_pipe_phv_in_data_466(mau_7_io_pipe_phv_in_data_466),
    .io_pipe_phv_in_data_467(mau_7_io_pipe_phv_in_data_467),
    .io_pipe_phv_in_data_468(mau_7_io_pipe_phv_in_data_468),
    .io_pipe_phv_in_data_469(mau_7_io_pipe_phv_in_data_469),
    .io_pipe_phv_in_data_470(mau_7_io_pipe_phv_in_data_470),
    .io_pipe_phv_in_data_471(mau_7_io_pipe_phv_in_data_471),
    .io_pipe_phv_in_data_472(mau_7_io_pipe_phv_in_data_472),
    .io_pipe_phv_in_data_473(mau_7_io_pipe_phv_in_data_473),
    .io_pipe_phv_in_data_474(mau_7_io_pipe_phv_in_data_474),
    .io_pipe_phv_in_data_475(mau_7_io_pipe_phv_in_data_475),
    .io_pipe_phv_in_data_476(mau_7_io_pipe_phv_in_data_476),
    .io_pipe_phv_in_data_477(mau_7_io_pipe_phv_in_data_477),
    .io_pipe_phv_in_data_478(mau_7_io_pipe_phv_in_data_478),
    .io_pipe_phv_in_data_479(mau_7_io_pipe_phv_in_data_479),
    .io_pipe_phv_in_data_480(mau_7_io_pipe_phv_in_data_480),
    .io_pipe_phv_in_data_481(mau_7_io_pipe_phv_in_data_481),
    .io_pipe_phv_in_data_482(mau_7_io_pipe_phv_in_data_482),
    .io_pipe_phv_in_data_483(mau_7_io_pipe_phv_in_data_483),
    .io_pipe_phv_in_data_484(mau_7_io_pipe_phv_in_data_484),
    .io_pipe_phv_in_data_485(mau_7_io_pipe_phv_in_data_485),
    .io_pipe_phv_in_data_486(mau_7_io_pipe_phv_in_data_486),
    .io_pipe_phv_in_data_487(mau_7_io_pipe_phv_in_data_487),
    .io_pipe_phv_in_data_488(mau_7_io_pipe_phv_in_data_488),
    .io_pipe_phv_in_data_489(mau_7_io_pipe_phv_in_data_489),
    .io_pipe_phv_in_data_490(mau_7_io_pipe_phv_in_data_490),
    .io_pipe_phv_in_data_491(mau_7_io_pipe_phv_in_data_491),
    .io_pipe_phv_in_data_492(mau_7_io_pipe_phv_in_data_492),
    .io_pipe_phv_in_data_493(mau_7_io_pipe_phv_in_data_493),
    .io_pipe_phv_in_data_494(mau_7_io_pipe_phv_in_data_494),
    .io_pipe_phv_in_data_495(mau_7_io_pipe_phv_in_data_495),
    .io_pipe_phv_in_data_496(mau_7_io_pipe_phv_in_data_496),
    .io_pipe_phv_in_data_497(mau_7_io_pipe_phv_in_data_497),
    .io_pipe_phv_in_data_498(mau_7_io_pipe_phv_in_data_498),
    .io_pipe_phv_in_data_499(mau_7_io_pipe_phv_in_data_499),
    .io_pipe_phv_in_data_500(mau_7_io_pipe_phv_in_data_500),
    .io_pipe_phv_in_data_501(mau_7_io_pipe_phv_in_data_501),
    .io_pipe_phv_in_data_502(mau_7_io_pipe_phv_in_data_502),
    .io_pipe_phv_in_data_503(mau_7_io_pipe_phv_in_data_503),
    .io_pipe_phv_in_data_504(mau_7_io_pipe_phv_in_data_504),
    .io_pipe_phv_in_data_505(mau_7_io_pipe_phv_in_data_505),
    .io_pipe_phv_in_data_506(mau_7_io_pipe_phv_in_data_506),
    .io_pipe_phv_in_data_507(mau_7_io_pipe_phv_in_data_507),
    .io_pipe_phv_in_data_508(mau_7_io_pipe_phv_in_data_508),
    .io_pipe_phv_in_data_509(mau_7_io_pipe_phv_in_data_509),
    .io_pipe_phv_in_data_510(mau_7_io_pipe_phv_in_data_510),
    .io_pipe_phv_in_data_511(mau_7_io_pipe_phv_in_data_511),
    .io_pipe_phv_in_header_0(mau_7_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(mau_7_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(mau_7_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(mau_7_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(mau_7_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(mau_7_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(mau_7_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(mau_7_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(mau_7_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(mau_7_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(mau_7_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(mau_7_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(mau_7_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(mau_7_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(mau_7_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(mau_7_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(mau_7_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(mau_7_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(mau_7_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(mau_7_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(mau_7_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(mau_7_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(mau_7_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(mau_7_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(mau_7_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(mau_7_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(mau_7_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(mau_7_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(mau_7_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(mau_7_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(mau_7_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(mau_7_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(mau_7_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(mau_7_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(mau_7_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(mau_7_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(mau_7_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(mau_7_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(mau_7_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(mau_7_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(mau_7_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(mau_7_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(mau_7_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(mau_7_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(mau_7_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(mau_7_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(mau_7_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(mau_7_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(mau_7_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(mau_7_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(mau_7_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(mau_7_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(mau_7_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(mau_7_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(mau_7_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(mau_7_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(mau_7_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(mau_7_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(mau_7_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(mau_7_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(mau_7_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(mau_7_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(mau_7_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(mau_7_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(mau_7_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(mau_7_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(mau_7_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(mau_7_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(mau_7_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(mau_7_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(mau_7_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(mau_7_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(mau_7_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(mau_7_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(mau_7_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(mau_7_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(mau_7_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(mau_7_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(mau_7_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(mau_7_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(mau_7_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(mau_7_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(mau_7_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(mau_7_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(mau_7_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(mau_7_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(mau_7_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(mau_7_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(mau_7_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(mau_7_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(mau_7_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(mau_7_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(mau_7_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(mau_7_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(mau_7_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(mau_7_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(mau_7_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(mau_7_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(mau_7_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(mau_7_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(mau_7_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(mau_7_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(mau_7_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(mau_7_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(mau_7_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(mau_7_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(mau_7_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(mau_7_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(mau_7_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(mau_7_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(mau_7_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(mau_7_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(mau_7_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(mau_7_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(mau_7_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(mau_7_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(mau_7_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(mau_7_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(mau_7_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(mau_7_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(mau_7_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(mau_7_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(mau_7_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(mau_7_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(mau_7_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(mau_7_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(mau_7_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(mau_7_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(mau_7_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(mau_7_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(mau_7_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(mau_7_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(mau_7_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(mau_7_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(mau_7_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(mau_7_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(mau_7_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(mau_7_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(mau_7_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(mau_7_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(mau_7_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(mau_7_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(mau_7_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(mau_7_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(mau_7_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(mau_7_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(mau_7_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(mau_7_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(mau_7_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(mau_7_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(mau_7_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(mau_7_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(mau_7_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(mau_7_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(mau_7_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(mau_7_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(mau_7_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(mau_7_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(mau_7_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(mau_7_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(mau_7_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(mau_7_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(mau_7_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(mau_7_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(mau_7_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(mau_7_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(mau_7_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(mau_7_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(mau_7_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(mau_7_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(mau_7_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(mau_7_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(mau_7_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(mau_7_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(mau_7_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(mau_7_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(mau_7_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(mau_7_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(mau_7_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(mau_7_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(mau_7_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(mau_7_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(mau_7_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(mau_7_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(mau_7_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(mau_7_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(mau_7_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(mau_7_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(mau_7_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(mau_7_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(mau_7_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(mau_7_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(mau_7_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(mau_7_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(mau_7_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(mau_7_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(mau_7_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(mau_7_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(mau_7_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(mau_7_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(mau_7_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(mau_7_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(mau_7_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(mau_7_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(mau_7_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(mau_7_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(mau_7_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(mau_7_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(mau_7_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(mau_7_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(mau_7_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(mau_7_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(mau_7_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(mau_7_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(mau_7_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(mau_7_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(mau_7_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(mau_7_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(mau_7_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(mau_7_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(mau_7_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(mau_7_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(mau_7_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(mau_7_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(mau_7_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(mau_7_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(mau_7_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(mau_7_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(mau_7_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(mau_7_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(mau_7_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(mau_7_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(mau_7_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(mau_7_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(mau_7_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(mau_7_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(mau_7_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(mau_7_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(mau_7_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(mau_7_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(mau_7_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(mau_7_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(mau_7_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(mau_7_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(mau_7_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(mau_7_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(mau_7_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(mau_7_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(mau_7_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(mau_7_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(mau_7_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(mau_7_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(mau_7_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(mau_7_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(mau_7_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(mau_7_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(mau_7_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(mau_7_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(mau_7_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(mau_7_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(mau_7_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(mau_7_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(mau_7_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(mau_7_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(mau_7_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(mau_7_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(mau_7_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(mau_7_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(mau_7_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(mau_7_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(mau_7_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(mau_7_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(mau_7_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(mau_7_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(mau_7_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(mau_7_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(mau_7_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(mau_7_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_data_256(mau_7_io_pipe_phv_out_data_256),
    .io_pipe_phv_out_data_257(mau_7_io_pipe_phv_out_data_257),
    .io_pipe_phv_out_data_258(mau_7_io_pipe_phv_out_data_258),
    .io_pipe_phv_out_data_259(mau_7_io_pipe_phv_out_data_259),
    .io_pipe_phv_out_data_260(mau_7_io_pipe_phv_out_data_260),
    .io_pipe_phv_out_data_261(mau_7_io_pipe_phv_out_data_261),
    .io_pipe_phv_out_data_262(mau_7_io_pipe_phv_out_data_262),
    .io_pipe_phv_out_data_263(mau_7_io_pipe_phv_out_data_263),
    .io_pipe_phv_out_data_264(mau_7_io_pipe_phv_out_data_264),
    .io_pipe_phv_out_data_265(mau_7_io_pipe_phv_out_data_265),
    .io_pipe_phv_out_data_266(mau_7_io_pipe_phv_out_data_266),
    .io_pipe_phv_out_data_267(mau_7_io_pipe_phv_out_data_267),
    .io_pipe_phv_out_data_268(mau_7_io_pipe_phv_out_data_268),
    .io_pipe_phv_out_data_269(mau_7_io_pipe_phv_out_data_269),
    .io_pipe_phv_out_data_270(mau_7_io_pipe_phv_out_data_270),
    .io_pipe_phv_out_data_271(mau_7_io_pipe_phv_out_data_271),
    .io_pipe_phv_out_data_272(mau_7_io_pipe_phv_out_data_272),
    .io_pipe_phv_out_data_273(mau_7_io_pipe_phv_out_data_273),
    .io_pipe_phv_out_data_274(mau_7_io_pipe_phv_out_data_274),
    .io_pipe_phv_out_data_275(mau_7_io_pipe_phv_out_data_275),
    .io_pipe_phv_out_data_276(mau_7_io_pipe_phv_out_data_276),
    .io_pipe_phv_out_data_277(mau_7_io_pipe_phv_out_data_277),
    .io_pipe_phv_out_data_278(mau_7_io_pipe_phv_out_data_278),
    .io_pipe_phv_out_data_279(mau_7_io_pipe_phv_out_data_279),
    .io_pipe_phv_out_data_280(mau_7_io_pipe_phv_out_data_280),
    .io_pipe_phv_out_data_281(mau_7_io_pipe_phv_out_data_281),
    .io_pipe_phv_out_data_282(mau_7_io_pipe_phv_out_data_282),
    .io_pipe_phv_out_data_283(mau_7_io_pipe_phv_out_data_283),
    .io_pipe_phv_out_data_284(mau_7_io_pipe_phv_out_data_284),
    .io_pipe_phv_out_data_285(mau_7_io_pipe_phv_out_data_285),
    .io_pipe_phv_out_data_286(mau_7_io_pipe_phv_out_data_286),
    .io_pipe_phv_out_data_287(mau_7_io_pipe_phv_out_data_287),
    .io_pipe_phv_out_data_288(mau_7_io_pipe_phv_out_data_288),
    .io_pipe_phv_out_data_289(mau_7_io_pipe_phv_out_data_289),
    .io_pipe_phv_out_data_290(mau_7_io_pipe_phv_out_data_290),
    .io_pipe_phv_out_data_291(mau_7_io_pipe_phv_out_data_291),
    .io_pipe_phv_out_data_292(mau_7_io_pipe_phv_out_data_292),
    .io_pipe_phv_out_data_293(mau_7_io_pipe_phv_out_data_293),
    .io_pipe_phv_out_data_294(mau_7_io_pipe_phv_out_data_294),
    .io_pipe_phv_out_data_295(mau_7_io_pipe_phv_out_data_295),
    .io_pipe_phv_out_data_296(mau_7_io_pipe_phv_out_data_296),
    .io_pipe_phv_out_data_297(mau_7_io_pipe_phv_out_data_297),
    .io_pipe_phv_out_data_298(mau_7_io_pipe_phv_out_data_298),
    .io_pipe_phv_out_data_299(mau_7_io_pipe_phv_out_data_299),
    .io_pipe_phv_out_data_300(mau_7_io_pipe_phv_out_data_300),
    .io_pipe_phv_out_data_301(mau_7_io_pipe_phv_out_data_301),
    .io_pipe_phv_out_data_302(mau_7_io_pipe_phv_out_data_302),
    .io_pipe_phv_out_data_303(mau_7_io_pipe_phv_out_data_303),
    .io_pipe_phv_out_data_304(mau_7_io_pipe_phv_out_data_304),
    .io_pipe_phv_out_data_305(mau_7_io_pipe_phv_out_data_305),
    .io_pipe_phv_out_data_306(mau_7_io_pipe_phv_out_data_306),
    .io_pipe_phv_out_data_307(mau_7_io_pipe_phv_out_data_307),
    .io_pipe_phv_out_data_308(mau_7_io_pipe_phv_out_data_308),
    .io_pipe_phv_out_data_309(mau_7_io_pipe_phv_out_data_309),
    .io_pipe_phv_out_data_310(mau_7_io_pipe_phv_out_data_310),
    .io_pipe_phv_out_data_311(mau_7_io_pipe_phv_out_data_311),
    .io_pipe_phv_out_data_312(mau_7_io_pipe_phv_out_data_312),
    .io_pipe_phv_out_data_313(mau_7_io_pipe_phv_out_data_313),
    .io_pipe_phv_out_data_314(mau_7_io_pipe_phv_out_data_314),
    .io_pipe_phv_out_data_315(mau_7_io_pipe_phv_out_data_315),
    .io_pipe_phv_out_data_316(mau_7_io_pipe_phv_out_data_316),
    .io_pipe_phv_out_data_317(mau_7_io_pipe_phv_out_data_317),
    .io_pipe_phv_out_data_318(mau_7_io_pipe_phv_out_data_318),
    .io_pipe_phv_out_data_319(mau_7_io_pipe_phv_out_data_319),
    .io_pipe_phv_out_data_320(mau_7_io_pipe_phv_out_data_320),
    .io_pipe_phv_out_data_321(mau_7_io_pipe_phv_out_data_321),
    .io_pipe_phv_out_data_322(mau_7_io_pipe_phv_out_data_322),
    .io_pipe_phv_out_data_323(mau_7_io_pipe_phv_out_data_323),
    .io_pipe_phv_out_data_324(mau_7_io_pipe_phv_out_data_324),
    .io_pipe_phv_out_data_325(mau_7_io_pipe_phv_out_data_325),
    .io_pipe_phv_out_data_326(mau_7_io_pipe_phv_out_data_326),
    .io_pipe_phv_out_data_327(mau_7_io_pipe_phv_out_data_327),
    .io_pipe_phv_out_data_328(mau_7_io_pipe_phv_out_data_328),
    .io_pipe_phv_out_data_329(mau_7_io_pipe_phv_out_data_329),
    .io_pipe_phv_out_data_330(mau_7_io_pipe_phv_out_data_330),
    .io_pipe_phv_out_data_331(mau_7_io_pipe_phv_out_data_331),
    .io_pipe_phv_out_data_332(mau_7_io_pipe_phv_out_data_332),
    .io_pipe_phv_out_data_333(mau_7_io_pipe_phv_out_data_333),
    .io_pipe_phv_out_data_334(mau_7_io_pipe_phv_out_data_334),
    .io_pipe_phv_out_data_335(mau_7_io_pipe_phv_out_data_335),
    .io_pipe_phv_out_data_336(mau_7_io_pipe_phv_out_data_336),
    .io_pipe_phv_out_data_337(mau_7_io_pipe_phv_out_data_337),
    .io_pipe_phv_out_data_338(mau_7_io_pipe_phv_out_data_338),
    .io_pipe_phv_out_data_339(mau_7_io_pipe_phv_out_data_339),
    .io_pipe_phv_out_data_340(mau_7_io_pipe_phv_out_data_340),
    .io_pipe_phv_out_data_341(mau_7_io_pipe_phv_out_data_341),
    .io_pipe_phv_out_data_342(mau_7_io_pipe_phv_out_data_342),
    .io_pipe_phv_out_data_343(mau_7_io_pipe_phv_out_data_343),
    .io_pipe_phv_out_data_344(mau_7_io_pipe_phv_out_data_344),
    .io_pipe_phv_out_data_345(mau_7_io_pipe_phv_out_data_345),
    .io_pipe_phv_out_data_346(mau_7_io_pipe_phv_out_data_346),
    .io_pipe_phv_out_data_347(mau_7_io_pipe_phv_out_data_347),
    .io_pipe_phv_out_data_348(mau_7_io_pipe_phv_out_data_348),
    .io_pipe_phv_out_data_349(mau_7_io_pipe_phv_out_data_349),
    .io_pipe_phv_out_data_350(mau_7_io_pipe_phv_out_data_350),
    .io_pipe_phv_out_data_351(mau_7_io_pipe_phv_out_data_351),
    .io_pipe_phv_out_data_352(mau_7_io_pipe_phv_out_data_352),
    .io_pipe_phv_out_data_353(mau_7_io_pipe_phv_out_data_353),
    .io_pipe_phv_out_data_354(mau_7_io_pipe_phv_out_data_354),
    .io_pipe_phv_out_data_355(mau_7_io_pipe_phv_out_data_355),
    .io_pipe_phv_out_data_356(mau_7_io_pipe_phv_out_data_356),
    .io_pipe_phv_out_data_357(mau_7_io_pipe_phv_out_data_357),
    .io_pipe_phv_out_data_358(mau_7_io_pipe_phv_out_data_358),
    .io_pipe_phv_out_data_359(mau_7_io_pipe_phv_out_data_359),
    .io_pipe_phv_out_data_360(mau_7_io_pipe_phv_out_data_360),
    .io_pipe_phv_out_data_361(mau_7_io_pipe_phv_out_data_361),
    .io_pipe_phv_out_data_362(mau_7_io_pipe_phv_out_data_362),
    .io_pipe_phv_out_data_363(mau_7_io_pipe_phv_out_data_363),
    .io_pipe_phv_out_data_364(mau_7_io_pipe_phv_out_data_364),
    .io_pipe_phv_out_data_365(mau_7_io_pipe_phv_out_data_365),
    .io_pipe_phv_out_data_366(mau_7_io_pipe_phv_out_data_366),
    .io_pipe_phv_out_data_367(mau_7_io_pipe_phv_out_data_367),
    .io_pipe_phv_out_data_368(mau_7_io_pipe_phv_out_data_368),
    .io_pipe_phv_out_data_369(mau_7_io_pipe_phv_out_data_369),
    .io_pipe_phv_out_data_370(mau_7_io_pipe_phv_out_data_370),
    .io_pipe_phv_out_data_371(mau_7_io_pipe_phv_out_data_371),
    .io_pipe_phv_out_data_372(mau_7_io_pipe_phv_out_data_372),
    .io_pipe_phv_out_data_373(mau_7_io_pipe_phv_out_data_373),
    .io_pipe_phv_out_data_374(mau_7_io_pipe_phv_out_data_374),
    .io_pipe_phv_out_data_375(mau_7_io_pipe_phv_out_data_375),
    .io_pipe_phv_out_data_376(mau_7_io_pipe_phv_out_data_376),
    .io_pipe_phv_out_data_377(mau_7_io_pipe_phv_out_data_377),
    .io_pipe_phv_out_data_378(mau_7_io_pipe_phv_out_data_378),
    .io_pipe_phv_out_data_379(mau_7_io_pipe_phv_out_data_379),
    .io_pipe_phv_out_data_380(mau_7_io_pipe_phv_out_data_380),
    .io_pipe_phv_out_data_381(mau_7_io_pipe_phv_out_data_381),
    .io_pipe_phv_out_data_382(mau_7_io_pipe_phv_out_data_382),
    .io_pipe_phv_out_data_383(mau_7_io_pipe_phv_out_data_383),
    .io_pipe_phv_out_data_384(mau_7_io_pipe_phv_out_data_384),
    .io_pipe_phv_out_data_385(mau_7_io_pipe_phv_out_data_385),
    .io_pipe_phv_out_data_386(mau_7_io_pipe_phv_out_data_386),
    .io_pipe_phv_out_data_387(mau_7_io_pipe_phv_out_data_387),
    .io_pipe_phv_out_data_388(mau_7_io_pipe_phv_out_data_388),
    .io_pipe_phv_out_data_389(mau_7_io_pipe_phv_out_data_389),
    .io_pipe_phv_out_data_390(mau_7_io_pipe_phv_out_data_390),
    .io_pipe_phv_out_data_391(mau_7_io_pipe_phv_out_data_391),
    .io_pipe_phv_out_data_392(mau_7_io_pipe_phv_out_data_392),
    .io_pipe_phv_out_data_393(mau_7_io_pipe_phv_out_data_393),
    .io_pipe_phv_out_data_394(mau_7_io_pipe_phv_out_data_394),
    .io_pipe_phv_out_data_395(mau_7_io_pipe_phv_out_data_395),
    .io_pipe_phv_out_data_396(mau_7_io_pipe_phv_out_data_396),
    .io_pipe_phv_out_data_397(mau_7_io_pipe_phv_out_data_397),
    .io_pipe_phv_out_data_398(mau_7_io_pipe_phv_out_data_398),
    .io_pipe_phv_out_data_399(mau_7_io_pipe_phv_out_data_399),
    .io_pipe_phv_out_data_400(mau_7_io_pipe_phv_out_data_400),
    .io_pipe_phv_out_data_401(mau_7_io_pipe_phv_out_data_401),
    .io_pipe_phv_out_data_402(mau_7_io_pipe_phv_out_data_402),
    .io_pipe_phv_out_data_403(mau_7_io_pipe_phv_out_data_403),
    .io_pipe_phv_out_data_404(mau_7_io_pipe_phv_out_data_404),
    .io_pipe_phv_out_data_405(mau_7_io_pipe_phv_out_data_405),
    .io_pipe_phv_out_data_406(mau_7_io_pipe_phv_out_data_406),
    .io_pipe_phv_out_data_407(mau_7_io_pipe_phv_out_data_407),
    .io_pipe_phv_out_data_408(mau_7_io_pipe_phv_out_data_408),
    .io_pipe_phv_out_data_409(mau_7_io_pipe_phv_out_data_409),
    .io_pipe_phv_out_data_410(mau_7_io_pipe_phv_out_data_410),
    .io_pipe_phv_out_data_411(mau_7_io_pipe_phv_out_data_411),
    .io_pipe_phv_out_data_412(mau_7_io_pipe_phv_out_data_412),
    .io_pipe_phv_out_data_413(mau_7_io_pipe_phv_out_data_413),
    .io_pipe_phv_out_data_414(mau_7_io_pipe_phv_out_data_414),
    .io_pipe_phv_out_data_415(mau_7_io_pipe_phv_out_data_415),
    .io_pipe_phv_out_data_416(mau_7_io_pipe_phv_out_data_416),
    .io_pipe_phv_out_data_417(mau_7_io_pipe_phv_out_data_417),
    .io_pipe_phv_out_data_418(mau_7_io_pipe_phv_out_data_418),
    .io_pipe_phv_out_data_419(mau_7_io_pipe_phv_out_data_419),
    .io_pipe_phv_out_data_420(mau_7_io_pipe_phv_out_data_420),
    .io_pipe_phv_out_data_421(mau_7_io_pipe_phv_out_data_421),
    .io_pipe_phv_out_data_422(mau_7_io_pipe_phv_out_data_422),
    .io_pipe_phv_out_data_423(mau_7_io_pipe_phv_out_data_423),
    .io_pipe_phv_out_data_424(mau_7_io_pipe_phv_out_data_424),
    .io_pipe_phv_out_data_425(mau_7_io_pipe_phv_out_data_425),
    .io_pipe_phv_out_data_426(mau_7_io_pipe_phv_out_data_426),
    .io_pipe_phv_out_data_427(mau_7_io_pipe_phv_out_data_427),
    .io_pipe_phv_out_data_428(mau_7_io_pipe_phv_out_data_428),
    .io_pipe_phv_out_data_429(mau_7_io_pipe_phv_out_data_429),
    .io_pipe_phv_out_data_430(mau_7_io_pipe_phv_out_data_430),
    .io_pipe_phv_out_data_431(mau_7_io_pipe_phv_out_data_431),
    .io_pipe_phv_out_data_432(mau_7_io_pipe_phv_out_data_432),
    .io_pipe_phv_out_data_433(mau_7_io_pipe_phv_out_data_433),
    .io_pipe_phv_out_data_434(mau_7_io_pipe_phv_out_data_434),
    .io_pipe_phv_out_data_435(mau_7_io_pipe_phv_out_data_435),
    .io_pipe_phv_out_data_436(mau_7_io_pipe_phv_out_data_436),
    .io_pipe_phv_out_data_437(mau_7_io_pipe_phv_out_data_437),
    .io_pipe_phv_out_data_438(mau_7_io_pipe_phv_out_data_438),
    .io_pipe_phv_out_data_439(mau_7_io_pipe_phv_out_data_439),
    .io_pipe_phv_out_data_440(mau_7_io_pipe_phv_out_data_440),
    .io_pipe_phv_out_data_441(mau_7_io_pipe_phv_out_data_441),
    .io_pipe_phv_out_data_442(mau_7_io_pipe_phv_out_data_442),
    .io_pipe_phv_out_data_443(mau_7_io_pipe_phv_out_data_443),
    .io_pipe_phv_out_data_444(mau_7_io_pipe_phv_out_data_444),
    .io_pipe_phv_out_data_445(mau_7_io_pipe_phv_out_data_445),
    .io_pipe_phv_out_data_446(mau_7_io_pipe_phv_out_data_446),
    .io_pipe_phv_out_data_447(mau_7_io_pipe_phv_out_data_447),
    .io_pipe_phv_out_data_448(mau_7_io_pipe_phv_out_data_448),
    .io_pipe_phv_out_data_449(mau_7_io_pipe_phv_out_data_449),
    .io_pipe_phv_out_data_450(mau_7_io_pipe_phv_out_data_450),
    .io_pipe_phv_out_data_451(mau_7_io_pipe_phv_out_data_451),
    .io_pipe_phv_out_data_452(mau_7_io_pipe_phv_out_data_452),
    .io_pipe_phv_out_data_453(mau_7_io_pipe_phv_out_data_453),
    .io_pipe_phv_out_data_454(mau_7_io_pipe_phv_out_data_454),
    .io_pipe_phv_out_data_455(mau_7_io_pipe_phv_out_data_455),
    .io_pipe_phv_out_data_456(mau_7_io_pipe_phv_out_data_456),
    .io_pipe_phv_out_data_457(mau_7_io_pipe_phv_out_data_457),
    .io_pipe_phv_out_data_458(mau_7_io_pipe_phv_out_data_458),
    .io_pipe_phv_out_data_459(mau_7_io_pipe_phv_out_data_459),
    .io_pipe_phv_out_data_460(mau_7_io_pipe_phv_out_data_460),
    .io_pipe_phv_out_data_461(mau_7_io_pipe_phv_out_data_461),
    .io_pipe_phv_out_data_462(mau_7_io_pipe_phv_out_data_462),
    .io_pipe_phv_out_data_463(mau_7_io_pipe_phv_out_data_463),
    .io_pipe_phv_out_data_464(mau_7_io_pipe_phv_out_data_464),
    .io_pipe_phv_out_data_465(mau_7_io_pipe_phv_out_data_465),
    .io_pipe_phv_out_data_466(mau_7_io_pipe_phv_out_data_466),
    .io_pipe_phv_out_data_467(mau_7_io_pipe_phv_out_data_467),
    .io_pipe_phv_out_data_468(mau_7_io_pipe_phv_out_data_468),
    .io_pipe_phv_out_data_469(mau_7_io_pipe_phv_out_data_469),
    .io_pipe_phv_out_data_470(mau_7_io_pipe_phv_out_data_470),
    .io_pipe_phv_out_data_471(mau_7_io_pipe_phv_out_data_471),
    .io_pipe_phv_out_data_472(mau_7_io_pipe_phv_out_data_472),
    .io_pipe_phv_out_data_473(mau_7_io_pipe_phv_out_data_473),
    .io_pipe_phv_out_data_474(mau_7_io_pipe_phv_out_data_474),
    .io_pipe_phv_out_data_475(mau_7_io_pipe_phv_out_data_475),
    .io_pipe_phv_out_data_476(mau_7_io_pipe_phv_out_data_476),
    .io_pipe_phv_out_data_477(mau_7_io_pipe_phv_out_data_477),
    .io_pipe_phv_out_data_478(mau_7_io_pipe_phv_out_data_478),
    .io_pipe_phv_out_data_479(mau_7_io_pipe_phv_out_data_479),
    .io_pipe_phv_out_data_480(mau_7_io_pipe_phv_out_data_480),
    .io_pipe_phv_out_data_481(mau_7_io_pipe_phv_out_data_481),
    .io_pipe_phv_out_data_482(mau_7_io_pipe_phv_out_data_482),
    .io_pipe_phv_out_data_483(mau_7_io_pipe_phv_out_data_483),
    .io_pipe_phv_out_data_484(mau_7_io_pipe_phv_out_data_484),
    .io_pipe_phv_out_data_485(mau_7_io_pipe_phv_out_data_485),
    .io_pipe_phv_out_data_486(mau_7_io_pipe_phv_out_data_486),
    .io_pipe_phv_out_data_487(mau_7_io_pipe_phv_out_data_487),
    .io_pipe_phv_out_data_488(mau_7_io_pipe_phv_out_data_488),
    .io_pipe_phv_out_data_489(mau_7_io_pipe_phv_out_data_489),
    .io_pipe_phv_out_data_490(mau_7_io_pipe_phv_out_data_490),
    .io_pipe_phv_out_data_491(mau_7_io_pipe_phv_out_data_491),
    .io_pipe_phv_out_data_492(mau_7_io_pipe_phv_out_data_492),
    .io_pipe_phv_out_data_493(mau_7_io_pipe_phv_out_data_493),
    .io_pipe_phv_out_data_494(mau_7_io_pipe_phv_out_data_494),
    .io_pipe_phv_out_data_495(mau_7_io_pipe_phv_out_data_495),
    .io_pipe_phv_out_data_496(mau_7_io_pipe_phv_out_data_496),
    .io_pipe_phv_out_data_497(mau_7_io_pipe_phv_out_data_497),
    .io_pipe_phv_out_data_498(mau_7_io_pipe_phv_out_data_498),
    .io_pipe_phv_out_data_499(mau_7_io_pipe_phv_out_data_499),
    .io_pipe_phv_out_data_500(mau_7_io_pipe_phv_out_data_500),
    .io_pipe_phv_out_data_501(mau_7_io_pipe_phv_out_data_501),
    .io_pipe_phv_out_data_502(mau_7_io_pipe_phv_out_data_502),
    .io_pipe_phv_out_data_503(mau_7_io_pipe_phv_out_data_503),
    .io_pipe_phv_out_data_504(mau_7_io_pipe_phv_out_data_504),
    .io_pipe_phv_out_data_505(mau_7_io_pipe_phv_out_data_505),
    .io_pipe_phv_out_data_506(mau_7_io_pipe_phv_out_data_506),
    .io_pipe_phv_out_data_507(mau_7_io_pipe_phv_out_data_507),
    .io_pipe_phv_out_data_508(mau_7_io_pipe_phv_out_data_508),
    .io_pipe_phv_out_data_509(mau_7_io_pipe_phv_out_data_509),
    .io_pipe_phv_out_data_510(mau_7_io_pipe_phv_out_data_510),
    .io_pipe_phv_out_data_511(mau_7_io_pipe_phv_out_data_511),
    .io_pipe_phv_out_header_0(mau_7_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(mau_7_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(mau_7_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(mau_7_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(mau_7_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(mau_7_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(mau_7_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(mau_7_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(mau_7_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(mau_7_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(mau_7_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(mau_7_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(mau_7_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(mau_7_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(mau_7_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(mau_7_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(mau_7_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(mau_7_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(mau_7_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(mau_7_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(mau_7_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(mau_7_io_pipe_phv_out_is_valid_processor),
    .io_mod_state_id_mod(mau_7_io_mod_state_id_mod),
    .io_mod_state_id(mau_7_io_mod_state_id),
    .io_mod_sram_w_cs(mau_7_io_mod_sram_w_cs),
    .io_mod_sram_w_en(mau_7_io_mod_sram_w_en),
    .io_mod_sram_w_addr(mau_7_io_mod_sram_w_addr),
    .io_mod_sram_w_data(mau_7_io_mod_sram_w_data)
  );
  assign io_pipe_phv_out_data_0 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_0 : _GEN_2692; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_1 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_1 : _GEN_2693; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_2 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_2 : _GEN_2694; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_3 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_3 : _GEN_2695; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_4 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_4 : _GEN_2696; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_5 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_5 : _GEN_2697; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_6 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_6 : _GEN_2698; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_7 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_7 : _GEN_2699; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_8 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_8 : _GEN_2700; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_9 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_9 : _GEN_2701; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_10 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_10 : _GEN_2702; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_11 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_11 : _GEN_2703; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_12 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_12 : _GEN_2704; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_13 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_13 : _GEN_2705; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_14 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_14 : _GEN_2706; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_15 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_15 : _GEN_2707; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_16 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_16 : _GEN_2708; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_17 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_17 : _GEN_2709; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_18 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_18 : _GEN_2710; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_19 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_19 : _GEN_2711; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_20 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_20 : _GEN_2712; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_21 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_21 : _GEN_2713; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_22 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_22 : _GEN_2714; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_23 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_23 : _GEN_2715; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_24 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_24 : _GEN_2716; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_25 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_25 : _GEN_2717; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_26 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_26 : _GEN_2718; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_27 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_27 : _GEN_2719; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_28 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_28 : _GEN_2720; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_29 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_29 : _GEN_2721; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_30 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_30 : _GEN_2722; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_31 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_31 : _GEN_2723; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_32 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_32 : _GEN_2724; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_33 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_33 : _GEN_2725; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_34 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_34 : _GEN_2726; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_35 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_35 : _GEN_2727; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_36 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_36 : _GEN_2728; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_37 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_37 : _GEN_2729; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_38 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_38 : _GEN_2730; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_39 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_39 : _GEN_2731; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_40 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_40 : _GEN_2732; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_41 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_41 : _GEN_2733; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_42 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_42 : _GEN_2734; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_43 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_43 : _GEN_2735; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_44 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_44 : _GEN_2736; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_45 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_45 : _GEN_2737; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_46 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_46 : _GEN_2738; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_47 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_47 : _GEN_2739; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_48 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_48 : _GEN_2740; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_49 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_49 : _GEN_2741; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_50 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_50 : _GEN_2742; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_51 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_51 : _GEN_2743; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_52 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_52 : _GEN_2744; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_53 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_53 : _GEN_2745; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_54 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_54 : _GEN_2746; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_55 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_55 : _GEN_2747; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_56 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_56 : _GEN_2748; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_57 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_57 : _GEN_2749; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_58 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_58 : _GEN_2750; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_59 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_59 : _GEN_2751; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_60 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_60 : _GEN_2752; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_61 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_61 : _GEN_2753; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_62 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_62 : _GEN_2754; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_63 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_63 : _GEN_2755; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_64 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_64 : _GEN_2756; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_65 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_65 : _GEN_2757; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_66 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_66 : _GEN_2758; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_67 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_67 : _GEN_2759; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_68 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_68 : _GEN_2760; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_69 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_69 : _GEN_2761; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_70 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_70 : _GEN_2762; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_71 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_71 : _GEN_2763; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_72 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_72 : _GEN_2764; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_73 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_73 : _GEN_2765; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_74 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_74 : _GEN_2766; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_75 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_75 : _GEN_2767; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_76 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_76 : _GEN_2768; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_77 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_77 : _GEN_2769; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_78 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_78 : _GEN_2770; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_79 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_79 : _GEN_2771; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_80 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_80 : _GEN_2772; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_81 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_81 : _GEN_2773; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_82 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_82 : _GEN_2774; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_83 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_83 : _GEN_2775; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_84 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_84 : _GEN_2776; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_85 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_85 : _GEN_2777; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_86 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_86 : _GEN_2778; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_87 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_87 : _GEN_2779; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_88 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_88 : _GEN_2780; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_89 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_89 : _GEN_2781; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_90 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_90 : _GEN_2782; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_91 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_91 : _GEN_2783; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_92 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_92 : _GEN_2784; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_93 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_93 : _GEN_2785; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_94 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_94 : _GEN_2786; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_95 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_95 : _GEN_2787; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_96 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_96 : _GEN_2788; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_97 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_97 : _GEN_2789; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_98 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_98 : _GEN_2790; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_99 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_99 : _GEN_2791; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_100 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_100 : _GEN_2792; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_101 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_101 : _GEN_2793; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_102 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_102 : _GEN_2794; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_103 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_103 : _GEN_2795; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_104 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_104 : _GEN_2796; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_105 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_105 : _GEN_2797; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_106 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_106 : _GEN_2798; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_107 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_107 : _GEN_2799; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_108 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_108 : _GEN_2800; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_109 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_109 : _GEN_2801; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_110 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_110 : _GEN_2802; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_111 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_111 : _GEN_2803; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_112 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_112 : _GEN_2804; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_113 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_113 : _GEN_2805; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_114 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_114 : _GEN_2806; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_115 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_115 : _GEN_2807; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_116 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_116 : _GEN_2808; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_117 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_117 : _GEN_2809; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_118 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_118 : _GEN_2810; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_119 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_119 : _GEN_2811; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_120 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_120 : _GEN_2812; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_121 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_121 : _GEN_2813; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_122 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_122 : _GEN_2814; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_123 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_123 : _GEN_2815; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_124 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_124 : _GEN_2816; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_125 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_125 : _GEN_2817; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_126 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_126 : _GEN_2818; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_127 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_127 : _GEN_2819; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_128 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_128 : _GEN_2820; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_129 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_129 : _GEN_2821; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_130 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_130 : _GEN_2822; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_131 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_131 : _GEN_2823; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_132 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_132 : _GEN_2824; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_133 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_133 : _GEN_2825; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_134 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_134 : _GEN_2826; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_135 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_135 : _GEN_2827; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_136 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_136 : _GEN_2828; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_137 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_137 : _GEN_2829; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_138 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_138 : _GEN_2830; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_139 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_139 : _GEN_2831; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_140 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_140 : _GEN_2832; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_141 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_141 : _GEN_2833; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_142 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_142 : _GEN_2834; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_143 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_143 : _GEN_2835; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_144 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_144 : _GEN_2836; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_145 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_145 : _GEN_2837; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_146 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_146 : _GEN_2838; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_147 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_147 : _GEN_2839; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_148 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_148 : _GEN_2840; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_149 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_149 : _GEN_2841; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_150 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_150 : _GEN_2842; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_151 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_151 : _GEN_2843; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_152 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_152 : _GEN_2844; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_153 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_153 : _GEN_2845; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_154 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_154 : _GEN_2846; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_155 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_155 : _GEN_2847; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_156 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_156 : _GEN_2848; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_157 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_157 : _GEN_2849; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_158 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_158 : _GEN_2850; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_159 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_159 : _GEN_2851; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_160 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_160 : _GEN_2852; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_161 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_161 : _GEN_2853; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_162 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_162 : _GEN_2854; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_163 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_163 : _GEN_2855; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_164 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_164 : _GEN_2856; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_165 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_165 : _GEN_2857; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_166 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_166 : _GEN_2858; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_167 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_167 : _GEN_2859; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_168 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_168 : _GEN_2860; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_169 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_169 : _GEN_2861; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_170 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_170 : _GEN_2862; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_171 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_171 : _GEN_2863; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_172 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_172 : _GEN_2864; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_173 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_173 : _GEN_2865; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_174 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_174 : _GEN_2866; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_175 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_175 : _GEN_2867; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_176 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_176 : _GEN_2868; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_177 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_177 : _GEN_2869; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_178 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_178 : _GEN_2870; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_179 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_179 : _GEN_2871; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_180 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_180 : _GEN_2872; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_181 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_181 : _GEN_2873; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_182 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_182 : _GEN_2874; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_183 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_183 : _GEN_2875; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_184 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_184 : _GEN_2876; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_185 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_185 : _GEN_2877; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_186 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_186 : _GEN_2878; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_187 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_187 : _GEN_2879; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_188 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_188 : _GEN_2880; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_189 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_189 : _GEN_2881; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_190 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_190 : _GEN_2882; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_191 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_191 : _GEN_2883; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_192 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_192 : _GEN_2884; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_193 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_193 : _GEN_2885; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_194 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_194 : _GEN_2886; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_195 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_195 : _GEN_2887; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_196 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_196 : _GEN_2888; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_197 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_197 : _GEN_2889; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_198 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_198 : _GEN_2890; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_199 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_199 : _GEN_2891; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_200 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_200 : _GEN_2892; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_201 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_201 : _GEN_2893; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_202 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_202 : _GEN_2894; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_203 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_203 : _GEN_2895; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_204 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_204 : _GEN_2896; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_205 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_205 : _GEN_2897; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_206 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_206 : _GEN_2898; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_207 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_207 : _GEN_2899; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_208 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_208 : _GEN_2900; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_209 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_209 : _GEN_2901; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_210 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_210 : _GEN_2902; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_211 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_211 : _GEN_2903; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_212 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_212 : _GEN_2904; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_213 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_213 : _GEN_2905; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_214 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_214 : _GEN_2906; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_215 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_215 : _GEN_2907; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_216 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_216 : _GEN_2908; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_217 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_217 : _GEN_2909; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_218 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_218 : _GEN_2910; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_219 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_219 : _GEN_2911; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_220 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_220 : _GEN_2912; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_221 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_221 : _GEN_2913; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_222 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_222 : _GEN_2914; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_223 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_223 : _GEN_2915; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_224 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_224 : _GEN_2916; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_225 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_225 : _GEN_2917; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_226 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_226 : _GEN_2918; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_227 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_227 : _GEN_2919; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_228 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_228 : _GEN_2920; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_229 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_229 : _GEN_2921; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_230 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_230 : _GEN_2922; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_231 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_231 : _GEN_2923; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_232 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_232 : _GEN_2924; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_233 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_233 : _GEN_2925; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_234 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_234 : _GEN_2926; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_235 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_235 : _GEN_2927; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_236 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_236 : _GEN_2928; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_237 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_237 : _GEN_2929; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_238 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_238 : _GEN_2930; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_239 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_239 : _GEN_2931; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_240 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_240 : _GEN_2932; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_241 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_241 : _GEN_2933; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_242 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_242 : _GEN_2934; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_243 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_243 : _GEN_2935; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_244 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_244 : _GEN_2936; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_245 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_245 : _GEN_2937; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_246 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_246 : _GEN_2938; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_247 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_247 : _GEN_2939; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_248 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_248 : _GEN_2940; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_249 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_249 : _GEN_2941; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_250 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_250 : _GEN_2942; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_251 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_251 : _GEN_2943; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_252 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_252 : _GEN_2944; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_253 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_253 : _GEN_2945; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_254 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_254 : _GEN_2946; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_255 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_255 : _GEN_2947; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_256 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_256 : _GEN_2948; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_257 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_257 : _GEN_2949; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_258 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_258 : _GEN_2950; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_259 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_259 : _GEN_2951; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_260 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_260 : _GEN_2952; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_261 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_261 : _GEN_2953; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_262 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_262 : _GEN_2954; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_263 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_263 : _GEN_2955; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_264 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_264 : _GEN_2956; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_265 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_265 : _GEN_2957; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_266 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_266 : _GEN_2958; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_267 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_267 : _GEN_2959; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_268 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_268 : _GEN_2960; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_269 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_269 : _GEN_2961; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_270 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_270 : _GEN_2962; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_271 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_271 : _GEN_2963; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_272 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_272 : _GEN_2964; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_273 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_273 : _GEN_2965; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_274 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_274 : _GEN_2966; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_275 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_275 : _GEN_2967; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_276 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_276 : _GEN_2968; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_277 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_277 : _GEN_2969; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_278 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_278 : _GEN_2970; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_279 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_279 : _GEN_2971; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_280 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_280 : _GEN_2972; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_281 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_281 : _GEN_2973; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_282 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_282 : _GEN_2974; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_283 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_283 : _GEN_2975; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_284 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_284 : _GEN_2976; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_285 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_285 : _GEN_2977; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_286 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_286 : _GEN_2978; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_287 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_287 : _GEN_2979; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_288 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_288 : _GEN_2980; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_289 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_289 : _GEN_2981; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_290 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_290 : _GEN_2982; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_291 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_291 : _GEN_2983; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_292 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_292 : _GEN_2984; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_293 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_293 : _GEN_2985; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_294 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_294 : _GEN_2986; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_295 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_295 : _GEN_2987; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_296 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_296 : _GEN_2988; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_297 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_297 : _GEN_2989; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_298 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_298 : _GEN_2990; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_299 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_299 : _GEN_2991; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_300 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_300 : _GEN_2992; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_301 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_301 : _GEN_2993; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_302 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_302 : _GEN_2994; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_303 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_303 : _GEN_2995; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_304 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_304 : _GEN_2996; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_305 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_305 : _GEN_2997; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_306 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_306 : _GEN_2998; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_307 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_307 : _GEN_2999; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_308 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_308 : _GEN_3000; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_309 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_309 : _GEN_3001; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_310 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_310 : _GEN_3002; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_311 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_311 : _GEN_3003; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_312 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_312 : _GEN_3004; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_313 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_313 : _GEN_3005; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_314 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_314 : _GEN_3006; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_315 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_315 : _GEN_3007; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_316 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_316 : _GEN_3008; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_317 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_317 : _GEN_3009; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_318 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_318 : _GEN_3010; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_319 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_319 : _GEN_3011; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_320 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_320 : _GEN_3012; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_321 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_321 : _GEN_3013; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_322 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_322 : _GEN_3014; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_323 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_323 : _GEN_3015; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_324 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_324 : _GEN_3016; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_325 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_325 : _GEN_3017; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_326 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_326 : _GEN_3018; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_327 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_327 : _GEN_3019; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_328 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_328 : _GEN_3020; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_329 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_329 : _GEN_3021; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_330 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_330 : _GEN_3022; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_331 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_331 : _GEN_3023; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_332 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_332 : _GEN_3024; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_333 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_333 : _GEN_3025; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_334 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_334 : _GEN_3026; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_335 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_335 : _GEN_3027; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_336 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_336 : _GEN_3028; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_337 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_337 : _GEN_3029; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_338 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_338 : _GEN_3030; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_339 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_339 : _GEN_3031; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_340 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_340 : _GEN_3032; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_341 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_341 : _GEN_3033; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_342 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_342 : _GEN_3034; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_343 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_343 : _GEN_3035; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_344 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_344 : _GEN_3036; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_345 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_345 : _GEN_3037; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_346 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_346 : _GEN_3038; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_347 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_347 : _GEN_3039; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_348 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_348 : _GEN_3040; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_349 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_349 : _GEN_3041; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_350 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_350 : _GEN_3042; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_351 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_351 : _GEN_3043; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_352 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_352 : _GEN_3044; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_353 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_353 : _GEN_3045; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_354 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_354 : _GEN_3046; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_355 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_355 : _GEN_3047; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_356 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_356 : _GEN_3048; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_357 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_357 : _GEN_3049; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_358 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_358 : _GEN_3050; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_359 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_359 : _GEN_3051; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_360 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_360 : _GEN_3052; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_361 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_361 : _GEN_3053; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_362 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_362 : _GEN_3054; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_363 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_363 : _GEN_3055; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_364 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_364 : _GEN_3056; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_365 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_365 : _GEN_3057; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_366 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_366 : _GEN_3058; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_367 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_367 : _GEN_3059; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_368 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_368 : _GEN_3060; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_369 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_369 : _GEN_3061; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_370 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_370 : _GEN_3062; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_371 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_371 : _GEN_3063; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_372 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_372 : _GEN_3064; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_373 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_373 : _GEN_3065; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_374 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_374 : _GEN_3066; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_375 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_375 : _GEN_3067; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_376 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_376 : _GEN_3068; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_377 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_377 : _GEN_3069; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_378 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_378 : _GEN_3070; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_379 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_379 : _GEN_3071; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_380 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_380 : _GEN_3072; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_381 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_381 : _GEN_3073; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_382 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_382 : _GEN_3074; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_383 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_383 : _GEN_3075; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_384 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_384 : _GEN_3076; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_385 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_385 : _GEN_3077; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_386 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_386 : _GEN_3078; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_387 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_387 : _GEN_3079; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_388 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_388 : _GEN_3080; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_389 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_389 : _GEN_3081; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_390 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_390 : _GEN_3082; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_391 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_391 : _GEN_3083; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_392 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_392 : _GEN_3084; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_393 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_393 : _GEN_3085; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_394 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_394 : _GEN_3086; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_395 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_395 : _GEN_3087; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_396 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_396 : _GEN_3088; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_397 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_397 : _GEN_3089; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_398 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_398 : _GEN_3090; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_399 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_399 : _GEN_3091; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_400 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_400 : _GEN_3092; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_401 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_401 : _GEN_3093; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_402 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_402 : _GEN_3094; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_403 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_403 : _GEN_3095; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_404 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_404 : _GEN_3096; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_405 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_405 : _GEN_3097; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_406 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_406 : _GEN_3098; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_407 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_407 : _GEN_3099; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_408 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_408 : _GEN_3100; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_409 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_409 : _GEN_3101; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_410 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_410 : _GEN_3102; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_411 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_411 : _GEN_3103; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_412 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_412 : _GEN_3104; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_413 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_413 : _GEN_3105; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_414 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_414 : _GEN_3106; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_415 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_415 : _GEN_3107; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_416 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_416 : _GEN_3108; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_417 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_417 : _GEN_3109; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_418 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_418 : _GEN_3110; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_419 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_419 : _GEN_3111; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_420 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_420 : _GEN_3112; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_421 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_421 : _GEN_3113; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_422 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_422 : _GEN_3114; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_423 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_423 : _GEN_3115; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_424 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_424 : _GEN_3116; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_425 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_425 : _GEN_3117; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_426 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_426 : _GEN_3118; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_427 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_427 : _GEN_3119; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_428 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_428 : _GEN_3120; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_429 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_429 : _GEN_3121; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_430 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_430 : _GEN_3122; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_431 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_431 : _GEN_3123; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_432 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_432 : _GEN_3124; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_433 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_433 : _GEN_3125; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_434 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_434 : _GEN_3126; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_435 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_435 : _GEN_3127; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_436 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_436 : _GEN_3128; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_437 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_437 : _GEN_3129; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_438 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_438 : _GEN_3130; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_439 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_439 : _GEN_3131; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_440 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_440 : _GEN_3132; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_441 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_441 : _GEN_3133; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_442 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_442 : _GEN_3134; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_443 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_443 : _GEN_3135; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_444 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_444 : _GEN_3136; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_445 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_445 : _GEN_3137; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_446 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_446 : _GEN_3138; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_447 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_447 : _GEN_3139; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_448 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_448 : _GEN_3140; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_449 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_449 : _GEN_3141; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_450 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_450 : _GEN_3142; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_451 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_451 : _GEN_3143; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_452 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_452 : _GEN_3144; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_453 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_453 : _GEN_3145; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_454 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_454 : _GEN_3146; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_455 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_455 : _GEN_3147; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_456 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_456 : _GEN_3148; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_457 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_457 : _GEN_3149; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_458 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_458 : _GEN_3150; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_459 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_459 : _GEN_3151; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_460 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_460 : _GEN_3152; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_461 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_461 : _GEN_3153; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_462 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_462 : _GEN_3154; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_463 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_463 : _GEN_3155; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_464 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_464 : _GEN_3156; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_465 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_465 : _GEN_3157; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_466 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_466 : _GEN_3158; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_467 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_467 : _GEN_3159; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_468 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_468 : _GEN_3160; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_469 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_469 : _GEN_3161; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_470 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_470 : _GEN_3162; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_471 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_471 : _GEN_3163; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_472 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_472 : _GEN_3164; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_473 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_473 : _GEN_3165; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_474 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_474 : _GEN_3166; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_475 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_475 : _GEN_3167; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_476 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_476 : _GEN_3168; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_477 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_477 : _GEN_3169; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_478 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_478 : _GEN_3170; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_479 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_479 : _GEN_3171; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_480 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_480 : _GEN_3172; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_481 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_481 : _GEN_3173; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_482 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_482 : _GEN_3174; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_483 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_483 : _GEN_3175; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_484 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_484 : _GEN_3176; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_485 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_485 : _GEN_3177; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_486 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_486 : _GEN_3178; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_487 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_487 : _GEN_3179; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_488 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_488 : _GEN_3180; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_489 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_489 : _GEN_3181; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_490 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_490 : _GEN_3182; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_491 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_491 : _GEN_3183; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_492 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_492 : _GEN_3184; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_493 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_493 : _GEN_3185; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_494 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_494 : _GEN_3186; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_495 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_495 : _GEN_3187; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_496 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_496 : _GEN_3188; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_497 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_497 : _GEN_3189; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_498 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_498 : _GEN_3190; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_499 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_499 : _GEN_3191; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_500 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_500 : _GEN_3192; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_501 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_501 : _GEN_3193; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_502 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_502 : _GEN_3194; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_503 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_503 : _GEN_3195; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_504 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_504 : _GEN_3196; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_505 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_505 : _GEN_3197; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_506 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_506 : _GEN_3198; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_507 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_507 : _GEN_3199; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_508 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_508 : _GEN_3200; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_509 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_509 : _GEN_3201; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_510 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_510 : _GEN_3202; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_511 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_511 : _GEN_3203; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_next_processor_id = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_next_processor_id : _GEN_2672; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_next_config_id = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_next_config_id : _GEN_2671; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign mau_0_clock = clock;
  assign mau_0_io_pipe_phv_in_data_0 = io_pipe_phv_in_data_0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_1 = io_pipe_phv_in_data_1; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_2 = io_pipe_phv_in_data_2; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_3 = io_pipe_phv_in_data_3; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_4 = io_pipe_phv_in_data_4; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_5 = io_pipe_phv_in_data_5; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_6 = io_pipe_phv_in_data_6; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_7 = io_pipe_phv_in_data_7; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_8 = io_pipe_phv_in_data_8; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_9 = io_pipe_phv_in_data_9; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_10 = io_pipe_phv_in_data_10; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_11 = io_pipe_phv_in_data_11; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_12 = io_pipe_phv_in_data_12; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_13 = io_pipe_phv_in_data_13; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_14 = io_pipe_phv_in_data_14; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_15 = io_pipe_phv_in_data_15; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_16 = io_pipe_phv_in_data_16; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_17 = io_pipe_phv_in_data_17; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_18 = io_pipe_phv_in_data_18; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_19 = io_pipe_phv_in_data_19; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_20 = io_pipe_phv_in_data_20; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_21 = io_pipe_phv_in_data_21; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_22 = io_pipe_phv_in_data_22; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_23 = io_pipe_phv_in_data_23; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_24 = io_pipe_phv_in_data_24; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_25 = io_pipe_phv_in_data_25; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_26 = io_pipe_phv_in_data_26; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_27 = io_pipe_phv_in_data_27; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_28 = io_pipe_phv_in_data_28; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_29 = io_pipe_phv_in_data_29; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_30 = io_pipe_phv_in_data_30; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_31 = io_pipe_phv_in_data_31; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_32 = io_pipe_phv_in_data_32; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_33 = io_pipe_phv_in_data_33; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_34 = io_pipe_phv_in_data_34; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_35 = io_pipe_phv_in_data_35; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_36 = io_pipe_phv_in_data_36; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_37 = io_pipe_phv_in_data_37; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_38 = io_pipe_phv_in_data_38; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_39 = io_pipe_phv_in_data_39; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_40 = io_pipe_phv_in_data_40; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_41 = io_pipe_phv_in_data_41; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_42 = io_pipe_phv_in_data_42; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_43 = io_pipe_phv_in_data_43; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_44 = io_pipe_phv_in_data_44; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_45 = io_pipe_phv_in_data_45; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_46 = io_pipe_phv_in_data_46; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_47 = io_pipe_phv_in_data_47; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_48 = io_pipe_phv_in_data_48; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_49 = io_pipe_phv_in_data_49; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_50 = io_pipe_phv_in_data_50; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_51 = io_pipe_phv_in_data_51; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_52 = io_pipe_phv_in_data_52; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_53 = io_pipe_phv_in_data_53; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_54 = io_pipe_phv_in_data_54; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_55 = io_pipe_phv_in_data_55; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_56 = io_pipe_phv_in_data_56; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_57 = io_pipe_phv_in_data_57; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_58 = io_pipe_phv_in_data_58; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_59 = io_pipe_phv_in_data_59; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_60 = io_pipe_phv_in_data_60; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_61 = io_pipe_phv_in_data_61; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_62 = io_pipe_phv_in_data_62; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_63 = io_pipe_phv_in_data_63; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_64 = io_pipe_phv_in_data_64; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_65 = io_pipe_phv_in_data_65; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_66 = io_pipe_phv_in_data_66; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_67 = io_pipe_phv_in_data_67; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_68 = io_pipe_phv_in_data_68; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_69 = io_pipe_phv_in_data_69; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_70 = io_pipe_phv_in_data_70; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_71 = io_pipe_phv_in_data_71; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_72 = io_pipe_phv_in_data_72; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_73 = io_pipe_phv_in_data_73; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_74 = io_pipe_phv_in_data_74; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_75 = io_pipe_phv_in_data_75; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_76 = io_pipe_phv_in_data_76; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_77 = io_pipe_phv_in_data_77; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_78 = io_pipe_phv_in_data_78; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_79 = io_pipe_phv_in_data_79; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_80 = io_pipe_phv_in_data_80; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_81 = io_pipe_phv_in_data_81; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_82 = io_pipe_phv_in_data_82; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_83 = io_pipe_phv_in_data_83; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_84 = io_pipe_phv_in_data_84; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_85 = io_pipe_phv_in_data_85; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_86 = io_pipe_phv_in_data_86; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_87 = io_pipe_phv_in_data_87; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_88 = io_pipe_phv_in_data_88; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_89 = io_pipe_phv_in_data_89; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_90 = io_pipe_phv_in_data_90; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_91 = io_pipe_phv_in_data_91; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_92 = io_pipe_phv_in_data_92; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_93 = io_pipe_phv_in_data_93; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_94 = io_pipe_phv_in_data_94; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_95 = io_pipe_phv_in_data_95; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_96 = io_pipe_phv_in_data_96; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_97 = io_pipe_phv_in_data_97; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_98 = io_pipe_phv_in_data_98; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_99 = io_pipe_phv_in_data_99; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_100 = io_pipe_phv_in_data_100; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_101 = io_pipe_phv_in_data_101; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_102 = io_pipe_phv_in_data_102; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_103 = io_pipe_phv_in_data_103; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_104 = io_pipe_phv_in_data_104; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_105 = io_pipe_phv_in_data_105; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_106 = io_pipe_phv_in_data_106; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_107 = io_pipe_phv_in_data_107; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_108 = io_pipe_phv_in_data_108; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_109 = io_pipe_phv_in_data_109; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_110 = io_pipe_phv_in_data_110; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_111 = io_pipe_phv_in_data_111; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_112 = io_pipe_phv_in_data_112; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_113 = io_pipe_phv_in_data_113; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_114 = io_pipe_phv_in_data_114; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_115 = io_pipe_phv_in_data_115; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_116 = io_pipe_phv_in_data_116; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_117 = io_pipe_phv_in_data_117; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_118 = io_pipe_phv_in_data_118; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_119 = io_pipe_phv_in_data_119; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_120 = io_pipe_phv_in_data_120; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_121 = io_pipe_phv_in_data_121; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_122 = io_pipe_phv_in_data_122; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_123 = io_pipe_phv_in_data_123; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_124 = io_pipe_phv_in_data_124; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_125 = io_pipe_phv_in_data_125; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_126 = io_pipe_phv_in_data_126; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_127 = io_pipe_phv_in_data_127; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_128 = io_pipe_phv_in_data_128; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_129 = io_pipe_phv_in_data_129; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_130 = io_pipe_phv_in_data_130; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_131 = io_pipe_phv_in_data_131; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_132 = io_pipe_phv_in_data_132; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_133 = io_pipe_phv_in_data_133; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_134 = io_pipe_phv_in_data_134; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_135 = io_pipe_phv_in_data_135; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_136 = io_pipe_phv_in_data_136; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_137 = io_pipe_phv_in_data_137; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_138 = io_pipe_phv_in_data_138; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_139 = io_pipe_phv_in_data_139; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_140 = io_pipe_phv_in_data_140; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_141 = io_pipe_phv_in_data_141; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_142 = io_pipe_phv_in_data_142; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_143 = io_pipe_phv_in_data_143; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_144 = io_pipe_phv_in_data_144; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_145 = io_pipe_phv_in_data_145; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_146 = io_pipe_phv_in_data_146; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_147 = io_pipe_phv_in_data_147; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_148 = io_pipe_phv_in_data_148; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_149 = io_pipe_phv_in_data_149; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_150 = io_pipe_phv_in_data_150; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_151 = io_pipe_phv_in_data_151; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_152 = io_pipe_phv_in_data_152; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_153 = io_pipe_phv_in_data_153; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_154 = io_pipe_phv_in_data_154; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_155 = io_pipe_phv_in_data_155; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_156 = io_pipe_phv_in_data_156; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_157 = io_pipe_phv_in_data_157; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_158 = io_pipe_phv_in_data_158; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_159 = io_pipe_phv_in_data_159; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_160 = io_pipe_phv_in_data_160; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_161 = io_pipe_phv_in_data_161; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_162 = io_pipe_phv_in_data_162; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_163 = io_pipe_phv_in_data_163; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_164 = io_pipe_phv_in_data_164; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_165 = io_pipe_phv_in_data_165; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_166 = io_pipe_phv_in_data_166; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_167 = io_pipe_phv_in_data_167; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_168 = io_pipe_phv_in_data_168; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_169 = io_pipe_phv_in_data_169; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_170 = io_pipe_phv_in_data_170; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_171 = io_pipe_phv_in_data_171; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_172 = io_pipe_phv_in_data_172; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_173 = io_pipe_phv_in_data_173; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_174 = io_pipe_phv_in_data_174; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_175 = io_pipe_phv_in_data_175; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_176 = io_pipe_phv_in_data_176; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_177 = io_pipe_phv_in_data_177; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_178 = io_pipe_phv_in_data_178; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_179 = io_pipe_phv_in_data_179; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_180 = io_pipe_phv_in_data_180; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_181 = io_pipe_phv_in_data_181; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_182 = io_pipe_phv_in_data_182; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_183 = io_pipe_phv_in_data_183; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_184 = io_pipe_phv_in_data_184; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_185 = io_pipe_phv_in_data_185; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_186 = io_pipe_phv_in_data_186; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_187 = io_pipe_phv_in_data_187; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_188 = io_pipe_phv_in_data_188; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_189 = io_pipe_phv_in_data_189; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_190 = io_pipe_phv_in_data_190; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_191 = io_pipe_phv_in_data_191; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_192 = io_pipe_phv_in_data_192; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_193 = io_pipe_phv_in_data_193; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_194 = io_pipe_phv_in_data_194; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_195 = io_pipe_phv_in_data_195; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_196 = io_pipe_phv_in_data_196; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_197 = io_pipe_phv_in_data_197; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_198 = io_pipe_phv_in_data_198; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_199 = io_pipe_phv_in_data_199; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_200 = io_pipe_phv_in_data_200; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_201 = io_pipe_phv_in_data_201; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_202 = io_pipe_phv_in_data_202; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_203 = io_pipe_phv_in_data_203; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_204 = io_pipe_phv_in_data_204; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_205 = io_pipe_phv_in_data_205; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_206 = io_pipe_phv_in_data_206; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_207 = io_pipe_phv_in_data_207; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_208 = io_pipe_phv_in_data_208; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_209 = io_pipe_phv_in_data_209; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_210 = io_pipe_phv_in_data_210; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_211 = io_pipe_phv_in_data_211; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_212 = io_pipe_phv_in_data_212; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_213 = io_pipe_phv_in_data_213; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_214 = io_pipe_phv_in_data_214; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_215 = io_pipe_phv_in_data_215; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_216 = io_pipe_phv_in_data_216; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_217 = io_pipe_phv_in_data_217; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_218 = io_pipe_phv_in_data_218; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_219 = io_pipe_phv_in_data_219; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_220 = io_pipe_phv_in_data_220; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_221 = io_pipe_phv_in_data_221; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_222 = io_pipe_phv_in_data_222; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_223 = io_pipe_phv_in_data_223; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_224 = io_pipe_phv_in_data_224; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_225 = io_pipe_phv_in_data_225; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_226 = io_pipe_phv_in_data_226; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_227 = io_pipe_phv_in_data_227; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_228 = io_pipe_phv_in_data_228; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_229 = io_pipe_phv_in_data_229; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_230 = io_pipe_phv_in_data_230; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_231 = io_pipe_phv_in_data_231; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_232 = io_pipe_phv_in_data_232; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_233 = io_pipe_phv_in_data_233; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_234 = io_pipe_phv_in_data_234; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_235 = io_pipe_phv_in_data_235; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_236 = io_pipe_phv_in_data_236; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_237 = io_pipe_phv_in_data_237; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_238 = io_pipe_phv_in_data_238; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_239 = io_pipe_phv_in_data_239; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_240 = io_pipe_phv_in_data_240; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_241 = io_pipe_phv_in_data_241; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_242 = io_pipe_phv_in_data_242; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_243 = io_pipe_phv_in_data_243; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_244 = io_pipe_phv_in_data_244; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_245 = io_pipe_phv_in_data_245; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_246 = io_pipe_phv_in_data_246; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_247 = io_pipe_phv_in_data_247; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_248 = io_pipe_phv_in_data_248; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_249 = io_pipe_phv_in_data_249; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_250 = io_pipe_phv_in_data_250; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_251 = io_pipe_phv_in_data_251; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_252 = io_pipe_phv_in_data_252; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_253 = io_pipe_phv_in_data_253; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_254 = io_pipe_phv_in_data_254; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_255 = io_pipe_phv_in_data_255; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_256 = io_pipe_phv_in_data_256; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_257 = io_pipe_phv_in_data_257; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_258 = io_pipe_phv_in_data_258; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_259 = io_pipe_phv_in_data_259; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_260 = io_pipe_phv_in_data_260; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_261 = io_pipe_phv_in_data_261; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_262 = io_pipe_phv_in_data_262; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_263 = io_pipe_phv_in_data_263; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_264 = io_pipe_phv_in_data_264; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_265 = io_pipe_phv_in_data_265; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_266 = io_pipe_phv_in_data_266; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_267 = io_pipe_phv_in_data_267; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_268 = io_pipe_phv_in_data_268; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_269 = io_pipe_phv_in_data_269; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_270 = io_pipe_phv_in_data_270; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_271 = io_pipe_phv_in_data_271; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_272 = io_pipe_phv_in_data_272; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_273 = io_pipe_phv_in_data_273; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_274 = io_pipe_phv_in_data_274; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_275 = io_pipe_phv_in_data_275; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_276 = io_pipe_phv_in_data_276; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_277 = io_pipe_phv_in_data_277; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_278 = io_pipe_phv_in_data_278; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_279 = io_pipe_phv_in_data_279; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_280 = io_pipe_phv_in_data_280; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_281 = io_pipe_phv_in_data_281; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_282 = io_pipe_phv_in_data_282; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_283 = io_pipe_phv_in_data_283; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_284 = io_pipe_phv_in_data_284; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_285 = io_pipe_phv_in_data_285; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_286 = io_pipe_phv_in_data_286; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_287 = io_pipe_phv_in_data_287; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_288 = io_pipe_phv_in_data_288; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_289 = io_pipe_phv_in_data_289; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_290 = io_pipe_phv_in_data_290; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_291 = io_pipe_phv_in_data_291; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_292 = io_pipe_phv_in_data_292; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_293 = io_pipe_phv_in_data_293; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_294 = io_pipe_phv_in_data_294; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_295 = io_pipe_phv_in_data_295; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_296 = io_pipe_phv_in_data_296; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_297 = io_pipe_phv_in_data_297; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_298 = io_pipe_phv_in_data_298; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_299 = io_pipe_phv_in_data_299; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_300 = io_pipe_phv_in_data_300; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_301 = io_pipe_phv_in_data_301; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_302 = io_pipe_phv_in_data_302; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_303 = io_pipe_phv_in_data_303; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_304 = io_pipe_phv_in_data_304; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_305 = io_pipe_phv_in_data_305; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_306 = io_pipe_phv_in_data_306; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_307 = io_pipe_phv_in_data_307; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_308 = io_pipe_phv_in_data_308; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_309 = io_pipe_phv_in_data_309; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_310 = io_pipe_phv_in_data_310; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_311 = io_pipe_phv_in_data_311; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_312 = io_pipe_phv_in_data_312; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_313 = io_pipe_phv_in_data_313; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_314 = io_pipe_phv_in_data_314; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_315 = io_pipe_phv_in_data_315; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_316 = io_pipe_phv_in_data_316; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_317 = io_pipe_phv_in_data_317; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_318 = io_pipe_phv_in_data_318; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_319 = io_pipe_phv_in_data_319; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_320 = io_pipe_phv_in_data_320; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_321 = io_pipe_phv_in_data_321; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_322 = io_pipe_phv_in_data_322; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_323 = io_pipe_phv_in_data_323; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_324 = io_pipe_phv_in_data_324; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_325 = io_pipe_phv_in_data_325; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_326 = io_pipe_phv_in_data_326; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_327 = io_pipe_phv_in_data_327; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_328 = io_pipe_phv_in_data_328; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_329 = io_pipe_phv_in_data_329; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_330 = io_pipe_phv_in_data_330; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_331 = io_pipe_phv_in_data_331; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_332 = io_pipe_phv_in_data_332; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_333 = io_pipe_phv_in_data_333; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_334 = io_pipe_phv_in_data_334; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_335 = io_pipe_phv_in_data_335; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_336 = io_pipe_phv_in_data_336; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_337 = io_pipe_phv_in_data_337; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_338 = io_pipe_phv_in_data_338; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_339 = io_pipe_phv_in_data_339; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_340 = io_pipe_phv_in_data_340; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_341 = io_pipe_phv_in_data_341; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_342 = io_pipe_phv_in_data_342; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_343 = io_pipe_phv_in_data_343; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_344 = io_pipe_phv_in_data_344; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_345 = io_pipe_phv_in_data_345; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_346 = io_pipe_phv_in_data_346; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_347 = io_pipe_phv_in_data_347; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_348 = io_pipe_phv_in_data_348; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_349 = io_pipe_phv_in_data_349; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_350 = io_pipe_phv_in_data_350; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_351 = io_pipe_phv_in_data_351; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_352 = io_pipe_phv_in_data_352; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_353 = io_pipe_phv_in_data_353; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_354 = io_pipe_phv_in_data_354; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_355 = io_pipe_phv_in_data_355; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_356 = io_pipe_phv_in_data_356; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_357 = io_pipe_phv_in_data_357; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_358 = io_pipe_phv_in_data_358; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_359 = io_pipe_phv_in_data_359; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_360 = io_pipe_phv_in_data_360; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_361 = io_pipe_phv_in_data_361; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_362 = io_pipe_phv_in_data_362; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_363 = io_pipe_phv_in_data_363; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_364 = io_pipe_phv_in_data_364; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_365 = io_pipe_phv_in_data_365; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_366 = io_pipe_phv_in_data_366; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_367 = io_pipe_phv_in_data_367; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_368 = io_pipe_phv_in_data_368; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_369 = io_pipe_phv_in_data_369; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_370 = io_pipe_phv_in_data_370; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_371 = io_pipe_phv_in_data_371; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_372 = io_pipe_phv_in_data_372; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_373 = io_pipe_phv_in_data_373; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_374 = io_pipe_phv_in_data_374; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_375 = io_pipe_phv_in_data_375; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_376 = io_pipe_phv_in_data_376; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_377 = io_pipe_phv_in_data_377; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_378 = io_pipe_phv_in_data_378; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_379 = io_pipe_phv_in_data_379; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_380 = io_pipe_phv_in_data_380; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_381 = io_pipe_phv_in_data_381; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_382 = io_pipe_phv_in_data_382; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_383 = io_pipe_phv_in_data_383; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_384 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_385 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_386 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_387 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_388 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_389 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_390 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_391 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_392 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_393 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_394 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_395 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_396 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_397 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_398 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_399 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_400 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_401 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_402 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_403 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_404 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_405 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_406 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_407 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_408 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_409 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_410 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_411 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_412 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_413 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_414 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_415 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_416 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_417 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_418 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_419 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_420 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_421 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_422 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_423 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_424 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_425 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_426 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_427 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_428 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_429 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_430 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_431 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_432 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_433 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_434 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_435 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_436 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_437 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_438 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_439 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_440 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_441 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_442 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_443 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_444 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_445 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_446 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_447 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_448 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_449 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_450 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_451 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_452 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_453 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_454 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_455 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_456 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_457 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_458 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_459 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_460 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_461 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_462 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_463 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_464 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_465 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_466 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_467 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_468 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_469 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_470 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_471 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_472 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_473 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_474 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_475 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_476 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_477 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_478 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_479 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_480 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_481 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_482 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_483 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_484 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_485 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_486 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_487 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_488 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_489 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_490 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_491 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_492 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_493 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_494 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_495 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_496 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_497 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_498 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_499 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_500 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_501 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_502 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_503 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_504 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_505 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_506 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_507 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_508 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_509 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_510 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_511 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_header_0 = 16'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_header_1 = 16'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_header_2 = 16'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_header_3 = 16'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_header_4 = 16'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_header_5 = 16'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_header_6 = 16'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_header_7 = 16'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_header_8 = 16'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_header_9 = 16'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_header_10 = 16'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_header_11 = 16'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_header_12 = 16'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_header_13 = 16'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_header_14 = 16'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_header_15 = 16'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_parse_current_state = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_parse_current_offset = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_parse_transition_field = 16'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_next_processor_id = 4'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_next_config_id = 1'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_is_valid_processor = 1'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_mod_state_id_mod = io_mod_en ? io_mod_module_mod_state_id_mod & mod_j : io_mod_module_mod_state_id_mod
    ; // @[parser_pisa.scala 51:22 parser_pisa.scala 58:40 parser_pisa.scala 47:23]
  assign mau_0_io_mod_state_id = io_mod_module_mod_state_id; // @[parser_pisa.scala 47:23]
  assign mau_0_io_mod_sram_w_cs = io_mod_module_mod_sram_w_cs; // @[parser_pisa.scala 47:23]
  assign mau_0_io_mod_sram_w_en = io_mod_en ? io_mod_module_mod_sram_w_en & mod_j : io_mod_module_mod_sram_w_en; // @[parser_pisa.scala 51:22 parser_pisa.scala 57:40 parser_pisa.scala 47:23]
  assign mau_0_io_mod_sram_w_addr = io_mod_module_mod_sram_w_addr; // @[parser_pisa.scala 47:23]
  assign mau_0_io_mod_sram_w_data = io_mod_module_mod_sram_w_data; // @[parser_pisa.scala 47:23]
  assign mau_1_clock = clock;
  assign mau_1_io_pipe_phv_in_data_0 = mau_0_io_pipe_phv_out_data_0; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_1 = mau_0_io_pipe_phv_out_data_1; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_2 = mau_0_io_pipe_phv_out_data_2; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_3 = mau_0_io_pipe_phv_out_data_3; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_4 = mau_0_io_pipe_phv_out_data_4; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_5 = mau_0_io_pipe_phv_out_data_5; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_6 = mau_0_io_pipe_phv_out_data_6; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_7 = mau_0_io_pipe_phv_out_data_7; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_8 = mau_0_io_pipe_phv_out_data_8; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_9 = mau_0_io_pipe_phv_out_data_9; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_10 = mau_0_io_pipe_phv_out_data_10; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_11 = mau_0_io_pipe_phv_out_data_11; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_12 = mau_0_io_pipe_phv_out_data_12; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_13 = mau_0_io_pipe_phv_out_data_13; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_14 = mau_0_io_pipe_phv_out_data_14; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_15 = mau_0_io_pipe_phv_out_data_15; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_16 = mau_0_io_pipe_phv_out_data_16; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_17 = mau_0_io_pipe_phv_out_data_17; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_18 = mau_0_io_pipe_phv_out_data_18; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_19 = mau_0_io_pipe_phv_out_data_19; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_20 = mau_0_io_pipe_phv_out_data_20; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_21 = mau_0_io_pipe_phv_out_data_21; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_22 = mau_0_io_pipe_phv_out_data_22; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_23 = mau_0_io_pipe_phv_out_data_23; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_24 = mau_0_io_pipe_phv_out_data_24; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_25 = mau_0_io_pipe_phv_out_data_25; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_26 = mau_0_io_pipe_phv_out_data_26; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_27 = mau_0_io_pipe_phv_out_data_27; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_28 = mau_0_io_pipe_phv_out_data_28; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_29 = mau_0_io_pipe_phv_out_data_29; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_30 = mau_0_io_pipe_phv_out_data_30; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_31 = mau_0_io_pipe_phv_out_data_31; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_32 = mau_0_io_pipe_phv_out_data_32; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_33 = mau_0_io_pipe_phv_out_data_33; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_34 = mau_0_io_pipe_phv_out_data_34; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_35 = mau_0_io_pipe_phv_out_data_35; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_36 = mau_0_io_pipe_phv_out_data_36; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_37 = mau_0_io_pipe_phv_out_data_37; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_38 = mau_0_io_pipe_phv_out_data_38; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_39 = mau_0_io_pipe_phv_out_data_39; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_40 = mau_0_io_pipe_phv_out_data_40; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_41 = mau_0_io_pipe_phv_out_data_41; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_42 = mau_0_io_pipe_phv_out_data_42; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_43 = mau_0_io_pipe_phv_out_data_43; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_44 = mau_0_io_pipe_phv_out_data_44; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_45 = mau_0_io_pipe_phv_out_data_45; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_46 = mau_0_io_pipe_phv_out_data_46; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_47 = mau_0_io_pipe_phv_out_data_47; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_48 = mau_0_io_pipe_phv_out_data_48; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_49 = mau_0_io_pipe_phv_out_data_49; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_50 = mau_0_io_pipe_phv_out_data_50; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_51 = mau_0_io_pipe_phv_out_data_51; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_52 = mau_0_io_pipe_phv_out_data_52; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_53 = mau_0_io_pipe_phv_out_data_53; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_54 = mau_0_io_pipe_phv_out_data_54; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_55 = mau_0_io_pipe_phv_out_data_55; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_56 = mau_0_io_pipe_phv_out_data_56; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_57 = mau_0_io_pipe_phv_out_data_57; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_58 = mau_0_io_pipe_phv_out_data_58; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_59 = mau_0_io_pipe_phv_out_data_59; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_60 = mau_0_io_pipe_phv_out_data_60; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_61 = mau_0_io_pipe_phv_out_data_61; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_62 = mau_0_io_pipe_phv_out_data_62; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_63 = mau_0_io_pipe_phv_out_data_63; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_64 = mau_0_io_pipe_phv_out_data_64; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_65 = mau_0_io_pipe_phv_out_data_65; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_66 = mau_0_io_pipe_phv_out_data_66; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_67 = mau_0_io_pipe_phv_out_data_67; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_68 = mau_0_io_pipe_phv_out_data_68; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_69 = mau_0_io_pipe_phv_out_data_69; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_70 = mau_0_io_pipe_phv_out_data_70; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_71 = mau_0_io_pipe_phv_out_data_71; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_72 = mau_0_io_pipe_phv_out_data_72; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_73 = mau_0_io_pipe_phv_out_data_73; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_74 = mau_0_io_pipe_phv_out_data_74; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_75 = mau_0_io_pipe_phv_out_data_75; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_76 = mau_0_io_pipe_phv_out_data_76; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_77 = mau_0_io_pipe_phv_out_data_77; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_78 = mau_0_io_pipe_phv_out_data_78; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_79 = mau_0_io_pipe_phv_out_data_79; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_80 = mau_0_io_pipe_phv_out_data_80; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_81 = mau_0_io_pipe_phv_out_data_81; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_82 = mau_0_io_pipe_phv_out_data_82; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_83 = mau_0_io_pipe_phv_out_data_83; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_84 = mau_0_io_pipe_phv_out_data_84; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_85 = mau_0_io_pipe_phv_out_data_85; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_86 = mau_0_io_pipe_phv_out_data_86; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_87 = mau_0_io_pipe_phv_out_data_87; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_88 = mau_0_io_pipe_phv_out_data_88; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_89 = mau_0_io_pipe_phv_out_data_89; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_90 = mau_0_io_pipe_phv_out_data_90; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_91 = mau_0_io_pipe_phv_out_data_91; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_92 = mau_0_io_pipe_phv_out_data_92; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_93 = mau_0_io_pipe_phv_out_data_93; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_94 = mau_0_io_pipe_phv_out_data_94; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_95 = mau_0_io_pipe_phv_out_data_95; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_96 = mau_0_io_pipe_phv_out_data_96; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_97 = mau_0_io_pipe_phv_out_data_97; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_98 = mau_0_io_pipe_phv_out_data_98; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_99 = mau_0_io_pipe_phv_out_data_99; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_100 = mau_0_io_pipe_phv_out_data_100; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_101 = mau_0_io_pipe_phv_out_data_101; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_102 = mau_0_io_pipe_phv_out_data_102; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_103 = mau_0_io_pipe_phv_out_data_103; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_104 = mau_0_io_pipe_phv_out_data_104; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_105 = mau_0_io_pipe_phv_out_data_105; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_106 = mau_0_io_pipe_phv_out_data_106; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_107 = mau_0_io_pipe_phv_out_data_107; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_108 = mau_0_io_pipe_phv_out_data_108; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_109 = mau_0_io_pipe_phv_out_data_109; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_110 = mau_0_io_pipe_phv_out_data_110; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_111 = mau_0_io_pipe_phv_out_data_111; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_112 = mau_0_io_pipe_phv_out_data_112; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_113 = mau_0_io_pipe_phv_out_data_113; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_114 = mau_0_io_pipe_phv_out_data_114; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_115 = mau_0_io_pipe_phv_out_data_115; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_116 = mau_0_io_pipe_phv_out_data_116; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_117 = mau_0_io_pipe_phv_out_data_117; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_118 = mau_0_io_pipe_phv_out_data_118; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_119 = mau_0_io_pipe_phv_out_data_119; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_120 = mau_0_io_pipe_phv_out_data_120; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_121 = mau_0_io_pipe_phv_out_data_121; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_122 = mau_0_io_pipe_phv_out_data_122; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_123 = mau_0_io_pipe_phv_out_data_123; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_124 = mau_0_io_pipe_phv_out_data_124; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_125 = mau_0_io_pipe_phv_out_data_125; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_126 = mau_0_io_pipe_phv_out_data_126; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_127 = mau_0_io_pipe_phv_out_data_127; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_128 = mau_0_io_pipe_phv_out_data_128; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_129 = mau_0_io_pipe_phv_out_data_129; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_130 = mau_0_io_pipe_phv_out_data_130; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_131 = mau_0_io_pipe_phv_out_data_131; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_132 = mau_0_io_pipe_phv_out_data_132; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_133 = mau_0_io_pipe_phv_out_data_133; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_134 = mau_0_io_pipe_phv_out_data_134; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_135 = mau_0_io_pipe_phv_out_data_135; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_136 = mau_0_io_pipe_phv_out_data_136; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_137 = mau_0_io_pipe_phv_out_data_137; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_138 = mau_0_io_pipe_phv_out_data_138; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_139 = mau_0_io_pipe_phv_out_data_139; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_140 = mau_0_io_pipe_phv_out_data_140; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_141 = mau_0_io_pipe_phv_out_data_141; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_142 = mau_0_io_pipe_phv_out_data_142; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_143 = mau_0_io_pipe_phv_out_data_143; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_144 = mau_0_io_pipe_phv_out_data_144; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_145 = mau_0_io_pipe_phv_out_data_145; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_146 = mau_0_io_pipe_phv_out_data_146; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_147 = mau_0_io_pipe_phv_out_data_147; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_148 = mau_0_io_pipe_phv_out_data_148; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_149 = mau_0_io_pipe_phv_out_data_149; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_150 = mau_0_io_pipe_phv_out_data_150; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_151 = mau_0_io_pipe_phv_out_data_151; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_152 = mau_0_io_pipe_phv_out_data_152; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_153 = mau_0_io_pipe_phv_out_data_153; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_154 = mau_0_io_pipe_phv_out_data_154; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_155 = mau_0_io_pipe_phv_out_data_155; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_156 = mau_0_io_pipe_phv_out_data_156; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_157 = mau_0_io_pipe_phv_out_data_157; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_158 = mau_0_io_pipe_phv_out_data_158; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_159 = mau_0_io_pipe_phv_out_data_159; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_160 = mau_0_io_pipe_phv_out_data_160; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_161 = mau_0_io_pipe_phv_out_data_161; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_162 = mau_0_io_pipe_phv_out_data_162; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_163 = mau_0_io_pipe_phv_out_data_163; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_164 = mau_0_io_pipe_phv_out_data_164; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_165 = mau_0_io_pipe_phv_out_data_165; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_166 = mau_0_io_pipe_phv_out_data_166; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_167 = mau_0_io_pipe_phv_out_data_167; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_168 = mau_0_io_pipe_phv_out_data_168; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_169 = mau_0_io_pipe_phv_out_data_169; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_170 = mau_0_io_pipe_phv_out_data_170; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_171 = mau_0_io_pipe_phv_out_data_171; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_172 = mau_0_io_pipe_phv_out_data_172; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_173 = mau_0_io_pipe_phv_out_data_173; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_174 = mau_0_io_pipe_phv_out_data_174; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_175 = mau_0_io_pipe_phv_out_data_175; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_176 = mau_0_io_pipe_phv_out_data_176; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_177 = mau_0_io_pipe_phv_out_data_177; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_178 = mau_0_io_pipe_phv_out_data_178; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_179 = mau_0_io_pipe_phv_out_data_179; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_180 = mau_0_io_pipe_phv_out_data_180; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_181 = mau_0_io_pipe_phv_out_data_181; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_182 = mau_0_io_pipe_phv_out_data_182; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_183 = mau_0_io_pipe_phv_out_data_183; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_184 = mau_0_io_pipe_phv_out_data_184; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_185 = mau_0_io_pipe_phv_out_data_185; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_186 = mau_0_io_pipe_phv_out_data_186; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_187 = mau_0_io_pipe_phv_out_data_187; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_188 = mau_0_io_pipe_phv_out_data_188; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_189 = mau_0_io_pipe_phv_out_data_189; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_190 = mau_0_io_pipe_phv_out_data_190; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_191 = mau_0_io_pipe_phv_out_data_191; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_192 = mau_0_io_pipe_phv_out_data_192; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_193 = mau_0_io_pipe_phv_out_data_193; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_194 = mau_0_io_pipe_phv_out_data_194; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_195 = mau_0_io_pipe_phv_out_data_195; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_196 = mau_0_io_pipe_phv_out_data_196; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_197 = mau_0_io_pipe_phv_out_data_197; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_198 = mau_0_io_pipe_phv_out_data_198; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_199 = mau_0_io_pipe_phv_out_data_199; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_200 = mau_0_io_pipe_phv_out_data_200; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_201 = mau_0_io_pipe_phv_out_data_201; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_202 = mau_0_io_pipe_phv_out_data_202; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_203 = mau_0_io_pipe_phv_out_data_203; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_204 = mau_0_io_pipe_phv_out_data_204; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_205 = mau_0_io_pipe_phv_out_data_205; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_206 = mau_0_io_pipe_phv_out_data_206; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_207 = mau_0_io_pipe_phv_out_data_207; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_208 = mau_0_io_pipe_phv_out_data_208; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_209 = mau_0_io_pipe_phv_out_data_209; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_210 = mau_0_io_pipe_phv_out_data_210; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_211 = mau_0_io_pipe_phv_out_data_211; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_212 = mau_0_io_pipe_phv_out_data_212; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_213 = mau_0_io_pipe_phv_out_data_213; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_214 = mau_0_io_pipe_phv_out_data_214; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_215 = mau_0_io_pipe_phv_out_data_215; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_216 = mau_0_io_pipe_phv_out_data_216; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_217 = mau_0_io_pipe_phv_out_data_217; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_218 = mau_0_io_pipe_phv_out_data_218; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_219 = mau_0_io_pipe_phv_out_data_219; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_220 = mau_0_io_pipe_phv_out_data_220; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_221 = mau_0_io_pipe_phv_out_data_221; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_222 = mau_0_io_pipe_phv_out_data_222; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_223 = mau_0_io_pipe_phv_out_data_223; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_224 = mau_0_io_pipe_phv_out_data_224; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_225 = mau_0_io_pipe_phv_out_data_225; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_226 = mau_0_io_pipe_phv_out_data_226; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_227 = mau_0_io_pipe_phv_out_data_227; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_228 = mau_0_io_pipe_phv_out_data_228; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_229 = mau_0_io_pipe_phv_out_data_229; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_230 = mau_0_io_pipe_phv_out_data_230; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_231 = mau_0_io_pipe_phv_out_data_231; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_232 = mau_0_io_pipe_phv_out_data_232; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_233 = mau_0_io_pipe_phv_out_data_233; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_234 = mau_0_io_pipe_phv_out_data_234; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_235 = mau_0_io_pipe_phv_out_data_235; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_236 = mau_0_io_pipe_phv_out_data_236; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_237 = mau_0_io_pipe_phv_out_data_237; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_238 = mau_0_io_pipe_phv_out_data_238; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_239 = mau_0_io_pipe_phv_out_data_239; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_240 = mau_0_io_pipe_phv_out_data_240; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_241 = mau_0_io_pipe_phv_out_data_241; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_242 = mau_0_io_pipe_phv_out_data_242; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_243 = mau_0_io_pipe_phv_out_data_243; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_244 = mau_0_io_pipe_phv_out_data_244; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_245 = mau_0_io_pipe_phv_out_data_245; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_246 = mau_0_io_pipe_phv_out_data_246; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_247 = mau_0_io_pipe_phv_out_data_247; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_248 = mau_0_io_pipe_phv_out_data_248; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_249 = mau_0_io_pipe_phv_out_data_249; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_250 = mau_0_io_pipe_phv_out_data_250; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_251 = mau_0_io_pipe_phv_out_data_251; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_252 = mau_0_io_pipe_phv_out_data_252; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_253 = mau_0_io_pipe_phv_out_data_253; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_254 = mau_0_io_pipe_phv_out_data_254; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_255 = mau_0_io_pipe_phv_out_data_255; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_256 = mau_0_io_pipe_phv_out_data_256; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_257 = mau_0_io_pipe_phv_out_data_257; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_258 = mau_0_io_pipe_phv_out_data_258; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_259 = mau_0_io_pipe_phv_out_data_259; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_260 = mau_0_io_pipe_phv_out_data_260; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_261 = mau_0_io_pipe_phv_out_data_261; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_262 = mau_0_io_pipe_phv_out_data_262; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_263 = mau_0_io_pipe_phv_out_data_263; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_264 = mau_0_io_pipe_phv_out_data_264; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_265 = mau_0_io_pipe_phv_out_data_265; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_266 = mau_0_io_pipe_phv_out_data_266; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_267 = mau_0_io_pipe_phv_out_data_267; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_268 = mau_0_io_pipe_phv_out_data_268; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_269 = mau_0_io_pipe_phv_out_data_269; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_270 = mau_0_io_pipe_phv_out_data_270; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_271 = mau_0_io_pipe_phv_out_data_271; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_272 = mau_0_io_pipe_phv_out_data_272; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_273 = mau_0_io_pipe_phv_out_data_273; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_274 = mau_0_io_pipe_phv_out_data_274; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_275 = mau_0_io_pipe_phv_out_data_275; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_276 = mau_0_io_pipe_phv_out_data_276; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_277 = mau_0_io_pipe_phv_out_data_277; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_278 = mau_0_io_pipe_phv_out_data_278; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_279 = mau_0_io_pipe_phv_out_data_279; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_280 = mau_0_io_pipe_phv_out_data_280; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_281 = mau_0_io_pipe_phv_out_data_281; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_282 = mau_0_io_pipe_phv_out_data_282; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_283 = mau_0_io_pipe_phv_out_data_283; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_284 = mau_0_io_pipe_phv_out_data_284; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_285 = mau_0_io_pipe_phv_out_data_285; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_286 = mau_0_io_pipe_phv_out_data_286; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_287 = mau_0_io_pipe_phv_out_data_287; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_288 = mau_0_io_pipe_phv_out_data_288; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_289 = mau_0_io_pipe_phv_out_data_289; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_290 = mau_0_io_pipe_phv_out_data_290; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_291 = mau_0_io_pipe_phv_out_data_291; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_292 = mau_0_io_pipe_phv_out_data_292; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_293 = mau_0_io_pipe_phv_out_data_293; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_294 = mau_0_io_pipe_phv_out_data_294; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_295 = mau_0_io_pipe_phv_out_data_295; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_296 = mau_0_io_pipe_phv_out_data_296; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_297 = mau_0_io_pipe_phv_out_data_297; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_298 = mau_0_io_pipe_phv_out_data_298; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_299 = mau_0_io_pipe_phv_out_data_299; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_300 = mau_0_io_pipe_phv_out_data_300; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_301 = mau_0_io_pipe_phv_out_data_301; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_302 = mau_0_io_pipe_phv_out_data_302; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_303 = mau_0_io_pipe_phv_out_data_303; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_304 = mau_0_io_pipe_phv_out_data_304; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_305 = mau_0_io_pipe_phv_out_data_305; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_306 = mau_0_io_pipe_phv_out_data_306; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_307 = mau_0_io_pipe_phv_out_data_307; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_308 = mau_0_io_pipe_phv_out_data_308; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_309 = mau_0_io_pipe_phv_out_data_309; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_310 = mau_0_io_pipe_phv_out_data_310; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_311 = mau_0_io_pipe_phv_out_data_311; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_312 = mau_0_io_pipe_phv_out_data_312; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_313 = mau_0_io_pipe_phv_out_data_313; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_314 = mau_0_io_pipe_phv_out_data_314; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_315 = mau_0_io_pipe_phv_out_data_315; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_316 = mau_0_io_pipe_phv_out_data_316; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_317 = mau_0_io_pipe_phv_out_data_317; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_318 = mau_0_io_pipe_phv_out_data_318; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_319 = mau_0_io_pipe_phv_out_data_319; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_320 = mau_0_io_pipe_phv_out_data_320; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_321 = mau_0_io_pipe_phv_out_data_321; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_322 = mau_0_io_pipe_phv_out_data_322; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_323 = mau_0_io_pipe_phv_out_data_323; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_324 = mau_0_io_pipe_phv_out_data_324; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_325 = mau_0_io_pipe_phv_out_data_325; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_326 = mau_0_io_pipe_phv_out_data_326; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_327 = mau_0_io_pipe_phv_out_data_327; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_328 = mau_0_io_pipe_phv_out_data_328; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_329 = mau_0_io_pipe_phv_out_data_329; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_330 = mau_0_io_pipe_phv_out_data_330; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_331 = mau_0_io_pipe_phv_out_data_331; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_332 = mau_0_io_pipe_phv_out_data_332; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_333 = mau_0_io_pipe_phv_out_data_333; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_334 = mau_0_io_pipe_phv_out_data_334; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_335 = mau_0_io_pipe_phv_out_data_335; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_336 = mau_0_io_pipe_phv_out_data_336; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_337 = mau_0_io_pipe_phv_out_data_337; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_338 = mau_0_io_pipe_phv_out_data_338; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_339 = mau_0_io_pipe_phv_out_data_339; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_340 = mau_0_io_pipe_phv_out_data_340; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_341 = mau_0_io_pipe_phv_out_data_341; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_342 = mau_0_io_pipe_phv_out_data_342; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_343 = mau_0_io_pipe_phv_out_data_343; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_344 = mau_0_io_pipe_phv_out_data_344; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_345 = mau_0_io_pipe_phv_out_data_345; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_346 = mau_0_io_pipe_phv_out_data_346; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_347 = mau_0_io_pipe_phv_out_data_347; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_348 = mau_0_io_pipe_phv_out_data_348; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_349 = mau_0_io_pipe_phv_out_data_349; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_350 = mau_0_io_pipe_phv_out_data_350; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_351 = mau_0_io_pipe_phv_out_data_351; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_352 = mau_0_io_pipe_phv_out_data_352; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_353 = mau_0_io_pipe_phv_out_data_353; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_354 = mau_0_io_pipe_phv_out_data_354; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_355 = mau_0_io_pipe_phv_out_data_355; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_356 = mau_0_io_pipe_phv_out_data_356; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_357 = mau_0_io_pipe_phv_out_data_357; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_358 = mau_0_io_pipe_phv_out_data_358; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_359 = mau_0_io_pipe_phv_out_data_359; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_360 = mau_0_io_pipe_phv_out_data_360; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_361 = mau_0_io_pipe_phv_out_data_361; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_362 = mau_0_io_pipe_phv_out_data_362; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_363 = mau_0_io_pipe_phv_out_data_363; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_364 = mau_0_io_pipe_phv_out_data_364; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_365 = mau_0_io_pipe_phv_out_data_365; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_366 = mau_0_io_pipe_phv_out_data_366; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_367 = mau_0_io_pipe_phv_out_data_367; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_368 = mau_0_io_pipe_phv_out_data_368; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_369 = mau_0_io_pipe_phv_out_data_369; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_370 = mau_0_io_pipe_phv_out_data_370; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_371 = mau_0_io_pipe_phv_out_data_371; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_372 = mau_0_io_pipe_phv_out_data_372; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_373 = mau_0_io_pipe_phv_out_data_373; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_374 = mau_0_io_pipe_phv_out_data_374; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_375 = mau_0_io_pipe_phv_out_data_375; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_376 = mau_0_io_pipe_phv_out_data_376; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_377 = mau_0_io_pipe_phv_out_data_377; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_378 = mau_0_io_pipe_phv_out_data_378; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_379 = mau_0_io_pipe_phv_out_data_379; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_380 = mau_0_io_pipe_phv_out_data_380; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_381 = mau_0_io_pipe_phv_out_data_381; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_382 = mau_0_io_pipe_phv_out_data_382; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_383 = mau_0_io_pipe_phv_out_data_383; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_384 = mau_0_io_pipe_phv_out_data_384; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_385 = mau_0_io_pipe_phv_out_data_385; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_386 = mau_0_io_pipe_phv_out_data_386; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_387 = mau_0_io_pipe_phv_out_data_387; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_388 = mau_0_io_pipe_phv_out_data_388; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_389 = mau_0_io_pipe_phv_out_data_389; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_390 = mau_0_io_pipe_phv_out_data_390; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_391 = mau_0_io_pipe_phv_out_data_391; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_392 = mau_0_io_pipe_phv_out_data_392; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_393 = mau_0_io_pipe_phv_out_data_393; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_394 = mau_0_io_pipe_phv_out_data_394; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_395 = mau_0_io_pipe_phv_out_data_395; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_396 = mau_0_io_pipe_phv_out_data_396; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_397 = mau_0_io_pipe_phv_out_data_397; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_398 = mau_0_io_pipe_phv_out_data_398; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_399 = mau_0_io_pipe_phv_out_data_399; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_400 = mau_0_io_pipe_phv_out_data_400; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_401 = mau_0_io_pipe_phv_out_data_401; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_402 = mau_0_io_pipe_phv_out_data_402; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_403 = mau_0_io_pipe_phv_out_data_403; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_404 = mau_0_io_pipe_phv_out_data_404; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_405 = mau_0_io_pipe_phv_out_data_405; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_406 = mau_0_io_pipe_phv_out_data_406; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_407 = mau_0_io_pipe_phv_out_data_407; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_408 = mau_0_io_pipe_phv_out_data_408; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_409 = mau_0_io_pipe_phv_out_data_409; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_410 = mau_0_io_pipe_phv_out_data_410; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_411 = mau_0_io_pipe_phv_out_data_411; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_412 = mau_0_io_pipe_phv_out_data_412; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_413 = mau_0_io_pipe_phv_out_data_413; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_414 = mau_0_io_pipe_phv_out_data_414; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_415 = mau_0_io_pipe_phv_out_data_415; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_416 = mau_0_io_pipe_phv_out_data_416; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_417 = mau_0_io_pipe_phv_out_data_417; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_418 = mau_0_io_pipe_phv_out_data_418; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_419 = mau_0_io_pipe_phv_out_data_419; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_420 = mau_0_io_pipe_phv_out_data_420; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_421 = mau_0_io_pipe_phv_out_data_421; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_422 = mau_0_io_pipe_phv_out_data_422; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_423 = mau_0_io_pipe_phv_out_data_423; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_424 = mau_0_io_pipe_phv_out_data_424; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_425 = mau_0_io_pipe_phv_out_data_425; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_426 = mau_0_io_pipe_phv_out_data_426; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_427 = mau_0_io_pipe_phv_out_data_427; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_428 = mau_0_io_pipe_phv_out_data_428; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_429 = mau_0_io_pipe_phv_out_data_429; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_430 = mau_0_io_pipe_phv_out_data_430; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_431 = mau_0_io_pipe_phv_out_data_431; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_432 = mau_0_io_pipe_phv_out_data_432; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_433 = mau_0_io_pipe_phv_out_data_433; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_434 = mau_0_io_pipe_phv_out_data_434; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_435 = mau_0_io_pipe_phv_out_data_435; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_436 = mau_0_io_pipe_phv_out_data_436; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_437 = mau_0_io_pipe_phv_out_data_437; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_438 = mau_0_io_pipe_phv_out_data_438; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_439 = mau_0_io_pipe_phv_out_data_439; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_440 = mau_0_io_pipe_phv_out_data_440; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_441 = mau_0_io_pipe_phv_out_data_441; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_442 = mau_0_io_pipe_phv_out_data_442; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_443 = mau_0_io_pipe_phv_out_data_443; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_444 = mau_0_io_pipe_phv_out_data_444; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_445 = mau_0_io_pipe_phv_out_data_445; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_446 = mau_0_io_pipe_phv_out_data_446; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_447 = mau_0_io_pipe_phv_out_data_447; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_448 = mau_0_io_pipe_phv_out_data_448; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_449 = mau_0_io_pipe_phv_out_data_449; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_450 = mau_0_io_pipe_phv_out_data_450; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_451 = mau_0_io_pipe_phv_out_data_451; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_452 = mau_0_io_pipe_phv_out_data_452; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_453 = mau_0_io_pipe_phv_out_data_453; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_454 = mau_0_io_pipe_phv_out_data_454; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_455 = mau_0_io_pipe_phv_out_data_455; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_456 = mau_0_io_pipe_phv_out_data_456; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_457 = mau_0_io_pipe_phv_out_data_457; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_458 = mau_0_io_pipe_phv_out_data_458; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_459 = mau_0_io_pipe_phv_out_data_459; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_460 = mau_0_io_pipe_phv_out_data_460; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_461 = mau_0_io_pipe_phv_out_data_461; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_462 = mau_0_io_pipe_phv_out_data_462; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_463 = mau_0_io_pipe_phv_out_data_463; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_464 = mau_0_io_pipe_phv_out_data_464; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_465 = mau_0_io_pipe_phv_out_data_465; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_466 = mau_0_io_pipe_phv_out_data_466; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_467 = mau_0_io_pipe_phv_out_data_467; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_468 = mau_0_io_pipe_phv_out_data_468; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_469 = mau_0_io_pipe_phv_out_data_469; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_470 = mau_0_io_pipe_phv_out_data_470; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_471 = mau_0_io_pipe_phv_out_data_471; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_472 = mau_0_io_pipe_phv_out_data_472; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_473 = mau_0_io_pipe_phv_out_data_473; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_474 = mau_0_io_pipe_phv_out_data_474; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_475 = mau_0_io_pipe_phv_out_data_475; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_476 = mau_0_io_pipe_phv_out_data_476; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_477 = mau_0_io_pipe_phv_out_data_477; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_478 = mau_0_io_pipe_phv_out_data_478; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_479 = mau_0_io_pipe_phv_out_data_479; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_480 = mau_0_io_pipe_phv_out_data_480; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_481 = mau_0_io_pipe_phv_out_data_481; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_482 = mau_0_io_pipe_phv_out_data_482; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_483 = mau_0_io_pipe_phv_out_data_483; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_484 = mau_0_io_pipe_phv_out_data_484; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_485 = mau_0_io_pipe_phv_out_data_485; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_486 = mau_0_io_pipe_phv_out_data_486; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_487 = mau_0_io_pipe_phv_out_data_487; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_488 = mau_0_io_pipe_phv_out_data_488; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_489 = mau_0_io_pipe_phv_out_data_489; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_490 = mau_0_io_pipe_phv_out_data_490; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_491 = mau_0_io_pipe_phv_out_data_491; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_492 = mau_0_io_pipe_phv_out_data_492; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_493 = mau_0_io_pipe_phv_out_data_493; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_494 = mau_0_io_pipe_phv_out_data_494; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_495 = mau_0_io_pipe_phv_out_data_495; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_496 = mau_0_io_pipe_phv_out_data_496; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_497 = mau_0_io_pipe_phv_out_data_497; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_498 = mau_0_io_pipe_phv_out_data_498; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_499 = mau_0_io_pipe_phv_out_data_499; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_500 = mau_0_io_pipe_phv_out_data_500; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_501 = mau_0_io_pipe_phv_out_data_501; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_502 = mau_0_io_pipe_phv_out_data_502; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_503 = mau_0_io_pipe_phv_out_data_503; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_504 = mau_0_io_pipe_phv_out_data_504; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_505 = mau_0_io_pipe_phv_out_data_505; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_506 = mau_0_io_pipe_phv_out_data_506; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_507 = mau_0_io_pipe_phv_out_data_507; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_508 = mau_0_io_pipe_phv_out_data_508; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_509 = mau_0_io_pipe_phv_out_data_509; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_510 = mau_0_io_pipe_phv_out_data_510; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_511 = mau_0_io_pipe_phv_out_data_511; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_header_0 = mau_0_io_pipe_phv_out_header_0; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_header_1 = mau_0_io_pipe_phv_out_header_1; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_header_2 = mau_0_io_pipe_phv_out_header_2; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_header_3 = mau_0_io_pipe_phv_out_header_3; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_header_4 = mau_0_io_pipe_phv_out_header_4; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_header_5 = mau_0_io_pipe_phv_out_header_5; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_header_6 = mau_0_io_pipe_phv_out_header_6; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_header_7 = mau_0_io_pipe_phv_out_header_7; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_header_8 = mau_0_io_pipe_phv_out_header_8; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_header_9 = mau_0_io_pipe_phv_out_header_9; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_header_10 = mau_0_io_pipe_phv_out_header_10; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_header_11 = mau_0_io_pipe_phv_out_header_11; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_header_12 = mau_0_io_pipe_phv_out_header_12; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_header_13 = mau_0_io_pipe_phv_out_header_13; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_header_14 = mau_0_io_pipe_phv_out_header_14; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_header_15 = mau_0_io_pipe_phv_out_header_15; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_parse_current_state = mau_0_io_pipe_phv_out_parse_current_state; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_parse_current_offset = mau_0_io_pipe_phv_out_parse_current_offset; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_parse_transition_field = mau_0_io_pipe_phv_out_parse_transition_field; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_next_processor_id = mau_0_io_pipe_phv_out_next_processor_id; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_next_config_id = mau_0_io_pipe_phv_out_next_config_id; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_is_valid_processor = mau_0_io_pipe_phv_out_is_valid_processor; // @[parser_pisa.scala 42:35]
  assign mau_1_io_mod_state_id_mod = io_mod_en ? io_mod_module_mod_state_id_mod & mod_j_1 :
    io_mod_module_mod_state_id_mod; // @[parser_pisa.scala 51:22 parser_pisa.scala 58:40 parser_pisa.scala 47:23]
  assign mau_1_io_mod_state_id = io_mod_module_mod_state_id; // @[parser_pisa.scala 47:23]
  assign mau_1_io_mod_sram_w_cs = io_mod_module_mod_sram_w_cs; // @[parser_pisa.scala 47:23]
  assign mau_1_io_mod_sram_w_en = io_mod_en ? io_mod_module_mod_sram_w_en & mod_j_1 : io_mod_module_mod_sram_w_en; // @[parser_pisa.scala 51:22 parser_pisa.scala 57:40 parser_pisa.scala 47:23]
  assign mau_1_io_mod_sram_w_addr = io_mod_module_mod_sram_w_addr; // @[parser_pisa.scala 47:23]
  assign mau_1_io_mod_sram_w_data = io_mod_module_mod_sram_w_data; // @[parser_pisa.scala 47:23]
  assign mau_2_clock = clock;
  assign mau_2_io_pipe_phv_in_data_0 = mau_1_io_pipe_phv_out_data_0; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_1 = mau_1_io_pipe_phv_out_data_1; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_2 = mau_1_io_pipe_phv_out_data_2; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_3 = mau_1_io_pipe_phv_out_data_3; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_4 = mau_1_io_pipe_phv_out_data_4; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_5 = mau_1_io_pipe_phv_out_data_5; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_6 = mau_1_io_pipe_phv_out_data_6; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_7 = mau_1_io_pipe_phv_out_data_7; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_8 = mau_1_io_pipe_phv_out_data_8; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_9 = mau_1_io_pipe_phv_out_data_9; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_10 = mau_1_io_pipe_phv_out_data_10; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_11 = mau_1_io_pipe_phv_out_data_11; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_12 = mau_1_io_pipe_phv_out_data_12; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_13 = mau_1_io_pipe_phv_out_data_13; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_14 = mau_1_io_pipe_phv_out_data_14; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_15 = mau_1_io_pipe_phv_out_data_15; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_16 = mau_1_io_pipe_phv_out_data_16; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_17 = mau_1_io_pipe_phv_out_data_17; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_18 = mau_1_io_pipe_phv_out_data_18; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_19 = mau_1_io_pipe_phv_out_data_19; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_20 = mau_1_io_pipe_phv_out_data_20; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_21 = mau_1_io_pipe_phv_out_data_21; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_22 = mau_1_io_pipe_phv_out_data_22; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_23 = mau_1_io_pipe_phv_out_data_23; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_24 = mau_1_io_pipe_phv_out_data_24; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_25 = mau_1_io_pipe_phv_out_data_25; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_26 = mau_1_io_pipe_phv_out_data_26; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_27 = mau_1_io_pipe_phv_out_data_27; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_28 = mau_1_io_pipe_phv_out_data_28; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_29 = mau_1_io_pipe_phv_out_data_29; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_30 = mau_1_io_pipe_phv_out_data_30; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_31 = mau_1_io_pipe_phv_out_data_31; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_32 = mau_1_io_pipe_phv_out_data_32; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_33 = mau_1_io_pipe_phv_out_data_33; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_34 = mau_1_io_pipe_phv_out_data_34; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_35 = mau_1_io_pipe_phv_out_data_35; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_36 = mau_1_io_pipe_phv_out_data_36; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_37 = mau_1_io_pipe_phv_out_data_37; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_38 = mau_1_io_pipe_phv_out_data_38; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_39 = mau_1_io_pipe_phv_out_data_39; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_40 = mau_1_io_pipe_phv_out_data_40; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_41 = mau_1_io_pipe_phv_out_data_41; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_42 = mau_1_io_pipe_phv_out_data_42; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_43 = mau_1_io_pipe_phv_out_data_43; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_44 = mau_1_io_pipe_phv_out_data_44; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_45 = mau_1_io_pipe_phv_out_data_45; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_46 = mau_1_io_pipe_phv_out_data_46; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_47 = mau_1_io_pipe_phv_out_data_47; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_48 = mau_1_io_pipe_phv_out_data_48; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_49 = mau_1_io_pipe_phv_out_data_49; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_50 = mau_1_io_pipe_phv_out_data_50; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_51 = mau_1_io_pipe_phv_out_data_51; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_52 = mau_1_io_pipe_phv_out_data_52; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_53 = mau_1_io_pipe_phv_out_data_53; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_54 = mau_1_io_pipe_phv_out_data_54; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_55 = mau_1_io_pipe_phv_out_data_55; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_56 = mau_1_io_pipe_phv_out_data_56; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_57 = mau_1_io_pipe_phv_out_data_57; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_58 = mau_1_io_pipe_phv_out_data_58; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_59 = mau_1_io_pipe_phv_out_data_59; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_60 = mau_1_io_pipe_phv_out_data_60; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_61 = mau_1_io_pipe_phv_out_data_61; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_62 = mau_1_io_pipe_phv_out_data_62; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_63 = mau_1_io_pipe_phv_out_data_63; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_64 = mau_1_io_pipe_phv_out_data_64; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_65 = mau_1_io_pipe_phv_out_data_65; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_66 = mau_1_io_pipe_phv_out_data_66; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_67 = mau_1_io_pipe_phv_out_data_67; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_68 = mau_1_io_pipe_phv_out_data_68; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_69 = mau_1_io_pipe_phv_out_data_69; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_70 = mau_1_io_pipe_phv_out_data_70; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_71 = mau_1_io_pipe_phv_out_data_71; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_72 = mau_1_io_pipe_phv_out_data_72; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_73 = mau_1_io_pipe_phv_out_data_73; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_74 = mau_1_io_pipe_phv_out_data_74; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_75 = mau_1_io_pipe_phv_out_data_75; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_76 = mau_1_io_pipe_phv_out_data_76; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_77 = mau_1_io_pipe_phv_out_data_77; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_78 = mau_1_io_pipe_phv_out_data_78; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_79 = mau_1_io_pipe_phv_out_data_79; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_80 = mau_1_io_pipe_phv_out_data_80; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_81 = mau_1_io_pipe_phv_out_data_81; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_82 = mau_1_io_pipe_phv_out_data_82; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_83 = mau_1_io_pipe_phv_out_data_83; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_84 = mau_1_io_pipe_phv_out_data_84; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_85 = mau_1_io_pipe_phv_out_data_85; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_86 = mau_1_io_pipe_phv_out_data_86; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_87 = mau_1_io_pipe_phv_out_data_87; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_88 = mau_1_io_pipe_phv_out_data_88; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_89 = mau_1_io_pipe_phv_out_data_89; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_90 = mau_1_io_pipe_phv_out_data_90; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_91 = mau_1_io_pipe_phv_out_data_91; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_92 = mau_1_io_pipe_phv_out_data_92; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_93 = mau_1_io_pipe_phv_out_data_93; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_94 = mau_1_io_pipe_phv_out_data_94; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_95 = mau_1_io_pipe_phv_out_data_95; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_96 = mau_1_io_pipe_phv_out_data_96; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_97 = mau_1_io_pipe_phv_out_data_97; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_98 = mau_1_io_pipe_phv_out_data_98; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_99 = mau_1_io_pipe_phv_out_data_99; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_100 = mau_1_io_pipe_phv_out_data_100; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_101 = mau_1_io_pipe_phv_out_data_101; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_102 = mau_1_io_pipe_phv_out_data_102; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_103 = mau_1_io_pipe_phv_out_data_103; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_104 = mau_1_io_pipe_phv_out_data_104; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_105 = mau_1_io_pipe_phv_out_data_105; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_106 = mau_1_io_pipe_phv_out_data_106; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_107 = mau_1_io_pipe_phv_out_data_107; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_108 = mau_1_io_pipe_phv_out_data_108; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_109 = mau_1_io_pipe_phv_out_data_109; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_110 = mau_1_io_pipe_phv_out_data_110; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_111 = mau_1_io_pipe_phv_out_data_111; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_112 = mau_1_io_pipe_phv_out_data_112; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_113 = mau_1_io_pipe_phv_out_data_113; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_114 = mau_1_io_pipe_phv_out_data_114; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_115 = mau_1_io_pipe_phv_out_data_115; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_116 = mau_1_io_pipe_phv_out_data_116; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_117 = mau_1_io_pipe_phv_out_data_117; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_118 = mau_1_io_pipe_phv_out_data_118; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_119 = mau_1_io_pipe_phv_out_data_119; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_120 = mau_1_io_pipe_phv_out_data_120; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_121 = mau_1_io_pipe_phv_out_data_121; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_122 = mau_1_io_pipe_phv_out_data_122; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_123 = mau_1_io_pipe_phv_out_data_123; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_124 = mau_1_io_pipe_phv_out_data_124; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_125 = mau_1_io_pipe_phv_out_data_125; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_126 = mau_1_io_pipe_phv_out_data_126; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_127 = mau_1_io_pipe_phv_out_data_127; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_128 = mau_1_io_pipe_phv_out_data_128; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_129 = mau_1_io_pipe_phv_out_data_129; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_130 = mau_1_io_pipe_phv_out_data_130; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_131 = mau_1_io_pipe_phv_out_data_131; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_132 = mau_1_io_pipe_phv_out_data_132; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_133 = mau_1_io_pipe_phv_out_data_133; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_134 = mau_1_io_pipe_phv_out_data_134; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_135 = mau_1_io_pipe_phv_out_data_135; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_136 = mau_1_io_pipe_phv_out_data_136; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_137 = mau_1_io_pipe_phv_out_data_137; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_138 = mau_1_io_pipe_phv_out_data_138; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_139 = mau_1_io_pipe_phv_out_data_139; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_140 = mau_1_io_pipe_phv_out_data_140; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_141 = mau_1_io_pipe_phv_out_data_141; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_142 = mau_1_io_pipe_phv_out_data_142; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_143 = mau_1_io_pipe_phv_out_data_143; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_144 = mau_1_io_pipe_phv_out_data_144; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_145 = mau_1_io_pipe_phv_out_data_145; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_146 = mau_1_io_pipe_phv_out_data_146; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_147 = mau_1_io_pipe_phv_out_data_147; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_148 = mau_1_io_pipe_phv_out_data_148; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_149 = mau_1_io_pipe_phv_out_data_149; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_150 = mau_1_io_pipe_phv_out_data_150; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_151 = mau_1_io_pipe_phv_out_data_151; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_152 = mau_1_io_pipe_phv_out_data_152; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_153 = mau_1_io_pipe_phv_out_data_153; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_154 = mau_1_io_pipe_phv_out_data_154; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_155 = mau_1_io_pipe_phv_out_data_155; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_156 = mau_1_io_pipe_phv_out_data_156; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_157 = mau_1_io_pipe_phv_out_data_157; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_158 = mau_1_io_pipe_phv_out_data_158; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_159 = mau_1_io_pipe_phv_out_data_159; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_160 = mau_1_io_pipe_phv_out_data_160; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_161 = mau_1_io_pipe_phv_out_data_161; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_162 = mau_1_io_pipe_phv_out_data_162; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_163 = mau_1_io_pipe_phv_out_data_163; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_164 = mau_1_io_pipe_phv_out_data_164; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_165 = mau_1_io_pipe_phv_out_data_165; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_166 = mau_1_io_pipe_phv_out_data_166; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_167 = mau_1_io_pipe_phv_out_data_167; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_168 = mau_1_io_pipe_phv_out_data_168; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_169 = mau_1_io_pipe_phv_out_data_169; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_170 = mau_1_io_pipe_phv_out_data_170; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_171 = mau_1_io_pipe_phv_out_data_171; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_172 = mau_1_io_pipe_phv_out_data_172; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_173 = mau_1_io_pipe_phv_out_data_173; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_174 = mau_1_io_pipe_phv_out_data_174; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_175 = mau_1_io_pipe_phv_out_data_175; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_176 = mau_1_io_pipe_phv_out_data_176; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_177 = mau_1_io_pipe_phv_out_data_177; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_178 = mau_1_io_pipe_phv_out_data_178; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_179 = mau_1_io_pipe_phv_out_data_179; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_180 = mau_1_io_pipe_phv_out_data_180; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_181 = mau_1_io_pipe_phv_out_data_181; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_182 = mau_1_io_pipe_phv_out_data_182; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_183 = mau_1_io_pipe_phv_out_data_183; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_184 = mau_1_io_pipe_phv_out_data_184; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_185 = mau_1_io_pipe_phv_out_data_185; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_186 = mau_1_io_pipe_phv_out_data_186; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_187 = mau_1_io_pipe_phv_out_data_187; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_188 = mau_1_io_pipe_phv_out_data_188; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_189 = mau_1_io_pipe_phv_out_data_189; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_190 = mau_1_io_pipe_phv_out_data_190; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_191 = mau_1_io_pipe_phv_out_data_191; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_192 = mau_1_io_pipe_phv_out_data_192; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_193 = mau_1_io_pipe_phv_out_data_193; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_194 = mau_1_io_pipe_phv_out_data_194; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_195 = mau_1_io_pipe_phv_out_data_195; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_196 = mau_1_io_pipe_phv_out_data_196; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_197 = mau_1_io_pipe_phv_out_data_197; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_198 = mau_1_io_pipe_phv_out_data_198; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_199 = mau_1_io_pipe_phv_out_data_199; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_200 = mau_1_io_pipe_phv_out_data_200; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_201 = mau_1_io_pipe_phv_out_data_201; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_202 = mau_1_io_pipe_phv_out_data_202; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_203 = mau_1_io_pipe_phv_out_data_203; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_204 = mau_1_io_pipe_phv_out_data_204; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_205 = mau_1_io_pipe_phv_out_data_205; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_206 = mau_1_io_pipe_phv_out_data_206; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_207 = mau_1_io_pipe_phv_out_data_207; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_208 = mau_1_io_pipe_phv_out_data_208; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_209 = mau_1_io_pipe_phv_out_data_209; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_210 = mau_1_io_pipe_phv_out_data_210; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_211 = mau_1_io_pipe_phv_out_data_211; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_212 = mau_1_io_pipe_phv_out_data_212; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_213 = mau_1_io_pipe_phv_out_data_213; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_214 = mau_1_io_pipe_phv_out_data_214; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_215 = mau_1_io_pipe_phv_out_data_215; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_216 = mau_1_io_pipe_phv_out_data_216; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_217 = mau_1_io_pipe_phv_out_data_217; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_218 = mau_1_io_pipe_phv_out_data_218; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_219 = mau_1_io_pipe_phv_out_data_219; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_220 = mau_1_io_pipe_phv_out_data_220; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_221 = mau_1_io_pipe_phv_out_data_221; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_222 = mau_1_io_pipe_phv_out_data_222; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_223 = mau_1_io_pipe_phv_out_data_223; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_224 = mau_1_io_pipe_phv_out_data_224; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_225 = mau_1_io_pipe_phv_out_data_225; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_226 = mau_1_io_pipe_phv_out_data_226; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_227 = mau_1_io_pipe_phv_out_data_227; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_228 = mau_1_io_pipe_phv_out_data_228; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_229 = mau_1_io_pipe_phv_out_data_229; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_230 = mau_1_io_pipe_phv_out_data_230; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_231 = mau_1_io_pipe_phv_out_data_231; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_232 = mau_1_io_pipe_phv_out_data_232; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_233 = mau_1_io_pipe_phv_out_data_233; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_234 = mau_1_io_pipe_phv_out_data_234; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_235 = mau_1_io_pipe_phv_out_data_235; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_236 = mau_1_io_pipe_phv_out_data_236; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_237 = mau_1_io_pipe_phv_out_data_237; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_238 = mau_1_io_pipe_phv_out_data_238; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_239 = mau_1_io_pipe_phv_out_data_239; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_240 = mau_1_io_pipe_phv_out_data_240; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_241 = mau_1_io_pipe_phv_out_data_241; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_242 = mau_1_io_pipe_phv_out_data_242; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_243 = mau_1_io_pipe_phv_out_data_243; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_244 = mau_1_io_pipe_phv_out_data_244; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_245 = mau_1_io_pipe_phv_out_data_245; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_246 = mau_1_io_pipe_phv_out_data_246; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_247 = mau_1_io_pipe_phv_out_data_247; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_248 = mau_1_io_pipe_phv_out_data_248; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_249 = mau_1_io_pipe_phv_out_data_249; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_250 = mau_1_io_pipe_phv_out_data_250; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_251 = mau_1_io_pipe_phv_out_data_251; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_252 = mau_1_io_pipe_phv_out_data_252; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_253 = mau_1_io_pipe_phv_out_data_253; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_254 = mau_1_io_pipe_phv_out_data_254; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_255 = mau_1_io_pipe_phv_out_data_255; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_256 = mau_1_io_pipe_phv_out_data_256; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_257 = mau_1_io_pipe_phv_out_data_257; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_258 = mau_1_io_pipe_phv_out_data_258; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_259 = mau_1_io_pipe_phv_out_data_259; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_260 = mau_1_io_pipe_phv_out_data_260; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_261 = mau_1_io_pipe_phv_out_data_261; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_262 = mau_1_io_pipe_phv_out_data_262; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_263 = mau_1_io_pipe_phv_out_data_263; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_264 = mau_1_io_pipe_phv_out_data_264; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_265 = mau_1_io_pipe_phv_out_data_265; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_266 = mau_1_io_pipe_phv_out_data_266; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_267 = mau_1_io_pipe_phv_out_data_267; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_268 = mau_1_io_pipe_phv_out_data_268; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_269 = mau_1_io_pipe_phv_out_data_269; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_270 = mau_1_io_pipe_phv_out_data_270; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_271 = mau_1_io_pipe_phv_out_data_271; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_272 = mau_1_io_pipe_phv_out_data_272; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_273 = mau_1_io_pipe_phv_out_data_273; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_274 = mau_1_io_pipe_phv_out_data_274; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_275 = mau_1_io_pipe_phv_out_data_275; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_276 = mau_1_io_pipe_phv_out_data_276; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_277 = mau_1_io_pipe_phv_out_data_277; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_278 = mau_1_io_pipe_phv_out_data_278; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_279 = mau_1_io_pipe_phv_out_data_279; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_280 = mau_1_io_pipe_phv_out_data_280; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_281 = mau_1_io_pipe_phv_out_data_281; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_282 = mau_1_io_pipe_phv_out_data_282; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_283 = mau_1_io_pipe_phv_out_data_283; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_284 = mau_1_io_pipe_phv_out_data_284; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_285 = mau_1_io_pipe_phv_out_data_285; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_286 = mau_1_io_pipe_phv_out_data_286; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_287 = mau_1_io_pipe_phv_out_data_287; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_288 = mau_1_io_pipe_phv_out_data_288; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_289 = mau_1_io_pipe_phv_out_data_289; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_290 = mau_1_io_pipe_phv_out_data_290; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_291 = mau_1_io_pipe_phv_out_data_291; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_292 = mau_1_io_pipe_phv_out_data_292; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_293 = mau_1_io_pipe_phv_out_data_293; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_294 = mau_1_io_pipe_phv_out_data_294; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_295 = mau_1_io_pipe_phv_out_data_295; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_296 = mau_1_io_pipe_phv_out_data_296; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_297 = mau_1_io_pipe_phv_out_data_297; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_298 = mau_1_io_pipe_phv_out_data_298; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_299 = mau_1_io_pipe_phv_out_data_299; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_300 = mau_1_io_pipe_phv_out_data_300; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_301 = mau_1_io_pipe_phv_out_data_301; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_302 = mau_1_io_pipe_phv_out_data_302; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_303 = mau_1_io_pipe_phv_out_data_303; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_304 = mau_1_io_pipe_phv_out_data_304; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_305 = mau_1_io_pipe_phv_out_data_305; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_306 = mau_1_io_pipe_phv_out_data_306; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_307 = mau_1_io_pipe_phv_out_data_307; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_308 = mau_1_io_pipe_phv_out_data_308; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_309 = mau_1_io_pipe_phv_out_data_309; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_310 = mau_1_io_pipe_phv_out_data_310; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_311 = mau_1_io_pipe_phv_out_data_311; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_312 = mau_1_io_pipe_phv_out_data_312; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_313 = mau_1_io_pipe_phv_out_data_313; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_314 = mau_1_io_pipe_phv_out_data_314; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_315 = mau_1_io_pipe_phv_out_data_315; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_316 = mau_1_io_pipe_phv_out_data_316; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_317 = mau_1_io_pipe_phv_out_data_317; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_318 = mau_1_io_pipe_phv_out_data_318; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_319 = mau_1_io_pipe_phv_out_data_319; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_320 = mau_1_io_pipe_phv_out_data_320; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_321 = mau_1_io_pipe_phv_out_data_321; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_322 = mau_1_io_pipe_phv_out_data_322; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_323 = mau_1_io_pipe_phv_out_data_323; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_324 = mau_1_io_pipe_phv_out_data_324; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_325 = mau_1_io_pipe_phv_out_data_325; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_326 = mau_1_io_pipe_phv_out_data_326; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_327 = mau_1_io_pipe_phv_out_data_327; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_328 = mau_1_io_pipe_phv_out_data_328; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_329 = mau_1_io_pipe_phv_out_data_329; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_330 = mau_1_io_pipe_phv_out_data_330; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_331 = mau_1_io_pipe_phv_out_data_331; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_332 = mau_1_io_pipe_phv_out_data_332; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_333 = mau_1_io_pipe_phv_out_data_333; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_334 = mau_1_io_pipe_phv_out_data_334; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_335 = mau_1_io_pipe_phv_out_data_335; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_336 = mau_1_io_pipe_phv_out_data_336; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_337 = mau_1_io_pipe_phv_out_data_337; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_338 = mau_1_io_pipe_phv_out_data_338; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_339 = mau_1_io_pipe_phv_out_data_339; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_340 = mau_1_io_pipe_phv_out_data_340; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_341 = mau_1_io_pipe_phv_out_data_341; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_342 = mau_1_io_pipe_phv_out_data_342; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_343 = mau_1_io_pipe_phv_out_data_343; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_344 = mau_1_io_pipe_phv_out_data_344; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_345 = mau_1_io_pipe_phv_out_data_345; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_346 = mau_1_io_pipe_phv_out_data_346; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_347 = mau_1_io_pipe_phv_out_data_347; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_348 = mau_1_io_pipe_phv_out_data_348; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_349 = mau_1_io_pipe_phv_out_data_349; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_350 = mau_1_io_pipe_phv_out_data_350; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_351 = mau_1_io_pipe_phv_out_data_351; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_352 = mau_1_io_pipe_phv_out_data_352; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_353 = mau_1_io_pipe_phv_out_data_353; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_354 = mau_1_io_pipe_phv_out_data_354; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_355 = mau_1_io_pipe_phv_out_data_355; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_356 = mau_1_io_pipe_phv_out_data_356; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_357 = mau_1_io_pipe_phv_out_data_357; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_358 = mau_1_io_pipe_phv_out_data_358; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_359 = mau_1_io_pipe_phv_out_data_359; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_360 = mau_1_io_pipe_phv_out_data_360; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_361 = mau_1_io_pipe_phv_out_data_361; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_362 = mau_1_io_pipe_phv_out_data_362; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_363 = mau_1_io_pipe_phv_out_data_363; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_364 = mau_1_io_pipe_phv_out_data_364; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_365 = mau_1_io_pipe_phv_out_data_365; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_366 = mau_1_io_pipe_phv_out_data_366; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_367 = mau_1_io_pipe_phv_out_data_367; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_368 = mau_1_io_pipe_phv_out_data_368; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_369 = mau_1_io_pipe_phv_out_data_369; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_370 = mau_1_io_pipe_phv_out_data_370; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_371 = mau_1_io_pipe_phv_out_data_371; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_372 = mau_1_io_pipe_phv_out_data_372; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_373 = mau_1_io_pipe_phv_out_data_373; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_374 = mau_1_io_pipe_phv_out_data_374; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_375 = mau_1_io_pipe_phv_out_data_375; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_376 = mau_1_io_pipe_phv_out_data_376; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_377 = mau_1_io_pipe_phv_out_data_377; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_378 = mau_1_io_pipe_phv_out_data_378; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_379 = mau_1_io_pipe_phv_out_data_379; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_380 = mau_1_io_pipe_phv_out_data_380; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_381 = mau_1_io_pipe_phv_out_data_381; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_382 = mau_1_io_pipe_phv_out_data_382; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_383 = mau_1_io_pipe_phv_out_data_383; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_384 = mau_1_io_pipe_phv_out_data_384; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_385 = mau_1_io_pipe_phv_out_data_385; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_386 = mau_1_io_pipe_phv_out_data_386; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_387 = mau_1_io_pipe_phv_out_data_387; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_388 = mau_1_io_pipe_phv_out_data_388; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_389 = mau_1_io_pipe_phv_out_data_389; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_390 = mau_1_io_pipe_phv_out_data_390; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_391 = mau_1_io_pipe_phv_out_data_391; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_392 = mau_1_io_pipe_phv_out_data_392; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_393 = mau_1_io_pipe_phv_out_data_393; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_394 = mau_1_io_pipe_phv_out_data_394; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_395 = mau_1_io_pipe_phv_out_data_395; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_396 = mau_1_io_pipe_phv_out_data_396; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_397 = mau_1_io_pipe_phv_out_data_397; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_398 = mau_1_io_pipe_phv_out_data_398; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_399 = mau_1_io_pipe_phv_out_data_399; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_400 = mau_1_io_pipe_phv_out_data_400; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_401 = mau_1_io_pipe_phv_out_data_401; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_402 = mau_1_io_pipe_phv_out_data_402; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_403 = mau_1_io_pipe_phv_out_data_403; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_404 = mau_1_io_pipe_phv_out_data_404; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_405 = mau_1_io_pipe_phv_out_data_405; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_406 = mau_1_io_pipe_phv_out_data_406; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_407 = mau_1_io_pipe_phv_out_data_407; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_408 = mau_1_io_pipe_phv_out_data_408; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_409 = mau_1_io_pipe_phv_out_data_409; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_410 = mau_1_io_pipe_phv_out_data_410; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_411 = mau_1_io_pipe_phv_out_data_411; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_412 = mau_1_io_pipe_phv_out_data_412; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_413 = mau_1_io_pipe_phv_out_data_413; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_414 = mau_1_io_pipe_phv_out_data_414; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_415 = mau_1_io_pipe_phv_out_data_415; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_416 = mau_1_io_pipe_phv_out_data_416; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_417 = mau_1_io_pipe_phv_out_data_417; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_418 = mau_1_io_pipe_phv_out_data_418; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_419 = mau_1_io_pipe_phv_out_data_419; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_420 = mau_1_io_pipe_phv_out_data_420; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_421 = mau_1_io_pipe_phv_out_data_421; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_422 = mau_1_io_pipe_phv_out_data_422; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_423 = mau_1_io_pipe_phv_out_data_423; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_424 = mau_1_io_pipe_phv_out_data_424; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_425 = mau_1_io_pipe_phv_out_data_425; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_426 = mau_1_io_pipe_phv_out_data_426; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_427 = mau_1_io_pipe_phv_out_data_427; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_428 = mau_1_io_pipe_phv_out_data_428; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_429 = mau_1_io_pipe_phv_out_data_429; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_430 = mau_1_io_pipe_phv_out_data_430; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_431 = mau_1_io_pipe_phv_out_data_431; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_432 = mau_1_io_pipe_phv_out_data_432; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_433 = mau_1_io_pipe_phv_out_data_433; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_434 = mau_1_io_pipe_phv_out_data_434; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_435 = mau_1_io_pipe_phv_out_data_435; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_436 = mau_1_io_pipe_phv_out_data_436; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_437 = mau_1_io_pipe_phv_out_data_437; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_438 = mau_1_io_pipe_phv_out_data_438; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_439 = mau_1_io_pipe_phv_out_data_439; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_440 = mau_1_io_pipe_phv_out_data_440; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_441 = mau_1_io_pipe_phv_out_data_441; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_442 = mau_1_io_pipe_phv_out_data_442; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_443 = mau_1_io_pipe_phv_out_data_443; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_444 = mau_1_io_pipe_phv_out_data_444; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_445 = mau_1_io_pipe_phv_out_data_445; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_446 = mau_1_io_pipe_phv_out_data_446; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_447 = mau_1_io_pipe_phv_out_data_447; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_448 = mau_1_io_pipe_phv_out_data_448; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_449 = mau_1_io_pipe_phv_out_data_449; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_450 = mau_1_io_pipe_phv_out_data_450; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_451 = mau_1_io_pipe_phv_out_data_451; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_452 = mau_1_io_pipe_phv_out_data_452; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_453 = mau_1_io_pipe_phv_out_data_453; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_454 = mau_1_io_pipe_phv_out_data_454; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_455 = mau_1_io_pipe_phv_out_data_455; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_456 = mau_1_io_pipe_phv_out_data_456; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_457 = mau_1_io_pipe_phv_out_data_457; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_458 = mau_1_io_pipe_phv_out_data_458; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_459 = mau_1_io_pipe_phv_out_data_459; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_460 = mau_1_io_pipe_phv_out_data_460; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_461 = mau_1_io_pipe_phv_out_data_461; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_462 = mau_1_io_pipe_phv_out_data_462; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_463 = mau_1_io_pipe_phv_out_data_463; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_464 = mau_1_io_pipe_phv_out_data_464; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_465 = mau_1_io_pipe_phv_out_data_465; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_466 = mau_1_io_pipe_phv_out_data_466; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_467 = mau_1_io_pipe_phv_out_data_467; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_468 = mau_1_io_pipe_phv_out_data_468; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_469 = mau_1_io_pipe_phv_out_data_469; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_470 = mau_1_io_pipe_phv_out_data_470; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_471 = mau_1_io_pipe_phv_out_data_471; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_472 = mau_1_io_pipe_phv_out_data_472; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_473 = mau_1_io_pipe_phv_out_data_473; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_474 = mau_1_io_pipe_phv_out_data_474; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_475 = mau_1_io_pipe_phv_out_data_475; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_476 = mau_1_io_pipe_phv_out_data_476; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_477 = mau_1_io_pipe_phv_out_data_477; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_478 = mau_1_io_pipe_phv_out_data_478; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_479 = mau_1_io_pipe_phv_out_data_479; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_480 = mau_1_io_pipe_phv_out_data_480; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_481 = mau_1_io_pipe_phv_out_data_481; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_482 = mau_1_io_pipe_phv_out_data_482; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_483 = mau_1_io_pipe_phv_out_data_483; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_484 = mau_1_io_pipe_phv_out_data_484; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_485 = mau_1_io_pipe_phv_out_data_485; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_486 = mau_1_io_pipe_phv_out_data_486; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_487 = mau_1_io_pipe_phv_out_data_487; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_488 = mau_1_io_pipe_phv_out_data_488; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_489 = mau_1_io_pipe_phv_out_data_489; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_490 = mau_1_io_pipe_phv_out_data_490; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_491 = mau_1_io_pipe_phv_out_data_491; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_492 = mau_1_io_pipe_phv_out_data_492; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_493 = mau_1_io_pipe_phv_out_data_493; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_494 = mau_1_io_pipe_phv_out_data_494; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_495 = mau_1_io_pipe_phv_out_data_495; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_496 = mau_1_io_pipe_phv_out_data_496; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_497 = mau_1_io_pipe_phv_out_data_497; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_498 = mau_1_io_pipe_phv_out_data_498; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_499 = mau_1_io_pipe_phv_out_data_499; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_500 = mau_1_io_pipe_phv_out_data_500; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_501 = mau_1_io_pipe_phv_out_data_501; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_502 = mau_1_io_pipe_phv_out_data_502; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_503 = mau_1_io_pipe_phv_out_data_503; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_504 = mau_1_io_pipe_phv_out_data_504; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_505 = mau_1_io_pipe_phv_out_data_505; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_506 = mau_1_io_pipe_phv_out_data_506; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_507 = mau_1_io_pipe_phv_out_data_507; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_508 = mau_1_io_pipe_phv_out_data_508; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_509 = mau_1_io_pipe_phv_out_data_509; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_510 = mau_1_io_pipe_phv_out_data_510; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_511 = mau_1_io_pipe_phv_out_data_511; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_header_0 = mau_1_io_pipe_phv_out_header_0; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_header_1 = mau_1_io_pipe_phv_out_header_1; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_header_2 = mau_1_io_pipe_phv_out_header_2; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_header_3 = mau_1_io_pipe_phv_out_header_3; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_header_4 = mau_1_io_pipe_phv_out_header_4; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_header_5 = mau_1_io_pipe_phv_out_header_5; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_header_6 = mau_1_io_pipe_phv_out_header_6; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_header_7 = mau_1_io_pipe_phv_out_header_7; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_header_8 = mau_1_io_pipe_phv_out_header_8; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_header_9 = mau_1_io_pipe_phv_out_header_9; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_header_10 = mau_1_io_pipe_phv_out_header_10; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_header_11 = mau_1_io_pipe_phv_out_header_11; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_header_12 = mau_1_io_pipe_phv_out_header_12; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_header_13 = mau_1_io_pipe_phv_out_header_13; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_header_14 = mau_1_io_pipe_phv_out_header_14; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_header_15 = mau_1_io_pipe_phv_out_header_15; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_parse_current_state = mau_1_io_pipe_phv_out_parse_current_state; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_parse_current_offset = mau_1_io_pipe_phv_out_parse_current_offset; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_parse_transition_field = mau_1_io_pipe_phv_out_parse_transition_field; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_next_processor_id = mau_1_io_pipe_phv_out_next_processor_id; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_next_config_id = mau_1_io_pipe_phv_out_next_config_id; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_is_valid_processor = mau_1_io_pipe_phv_out_is_valid_processor; // @[parser_pisa.scala 42:35]
  assign mau_2_io_mod_state_id_mod = io_mod_en ? io_mod_module_mod_state_id_mod & mod_j_2 :
    io_mod_module_mod_state_id_mod; // @[parser_pisa.scala 51:22 parser_pisa.scala 58:40 parser_pisa.scala 47:23]
  assign mau_2_io_mod_state_id = io_mod_module_mod_state_id; // @[parser_pisa.scala 47:23]
  assign mau_2_io_mod_sram_w_cs = io_mod_module_mod_sram_w_cs; // @[parser_pisa.scala 47:23]
  assign mau_2_io_mod_sram_w_en = io_mod_en ? io_mod_module_mod_sram_w_en & mod_j_2 : io_mod_module_mod_sram_w_en; // @[parser_pisa.scala 51:22 parser_pisa.scala 57:40 parser_pisa.scala 47:23]
  assign mau_2_io_mod_sram_w_addr = io_mod_module_mod_sram_w_addr; // @[parser_pisa.scala 47:23]
  assign mau_2_io_mod_sram_w_data = io_mod_module_mod_sram_w_data; // @[parser_pisa.scala 47:23]
  assign mau_3_clock = clock;
  assign mau_3_io_pipe_phv_in_data_0 = mau_2_io_pipe_phv_out_data_0; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_1 = mau_2_io_pipe_phv_out_data_1; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_2 = mau_2_io_pipe_phv_out_data_2; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_3 = mau_2_io_pipe_phv_out_data_3; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_4 = mau_2_io_pipe_phv_out_data_4; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_5 = mau_2_io_pipe_phv_out_data_5; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_6 = mau_2_io_pipe_phv_out_data_6; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_7 = mau_2_io_pipe_phv_out_data_7; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_8 = mau_2_io_pipe_phv_out_data_8; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_9 = mau_2_io_pipe_phv_out_data_9; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_10 = mau_2_io_pipe_phv_out_data_10; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_11 = mau_2_io_pipe_phv_out_data_11; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_12 = mau_2_io_pipe_phv_out_data_12; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_13 = mau_2_io_pipe_phv_out_data_13; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_14 = mau_2_io_pipe_phv_out_data_14; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_15 = mau_2_io_pipe_phv_out_data_15; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_16 = mau_2_io_pipe_phv_out_data_16; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_17 = mau_2_io_pipe_phv_out_data_17; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_18 = mau_2_io_pipe_phv_out_data_18; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_19 = mau_2_io_pipe_phv_out_data_19; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_20 = mau_2_io_pipe_phv_out_data_20; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_21 = mau_2_io_pipe_phv_out_data_21; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_22 = mau_2_io_pipe_phv_out_data_22; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_23 = mau_2_io_pipe_phv_out_data_23; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_24 = mau_2_io_pipe_phv_out_data_24; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_25 = mau_2_io_pipe_phv_out_data_25; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_26 = mau_2_io_pipe_phv_out_data_26; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_27 = mau_2_io_pipe_phv_out_data_27; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_28 = mau_2_io_pipe_phv_out_data_28; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_29 = mau_2_io_pipe_phv_out_data_29; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_30 = mau_2_io_pipe_phv_out_data_30; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_31 = mau_2_io_pipe_phv_out_data_31; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_32 = mau_2_io_pipe_phv_out_data_32; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_33 = mau_2_io_pipe_phv_out_data_33; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_34 = mau_2_io_pipe_phv_out_data_34; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_35 = mau_2_io_pipe_phv_out_data_35; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_36 = mau_2_io_pipe_phv_out_data_36; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_37 = mau_2_io_pipe_phv_out_data_37; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_38 = mau_2_io_pipe_phv_out_data_38; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_39 = mau_2_io_pipe_phv_out_data_39; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_40 = mau_2_io_pipe_phv_out_data_40; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_41 = mau_2_io_pipe_phv_out_data_41; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_42 = mau_2_io_pipe_phv_out_data_42; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_43 = mau_2_io_pipe_phv_out_data_43; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_44 = mau_2_io_pipe_phv_out_data_44; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_45 = mau_2_io_pipe_phv_out_data_45; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_46 = mau_2_io_pipe_phv_out_data_46; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_47 = mau_2_io_pipe_phv_out_data_47; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_48 = mau_2_io_pipe_phv_out_data_48; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_49 = mau_2_io_pipe_phv_out_data_49; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_50 = mau_2_io_pipe_phv_out_data_50; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_51 = mau_2_io_pipe_phv_out_data_51; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_52 = mau_2_io_pipe_phv_out_data_52; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_53 = mau_2_io_pipe_phv_out_data_53; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_54 = mau_2_io_pipe_phv_out_data_54; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_55 = mau_2_io_pipe_phv_out_data_55; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_56 = mau_2_io_pipe_phv_out_data_56; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_57 = mau_2_io_pipe_phv_out_data_57; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_58 = mau_2_io_pipe_phv_out_data_58; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_59 = mau_2_io_pipe_phv_out_data_59; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_60 = mau_2_io_pipe_phv_out_data_60; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_61 = mau_2_io_pipe_phv_out_data_61; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_62 = mau_2_io_pipe_phv_out_data_62; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_63 = mau_2_io_pipe_phv_out_data_63; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_64 = mau_2_io_pipe_phv_out_data_64; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_65 = mau_2_io_pipe_phv_out_data_65; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_66 = mau_2_io_pipe_phv_out_data_66; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_67 = mau_2_io_pipe_phv_out_data_67; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_68 = mau_2_io_pipe_phv_out_data_68; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_69 = mau_2_io_pipe_phv_out_data_69; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_70 = mau_2_io_pipe_phv_out_data_70; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_71 = mau_2_io_pipe_phv_out_data_71; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_72 = mau_2_io_pipe_phv_out_data_72; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_73 = mau_2_io_pipe_phv_out_data_73; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_74 = mau_2_io_pipe_phv_out_data_74; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_75 = mau_2_io_pipe_phv_out_data_75; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_76 = mau_2_io_pipe_phv_out_data_76; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_77 = mau_2_io_pipe_phv_out_data_77; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_78 = mau_2_io_pipe_phv_out_data_78; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_79 = mau_2_io_pipe_phv_out_data_79; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_80 = mau_2_io_pipe_phv_out_data_80; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_81 = mau_2_io_pipe_phv_out_data_81; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_82 = mau_2_io_pipe_phv_out_data_82; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_83 = mau_2_io_pipe_phv_out_data_83; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_84 = mau_2_io_pipe_phv_out_data_84; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_85 = mau_2_io_pipe_phv_out_data_85; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_86 = mau_2_io_pipe_phv_out_data_86; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_87 = mau_2_io_pipe_phv_out_data_87; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_88 = mau_2_io_pipe_phv_out_data_88; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_89 = mau_2_io_pipe_phv_out_data_89; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_90 = mau_2_io_pipe_phv_out_data_90; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_91 = mau_2_io_pipe_phv_out_data_91; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_92 = mau_2_io_pipe_phv_out_data_92; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_93 = mau_2_io_pipe_phv_out_data_93; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_94 = mau_2_io_pipe_phv_out_data_94; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_95 = mau_2_io_pipe_phv_out_data_95; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_96 = mau_2_io_pipe_phv_out_data_96; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_97 = mau_2_io_pipe_phv_out_data_97; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_98 = mau_2_io_pipe_phv_out_data_98; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_99 = mau_2_io_pipe_phv_out_data_99; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_100 = mau_2_io_pipe_phv_out_data_100; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_101 = mau_2_io_pipe_phv_out_data_101; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_102 = mau_2_io_pipe_phv_out_data_102; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_103 = mau_2_io_pipe_phv_out_data_103; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_104 = mau_2_io_pipe_phv_out_data_104; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_105 = mau_2_io_pipe_phv_out_data_105; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_106 = mau_2_io_pipe_phv_out_data_106; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_107 = mau_2_io_pipe_phv_out_data_107; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_108 = mau_2_io_pipe_phv_out_data_108; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_109 = mau_2_io_pipe_phv_out_data_109; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_110 = mau_2_io_pipe_phv_out_data_110; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_111 = mau_2_io_pipe_phv_out_data_111; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_112 = mau_2_io_pipe_phv_out_data_112; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_113 = mau_2_io_pipe_phv_out_data_113; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_114 = mau_2_io_pipe_phv_out_data_114; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_115 = mau_2_io_pipe_phv_out_data_115; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_116 = mau_2_io_pipe_phv_out_data_116; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_117 = mau_2_io_pipe_phv_out_data_117; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_118 = mau_2_io_pipe_phv_out_data_118; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_119 = mau_2_io_pipe_phv_out_data_119; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_120 = mau_2_io_pipe_phv_out_data_120; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_121 = mau_2_io_pipe_phv_out_data_121; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_122 = mau_2_io_pipe_phv_out_data_122; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_123 = mau_2_io_pipe_phv_out_data_123; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_124 = mau_2_io_pipe_phv_out_data_124; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_125 = mau_2_io_pipe_phv_out_data_125; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_126 = mau_2_io_pipe_phv_out_data_126; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_127 = mau_2_io_pipe_phv_out_data_127; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_128 = mau_2_io_pipe_phv_out_data_128; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_129 = mau_2_io_pipe_phv_out_data_129; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_130 = mau_2_io_pipe_phv_out_data_130; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_131 = mau_2_io_pipe_phv_out_data_131; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_132 = mau_2_io_pipe_phv_out_data_132; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_133 = mau_2_io_pipe_phv_out_data_133; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_134 = mau_2_io_pipe_phv_out_data_134; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_135 = mau_2_io_pipe_phv_out_data_135; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_136 = mau_2_io_pipe_phv_out_data_136; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_137 = mau_2_io_pipe_phv_out_data_137; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_138 = mau_2_io_pipe_phv_out_data_138; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_139 = mau_2_io_pipe_phv_out_data_139; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_140 = mau_2_io_pipe_phv_out_data_140; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_141 = mau_2_io_pipe_phv_out_data_141; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_142 = mau_2_io_pipe_phv_out_data_142; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_143 = mau_2_io_pipe_phv_out_data_143; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_144 = mau_2_io_pipe_phv_out_data_144; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_145 = mau_2_io_pipe_phv_out_data_145; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_146 = mau_2_io_pipe_phv_out_data_146; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_147 = mau_2_io_pipe_phv_out_data_147; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_148 = mau_2_io_pipe_phv_out_data_148; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_149 = mau_2_io_pipe_phv_out_data_149; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_150 = mau_2_io_pipe_phv_out_data_150; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_151 = mau_2_io_pipe_phv_out_data_151; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_152 = mau_2_io_pipe_phv_out_data_152; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_153 = mau_2_io_pipe_phv_out_data_153; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_154 = mau_2_io_pipe_phv_out_data_154; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_155 = mau_2_io_pipe_phv_out_data_155; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_156 = mau_2_io_pipe_phv_out_data_156; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_157 = mau_2_io_pipe_phv_out_data_157; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_158 = mau_2_io_pipe_phv_out_data_158; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_159 = mau_2_io_pipe_phv_out_data_159; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_160 = mau_2_io_pipe_phv_out_data_160; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_161 = mau_2_io_pipe_phv_out_data_161; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_162 = mau_2_io_pipe_phv_out_data_162; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_163 = mau_2_io_pipe_phv_out_data_163; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_164 = mau_2_io_pipe_phv_out_data_164; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_165 = mau_2_io_pipe_phv_out_data_165; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_166 = mau_2_io_pipe_phv_out_data_166; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_167 = mau_2_io_pipe_phv_out_data_167; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_168 = mau_2_io_pipe_phv_out_data_168; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_169 = mau_2_io_pipe_phv_out_data_169; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_170 = mau_2_io_pipe_phv_out_data_170; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_171 = mau_2_io_pipe_phv_out_data_171; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_172 = mau_2_io_pipe_phv_out_data_172; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_173 = mau_2_io_pipe_phv_out_data_173; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_174 = mau_2_io_pipe_phv_out_data_174; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_175 = mau_2_io_pipe_phv_out_data_175; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_176 = mau_2_io_pipe_phv_out_data_176; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_177 = mau_2_io_pipe_phv_out_data_177; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_178 = mau_2_io_pipe_phv_out_data_178; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_179 = mau_2_io_pipe_phv_out_data_179; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_180 = mau_2_io_pipe_phv_out_data_180; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_181 = mau_2_io_pipe_phv_out_data_181; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_182 = mau_2_io_pipe_phv_out_data_182; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_183 = mau_2_io_pipe_phv_out_data_183; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_184 = mau_2_io_pipe_phv_out_data_184; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_185 = mau_2_io_pipe_phv_out_data_185; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_186 = mau_2_io_pipe_phv_out_data_186; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_187 = mau_2_io_pipe_phv_out_data_187; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_188 = mau_2_io_pipe_phv_out_data_188; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_189 = mau_2_io_pipe_phv_out_data_189; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_190 = mau_2_io_pipe_phv_out_data_190; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_191 = mau_2_io_pipe_phv_out_data_191; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_192 = mau_2_io_pipe_phv_out_data_192; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_193 = mau_2_io_pipe_phv_out_data_193; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_194 = mau_2_io_pipe_phv_out_data_194; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_195 = mau_2_io_pipe_phv_out_data_195; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_196 = mau_2_io_pipe_phv_out_data_196; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_197 = mau_2_io_pipe_phv_out_data_197; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_198 = mau_2_io_pipe_phv_out_data_198; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_199 = mau_2_io_pipe_phv_out_data_199; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_200 = mau_2_io_pipe_phv_out_data_200; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_201 = mau_2_io_pipe_phv_out_data_201; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_202 = mau_2_io_pipe_phv_out_data_202; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_203 = mau_2_io_pipe_phv_out_data_203; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_204 = mau_2_io_pipe_phv_out_data_204; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_205 = mau_2_io_pipe_phv_out_data_205; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_206 = mau_2_io_pipe_phv_out_data_206; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_207 = mau_2_io_pipe_phv_out_data_207; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_208 = mau_2_io_pipe_phv_out_data_208; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_209 = mau_2_io_pipe_phv_out_data_209; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_210 = mau_2_io_pipe_phv_out_data_210; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_211 = mau_2_io_pipe_phv_out_data_211; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_212 = mau_2_io_pipe_phv_out_data_212; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_213 = mau_2_io_pipe_phv_out_data_213; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_214 = mau_2_io_pipe_phv_out_data_214; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_215 = mau_2_io_pipe_phv_out_data_215; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_216 = mau_2_io_pipe_phv_out_data_216; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_217 = mau_2_io_pipe_phv_out_data_217; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_218 = mau_2_io_pipe_phv_out_data_218; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_219 = mau_2_io_pipe_phv_out_data_219; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_220 = mau_2_io_pipe_phv_out_data_220; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_221 = mau_2_io_pipe_phv_out_data_221; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_222 = mau_2_io_pipe_phv_out_data_222; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_223 = mau_2_io_pipe_phv_out_data_223; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_224 = mau_2_io_pipe_phv_out_data_224; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_225 = mau_2_io_pipe_phv_out_data_225; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_226 = mau_2_io_pipe_phv_out_data_226; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_227 = mau_2_io_pipe_phv_out_data_227; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_228 = mau_2_io_pipe_phv_out_data_228; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_229 = mau_2_io_pipe_phv_out_data_229; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_230 = mau_2_io_pipe_phv_out_data_230; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_231 = mau_2_io_pipe_phv_out_data_231; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_232 = mau_2_io_pipe_phv_out_data_232; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_233 = mau_2_io_pipe_phv_out_data_233; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_234 = mau_2_io_pipe_phv_out_data_234; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_235 = mau_2_io_pipe_phv_out_data_235; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_236 = mau_2_io_pipe_phv_out_data_236; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_237 = mau_2_io_pipe_phv_out_data_237; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_238 = mau_2_io_pipe_phv_out_data_238; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_239 = mau_2_io_pipe_phv_out_data_239; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_240 = mau_2_io_pipe_phv_out_data_240; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_241 = mau_2_io_pipe_phv_out_data_241; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_242 = mau_2_io_pipe_phv_out_data_242; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_243 = mau_2_io_pipe_phv_out_data_243; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_244 = mau_2_io_pipe_phv_out_data_244; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_245 = mau_2_io_pipe_phv_out_data_245; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_246 = mau_2_io_pipe_phv_out_data_246; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_247 = mau_2_io_pipe_phv_out_data_247; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_248 = mau_2_io_pipe_phv_out_data_248; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_249 = mau_2_io_pipe_phv_out_data_249; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_250 = mau_2_io_pipe_phv_out_data_250; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_251 = mau_2_io_pipe_phv_out_data_251; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_252 = mau_2_io_pipe_phv_out_data_252; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_253 = mau_2_io_pipe_phv_out_data_253; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_254 = mau_2_io_pipe_phv_out_data_254; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_255 = mau_2_io_pipe_phv_out_data_255; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_256 = mau_2_io_pipe_phv_out_data_256; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_257 = mau_2_io_pipe_phv_out_data_257; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_258 = mau_2_io_pipe_phv_out_data_258; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_259 = mau_2_io_pipe_phv_out_data_259; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_260 = mau_2_io_pipe_phv_out_data_260; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_261 = mau_2_io_pipe_phv_out_data_261; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_262 = mau_2_io_pipe_phv_out_data_262; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_263 = mau_2_io_pipe_phv_out_data_263; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_264 = mau_2_io_pipe_phv_out_data_264; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_265 = mau_2_io_pipe_phv_out_data_265; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_266 = mau_2_io_pipe_phv_out_data_266; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_267 = mau_2_io_pipe_phv_out_data_267; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_268 = mau_2_io_pipe_phv_out_data_268; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_269 = mau_2_io_pipe_phv_out_data_269; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_270 = mau_2_io_pipe_phv_out_data_270; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_271 = mau_2_io_pipe_phv_out_data_271; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_272 = mau_2_io_pipe_phv_out_data_272; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_273 = mau_2_io_pipe_phv_out_data_273; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_274 = mau_2_io_pipe_phv_out_data_274; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_275 = mau_2_io_pipe_phv_out_data_275; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_276 = mau_2_io_pipe_phv_out_data_276; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_277 = mau_2_io_pipe_phv_out_data_277; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_278 = mau_2_io_pipe_phv_out_data_278; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_279 = mau_2_io_pipe_phv_out_data_279; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_280 = mau_2_io_pipe_phv_out_data_280; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_281 = mau_2_io_pipe_phv_out_data_281; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_282 = mau_2_io_pipe_phv_out_data_282; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_283 = mau_2_io_pipe_phv_out_data_283; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_284 = mau_2_io_pipe_phv_out_data_284; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_285 = mau_2_io_pipe_phv_out_data_285; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_286 = mau_2_io_pipe_phv_out_data_286; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_287 = mau_2_io_pipe_phv_out_data_287; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_288 = mau_2_io_pipe_phv_out_data_288; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_289 = mau_2_io_pipe_phv_out_data_289; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_290 = mau_2_io_pipe_phv_out_data_290; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_291 = mau_2_io_pipe_phv_out_data_291; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_292 = mau_2_io_pipe_phv_out_data_292; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_293 = mau_2_io_pipe_phv_out_data_293; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_294 = mau_2_io_pipe_phv_out_data_294; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_295 = mau_2_io_pipe_phv_out_data_295; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_296 = mau_2_io_pipe_phv_out_data_296; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_297 = mau_2_io_pipe_phv_out_data_297; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_298 = mau_2_io_pipe_phv_out_data_298; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_299 = mau_2_io_pipe_phv_out_data_299; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_300 = mau_2_io_pipe_phv_out_data_300; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_301 = mau_2_io_pipe_phv_out_data_301; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_302 = mau_2_io_pipe_phv_out_data_302; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_303 = mau_2_io_pipe_phv_out_data_303; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_304 = mau_2_io_pipe_phv_out_data_304; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_305 = mau_2_io_pipe_phv_out_data_305; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_306 = mau_2_io_pipe_phv_out_data_306; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_307 = mau_2_io_pipe_phv_out_data_307; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_308 = mau_2_io_pipe_phv_out_data_308; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_309 = mau_2_io_pipe_phv_out_data_309; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_310 = mau_2_io_pipe_phv_out_data_310; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_311 = mau_2_io_pipe_phv_out_data_311; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_312 = mau_2_io_pipe_phv_out_data_312; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_313 = mau_2_io_pipe_phv_out_data_313; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_314 = mau_2_io_pipe_phv_out_data_314; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_315 = mau_2_io_pipe_phv_out_data_315; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_316 = mau_2_io_pipe_phv_out_data_316; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_317 = mau_2_io_pipe_phv_out_data_317; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_318 = mau_2_io_pipe_phv_out_data_318; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_319 = mau_2_io_pipe_phv_out_data_319; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_320 = mau_2_io_pipe_phv_out_data_320; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_321 = mau_2_io_pipe_phv_out_data_321; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_322 = mau_2_io_pipe_phv_out_data_322; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_323 = mau_2_io_pipe_phv_out_data_323; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_324 = mau_2_io_pipe_phv_out_data_324; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_325 = mau_2_io_pipe_phv_out_data_325; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_326 = mau_2_io_pipe_phv_out_data_326; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_327 = mau_2_io_pipe_phv_out_data_327; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_328 = mau_2_io_pipe_phv_out_data_328; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_329 = mau_2_io_pipe_phv_out_data_329; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_330 = mau_2_io_pipe_phv_out_data_330; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_331 = mau_2_io_pipe_phv_out_data_331; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_332 = mau_2_io_pipe_phv_out_data_332; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_333 = mau_2_io_pipe_phv_out_data_333; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_334 = mau_2_io_pipe_phv_out_data_334; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_335 = mau_2_io_pipe_phv_out_data_335; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_336 = mau_2_io_pipe_phv_out_data_336; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_337 = mau_2_io_pipe_phv_out_data_337; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_338 = mau_2_io_pipe_phv_out_data_338; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_339 = mau_2_io_pipe_phv_out_data_339; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_340 = mau_2_io_pipe_phv_out_data_340; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_341 = mau_2_io_pipe_phv_out_data_341; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_342 = mau_2_io_pipe_phv_out_data_342; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_343 = mau_2_io_pipe_phv_out_data_343; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_344 = mau_2_io_pipe_phv_out_data_344; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_345 = mau_2_io_pipe_phv_out_data_345; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_346 = mau_2_io_pipe_phv_out_data_346; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_347 = mau_2_io_pipe_phv_out_data_347; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_348 = mau_2_io_pipe_phv_out_data_348; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_349 = mau_2_io_pipe_phv_out_data_349; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_350 = mau_2_io_pipe_phv_out_data_350; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_351 = mau_2_io_pipe_phv_out_data_351; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_352 = mau_2_io_pipe_phv_out_data_352; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_353 = mau_2_io_pipe_phv_out_data_353; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_354 = mau_2_io_pipe_phv_out_data_354; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_355 = mau_2_io_pipe_phv_out_data_355; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_356 = mau_2_io_pipe_phv_out_data_356; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_357 = mau_2_io_pipe_phv_out_data_357; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_358 = mau_2_io_pipe_phv_out_data_358; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_359 = mau_2_io_pipe_phv_out_data_359; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_360 = mau_2_io_pipe_phv_out_data_360; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_361 = mau_2_io_pipe_phv_out_data_361; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_362 = mau_2_io_pipe_phv_out_data_362; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_363 = mau_2_io_pipe_phv_out_data_363; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_364 = mau_2_io_pipe_phv_out_data_364; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_365 = mau_2_io_pipe_phv_out_data_365; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_366 = mau_2_io_pipe_phv_out_data_366; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_367 = mau_2_io_pipe_phv_out_data_367; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_368 = mau_2_io_pipe_phv_out_data_368; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_369 = mau_2_io_pipe_phv_out_data_369; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_370 = mau_2_io_pipe_phv_out_data_370; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_371 = mau_2_io_pipe_phv_out_data_371; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_372 = mau_2_io_pipe_phv_out_data_372; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_373 = mau_2_io_pipe_phv_out_data_373; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_374 = mau_2_io_pipe_phv_out_data_374; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_375 = mau_2_io_pipe_phv_out_data_375; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_376 = mau_2_io_pipe_phv_out_data_376; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_377 = mau_2_io_pipe_phv_out_data_377; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_378 = mau_2_io_pipe_phv_out_data_378; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_379 = mau_2_io_pipe_phv_out_data_379; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_380 = mau_2_io_pipe_phv_out_data_380; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_381 = mau_2_io_pipe_phv_out_data_381; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_382 = mau_2_io_pipe_phv_out_data_382; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_383 = mau_2_io_pipe_phv_out_data_383; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_384 = mau_2_io_pipe_phv_out_data_384; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_385 = mau_2_io_pipe_phv_out_data_385; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_386 = mau_2_io_pipe_phv_out_data_386; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_387 = mau_2_io_pipe_phv_out_data_387; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_388 = mau_2_io_pipe_phv_out_data_388; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_389 = mau_2_io_pipe_phv_out_data_389; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_390 = mau_2_io_pipe_phv_out_data_390; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_391 = mau_2_io_pipe_phv_out_data_391; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_392 = mau_2_io_pipe_phv_out_data_392; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_393 = mau_2_io_pipe_phv_out_data_393; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_394 = mau_2_io_pipe_phv_out_data_394; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_395 = mau_2_io_pipe_phv_out_data_395; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_396 = mau_2_io_pipe_phv_out_data_396; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_397 = mau_2_io_pipe_phv_out_data_397; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_398 = mau_2_io_pipe_phv_out_data_398; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_399 = mau_2_io_pipe_phv_out_data_399; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_400 = mau_2_io_pipe_phv_out_data_400; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_401 = mau_2_io_pipe_phv_out_data_401; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_402 = mau_2_io_pipe_phv_out_data_402; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_403 = mau_2_io_pipe_phv_out_data_403; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_404 = mau_2_io_pipe_phv_out_data_404; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_405 = mau_2_io_pipe_phv_out_data_405; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_406 = mau_2_io_pipe_phv_out_data_406; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_407 = mau_2_io_pipe_phv_out_data_407; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_408 = mau_2_io_pipe_phv_out_data_408; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_409 = mau_2_io_pipe_phv_out_data_409; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_410 = mau_2_io_pipe_phv_out_data_410; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_411 = mau_2_io_pipe_phv_out_data_411; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_412 = mau_2_io_pipe_phv_out_data_412; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_413 = mau_2_io_pipe_phv_out_data_413; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_414 = mau_2_io_pipe_phv_out_data_414; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_415 = mau_2_io_pipe_phv_out_data_415; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_416 = mau_2_io_pipe_phv_out_data_416; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_417 = mau_2_io_pipe_phv_out_data_417; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_418 = mau_2_io_pipe_phv_out_data_418; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_419 = mau_2_io_pipe_phv_out_data_419; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_420 = mau_2_io_pipe_phv_out_data_420; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_421 = mau_2_io_pipe_phv_out_data_421; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_422 = mau_2_io_pipe_phv_out_data_422; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_423 = mau_2_io_pipe_phv_out_data_423; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_424 = mau_2_io_pipe_phv_out_data_424; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_425 = mau_2_io_pipe_phv_out_data_425; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_426 = mau_2_io_pipe_phv_out_data_426; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_427 = mau_2_io_pipe_phv_out_data_427; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_428 = mau_2_io_pipe_phv_out_data_428; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_429 = mau_2_io_pipe_phv_out_data_429; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_430 = mau_2_io_pipe_phv_out_data_430; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_431 = mau_2_io_pipe_phv_out_data_431; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_432 = mau_2_io_pipe_phv_out_data_432; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_433 = mau_2_io_pipe_phv_out_data_433; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_434 = mau_2_io_pipe_phv_out_data_434; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_435 = mau_2_io_pipe_phv_out_data_435; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_436 = mau_2_io_pipe_phv_out_data_436; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_437 = mau_2_io_pipe_phv_out_data_437; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_438 = mau_2_io_pipe_phv_out_data_438; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_439 = mau_2_io_pipe_phv_out_data_439; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_440 = mau_2_io_pipe_phv_out_data_440; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_441 = mau_2_io_pipe_phv_out_data_441; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_442 = mau_2_io_pipe_phv_out_data_442; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_443 = mau_2_io_pipe_phv_out_data_443; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_444 = mau_2_io_pipe_phv_out_data_444; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_445 = mau_2_io_pipe_phv_out_data_445; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_446 = mau_2_io_pipe_phv_out_data_446; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_447 = mau_2_io_pipe_phv_out_data_447; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_448 = mau_2_io_pipe_phv_out_data_448; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_449 = mau_2_io_pipe_phv_out_data_449; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_450 = mau_2_io_pipe_phv_out_data_450; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_451 = mau_2_io_pipe_phv_out_data_451; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_452 = mau_2_io_pipe_phv_out_data_452; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_453 = mau_2_io_pipe_phv_out_data_453; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_454 = mau_2_io_pipe_phv_out_data_454; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_455 = mau_2_io_pipe_phv_out_data_455; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_456 = mau_2_io_pipe_phv_out_data_456; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_457 = mau_2_io_pipe_phv_out_data_457; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_458 = mau_2_io_pipe_phv_out_data_458; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_459 = mau_2_io_pipe_phv_out_data_459; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_460 = mau_2_io_pipe_phv_out_data_460; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_461 = mau_2_io_pipe_phv_out_data_461; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_462 = mau_2_io_pipe_phv_out_data_462; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_463 = mau_2_io_pipe_phv_out_data_463; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_464 = mau_2_io_pipe_phv_out_data_464; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_465 = mau_2_io_pipe_phv_out_data_465; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_466 = mau_2_io_pipe_phv_out_data_466; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_467 = mau_2_io_pipe_phv_out_data_467; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_468 = mau_2_io_pipe_phv_out_data_468; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_469 = mau_2_io_pipe_phv_out_data_469; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_470 = mau_2_io_pipe_phv_out_data_470; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_471 = mau_2_io_pipe_phv_out_data_471; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_472 = mau_2_io_pipe_phv_out_data_472; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_473 = mau_2_io_pipe_phv_out_data_473; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_474 = mau_2_io_pipe_phv_out_data_474; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_475 = mau_2_io_pipe_phv_out_data_475; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_476 = mau_2_io_pipe_phv_out_data_476; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_477 = mau_2_io_pipe_phv_out_data_477; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_478 = mau_2_io_pipe_phv_out_data_478; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_479 = mau_2_io_pipe_phv_out_data_479; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_480 = mau_2_io_pipe_phv_out_data_480; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_481 = mau_2_io_pipe_phv_out_data_481; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_482 = mau_2_io_pipe_phv_out_data_482; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_483 = mau_2_io_pipe_phv_out_data_483; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_484 = mau_2_io_pipe_phv_out_data_484; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_485 = mau_2_io_pipe_phv_out_data_485; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_486 = mau_2_io_pipe_phv_out_data_486; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_487 = mau_2_io_pipe_phv_out_data_487; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_488 = mau_2_io_pipe_phv_out_data_488; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_489 = mau_2_io_pipe_phv_out_data_489; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_490 = mau_2_io_pipe_phv_out_data_490; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_491 = mau_2_io_pipe_phv_out_data_491; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_492 = mau_2_io_pipe_phv_out_data_492; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_493 = mau_2_io_pipe_phv_out_data_493; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_494 = mau_2_io_pipe_phv_out_data_494; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_495 = mau_2_io_pipe_phv_out_data_495; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_496 = mau_2_io_pipe_phv_out_data_496; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_497 = mau_2_io_pipe_phv_out_data_497; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_498 = mau_2_io_pipe_phv_out_data_498; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_499 = mau_2_io_pipe_phv_out_data_499; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_500 = mau_2_io_pipe_phv_out_data_500; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_501 = mau_2_io_pipe_phv_out_data_501; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_502 = mau_2_io_pipe_phv_out_data_502; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_503 = mau_2_io_pipe_phv_out_data_503; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_504 = mau_2_io_pipe_phv_out_data_504; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_505 = mau_2_io_pipe_phv_out_data_505; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_506 = mau_2_io_pipe_phv_out_data_506; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_507 = mau_2_io_pipe_phv_out_data_507; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_508 = mau_2_io_pipe_phv_out_data_508; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_509 = mau_2_io_pipe_phv_out_data_509; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_510 = mau_2_io_pipe_phv_out_data_510; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_511 = mau_2_io_pipe_phv_out_data_511; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_header_0 = mau_2_io_pipe_phv_out_header_0; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_header_1 = mau_2_io_pipe_phv_out_header_1; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_header_2 = mau_2_io_pipe_phv_out_header_2; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_header_3 = mau_2_io_pipe_phv_out_header_3; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_header_4 = mau_2_io_pipe_phv_out_header_4; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_header_5 = mau_2_io_pipe_phv_out_header_5; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_header_6 = mau_2_io_pipe_phv_out_header_6; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_header_7 = mau_2_io_pipe_phv_out_header_7; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_header_8 = mau_2_io_pipe_phv_out_header_8; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_header_9 = mau_2_io_pipe_phv_out_header_9; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_header_10 = mau_2_io_pipe_phv_out_header_10; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_header_11 = mau_2_io_pipe_phv_out_header_11; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_header_12 = mau_2_io_pipe_phv_out_header_12; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_header_13 = mau_2_io_pipe_phv_out_header_13; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_header_14 = mau_2_io_pipe_phv_out_header_14; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_header_15 = mau_2_io_pipe_phv_out_header_15; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_parse_current_state = mau_2_io_pipe_phv_out_parse_current_state; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_parse_current_offset = mau_2_io_pipe_phv_out_parse_current_offset; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_parse_transition_field = mau_2_io_pipe_phv_out_parse_transition_field; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_next_processor_id = mau_2_io_pipe_phv_out_next_processor_id; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_next_config_id = mau_2_io_pipe_phv_out_next_config_id; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_is_valid_processor = mau_2_io_pipe_phv_out_is_valid_processor; // @[parser_pisa.scala 42:35]
  assign mau_3_io_mod_state_id_mod = io_mod_en ? io_mod_module_mod_state_id_mod & mod_j_3 :
    io_mod_module_mod_state_id_mod; // @[parser_pisa.scala 51:22 parser_pisa.scala 58:40 parser_pisa.scala 47:23]
  assign mau_3_io_mod_state_id = io_mod_module_mod_state_id; // @[parser_pisa.scala 47:23]
  assign mau_3_io_mod_sram_w_cs = io_mod_module_mod_sram_w_cs; // @[parser_pisa.scala 47:23]
  assign mau_3_io_mod_sram_w_en = io_mod_en ? io_mod_module_mod_sram_w_en & mod_j_3 : io_mod_module_mod_sram_w_en; // @[parser_pisa.scala 51:22 parser_pisa.scala 57:40 parser_pisa.scala 47:23]
  assign mau_3_io_mod_sram_w_addr = io_mod_module_mod_sram_w_addr; // @[parser_pisa.scala 47:23]
  assign mau_3_io_mod_sram_w_data = io_mod_module_mod_sram_w_data; // @[parser_pisa.scala 47:23]
  assign mau_4_clock = clock;
  assign mau_4_io_pipe_phv_in_data_0 = mau_3_io_pipe_phv_out_data_0; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_1 = mau_3_io_pipe_phv_out_data_1; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_2 = mau_3_io_pipe_phv_out_data_2; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_3 = mau_3_io_pipe_phv_out_data_3; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_4 = mau_3_io_pipe_phv_out_data_4; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_5 = mau_3_io_pipe_phv_out_data_5; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_6 = mau_3_io_pipe_phv_out_data_6; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_7 = mau_3_io_pipe_phv_out_data_7; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_8 = mau_3_io_pipe_phv_out_data_8; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_9 = mau_3_io_pipe_phv_out_data_9; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_10 = mau_3_io_pipe_phv_out_data_10; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_11 = mau_3_io_pipe_phv_out_data_11; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_12 = mau_3_io_pipe_phv_out_data_12; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_13 = mau_3_io_pipe_phv_out_data_13; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_14 = mau_3_io_pipe_phv_out_data_14; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_15 = mau_3_io_pipe_phv_out_data_15; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_16 = mau_3_io_pipe_phv_out_data_16; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_17 = mau_3_io_pipe_phv_out_data_17; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_18 = mau_3_io_pipe_phv_out_data_18; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_19 = mau_3_io_pipe_phv_out_data_19; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_20 = mau_3_io_pipe_phv_out_data_20; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_21 = mau_3_io_pipe_phv_out_data_21; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_22 = mau_3_io_pipe_phv_out_data_22; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_23 = mau_3_io_pipe_phv_out_data_23; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_24 = mau_3_io_pipe_phv_out_data_24; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_25 = mau_3_io_pipe_phv_out_data_25; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_26 = mau_3_io_pipe_phv_out_data_26; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_27 = mau_3_io_pipe_phv_out_data_27; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_28 = mau_3_io_pipe_phv_out_data_28; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_29 = mau_3_io_pipe_phv_out_data_29; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_30 = mau_3_io_pipe_phv_out_data_30; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_31 = mau_3_io_pipe_phv_out_data_31; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_32 = mau_3_io_pipe_phv_out_data_32; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_33 = mau_3_io_pipe_phv_out_data_33; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_34 = mau_3_io_pipe_phv_out_data_34; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_35 = mau_3_io_pipe_phv_out_data_35; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_36 = mau_3_io_pipe_phv_out_data_36; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_37 = mau_3_io_pipe_phv_out_data_37; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_38 = mau_3_io_pipe_phv_out_data_38; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_39 = mau_3_io_pipe_phv_out_data_39; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_40 = mau_3_io_pipe_phv_out_data_40; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_41 = mau_3_io_pipe_phv_out_data_41; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_42 = mau_3_io_pipe_phv_out_data_42; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_43 = mau_3_io_pipe_phv_out_data_43; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_44 = mau_3_io_pipe_phv_out_data_44; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_45 = mau_3_io_pipe_phv_out_data_45; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_46 = mau_3_io_pipe_phv_out_data_46; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_47 = mau_3_io_pipe_phv_out_data_47; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_48 = mau_3_io_pipe_phv_out_data_48; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_49 = mau_3_io_pipe_phv_out_data_49; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_50 = mau_3_io_pipe_phv_out_data_50; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_51 = mau_3_io_pipe_phv_out_data_51; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_52 = mau_3_io_pipe_phv_out_data_52; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_53 = mau_3_io_pipe_phv_out_data_53; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_54 = mau_3_io_pipe_phv_out_data_54; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_55 = mau_3_io_pipe_phv_out_data_55; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_56 = mau_3_io_pipe_phv_out_data_56; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_57 = mau_3_io_pipe_phv_out_data_57; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_58 = mau_3_io_pipe_phv_out_data_58; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_59 = mau_3_io_pipe_phv_out_data_59; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_60 = mau_3_io_pipe_phv_out_data_60; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_61 = mau_3_io_pipe_phv_out_data_61; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_62 = mau_3_io_pipe_phv_out_data_62; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_63 = mau_3_io_pipe_phv_out_data_63; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_64 = mau_3_io_pipe_phv_out_data_64; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_65 = mau_3_io_pipe_phv_out_data_65; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_66 = mau_3_io_pipe_phv_out_data_66; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_67 = mau_3_io_pipe_phv_out_data_67; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_68 = mau_3_io_pipe_phv_out_data_68; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_69 = mau_3_io_pipe_phv_out_data_69; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_70 = mau_3_io_pipe_phv_out_data_70; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_71 = mau_3_io_pipe_phv_out_data_71; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_72 = mau_3_io_pipe_phv_out_data_72; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_73 = mau_3_io_pipe_phv_out_data_73; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_74 = mau_3_io_pipe_phv_out_data_74; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_75 = mau_3_io_pipe_phv_out_data_75; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_76 = mau_3_io_pipe_phv_out_data_76; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_77 = mau_3_io_pipe_phv_out_data_77; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_78 = mau_3_io_pipe_phv_out_data_78; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_79 = mau_3_io_pipe_phv_out_data_79; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_80 = mau_3_io_pipe_phv_out_data_80; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_81 = mau_3_io_pipe_phv_out_data_81; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_82 = mau_3_io_pipe_phv_out_data_82; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_83 = mau_3_io_pipe_phv_out_data_83; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_84 = mau_3_io_pipe_phv_out_data_84; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_85 = mau_3_io_pipe_phv_out_data_85; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_86 = mau_3_io_pipe_phv_out_data_86; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_87 = mau_3_io_pipe_phv_out_data_87; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_88 = mau_3_io_pipe_phv_out_data_88; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_89 = mau_3_io_pipe_phv_out_data_89; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_90 = mau_3_io_pipe_phv_out_data_90; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_91 = mau_3_io_pipe_phv_out_data_91; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_92 = mau_3_io_pipe_phv_out_data_92; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_93 = mau_3_io_pipe_phv_out_data_93; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_94 = mau_3_io_pipe_phv_out_data_94; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_95 = mau_3_io_pipe_phv_out_data_95; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_96 = mau_3_io_pipe_phv_out_data_96; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_97 = mau_3_io_pipe_phv_out_data_97; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_98 = mau_3_io_pipe_phv_out_data_98; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_99 = mau_3_io_pipe_phv_out_data_99; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_100 = mau_3_io_pipe_phv_out_data_100; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_101 = mau_3_io_pipe_phv_out_data_101; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_102 = mau_3_io_pipe_phv_out_data_102; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_103 = mau_3_io_pipe_phv_out_data_103; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_104 = mau_3_io_pipe_phv_out_data_104; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_105 = mau_3_io_pipe_phv_out_data_105; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_106 = mau_3_io_pipe_phv_out_data_106; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_107 = mau_3_io_pipe_phv_out_data_107; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_108 = mau_3_io_pipe_phv_out_data_108; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_109 = mau_3_io_pipe_phv_out_data_109; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_110 = mau_3_io_pipe_phv_out_data_110; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_111 = mau_3_io_pipe_phv_out_data_111; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_112 = mau_3_io_pipe_phv_out_data_112; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_113 = mau_3_io_pipe_phv_out_data_113; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_114 = mau_3_io_pipe_phv_out_data_114; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_115 = mau_3_io_pipe_phv_out_data_115; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_116 = mau_3_io_pipe_phv_out_data_116; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_117 = mau_3_io_pipe_phv_out_data_117; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_118 = mau_3_io_pipe_phv_out_data_118; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_119 = mau_3_io_pipe_phv_out_data_119; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_120 = mau_3_io_pipe_phv_out_data_120; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_121 = mau_3_io_pipe_phv_out_data_121; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_122 = mau_3_io_pipe_phv_out_data_122; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_123 = mau_3_io_pipe_phv_out_data_123; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_124 = mau_3_io_pipe_phv_out_data_124; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_125 = mau_3_io_pipe_phv_out_data_125; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_126 = mau_3_io_pipe_phv_out_data_126; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_127 = mau_3_io_pipe_phv_out_data_127; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_128 = mau_3_io_pipe_phv_out_data_128; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_129 = mau_3_io_pipe_phv_out_data_129; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_130 = mau_3_io_pipe_phv_out_data_130; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_131 = mau_3_io_pipe_phv_out_data_131; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_132 = mau_3_io_pipe_phv_out_data_132; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_133 = mau_3_io_pipe_phv_out_data_133; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_134 = mau_3_io_pipe_phv_out_data_134; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_135 = mau_3_io_pipe_phv_out_data_135; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_136 = mau_3_io_pipe_phv_out_data_136; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_137 = mau_3_io_pipe_phv_out_data_137; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_138 = mau_3_io_pipe_phv_out_data_138; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_139 = mau_3_io_pipe_phv_out_data_139; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_140 = mau_3_io_pipe_phv_out_data_140; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_141 = mau_3_io_pipe_phv_out_data_141; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_142 = mau_3_io_pipe_phv_out_data_142; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_143 = mau_3_io_pipe_phv_out_data_143; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_144 = mau_3_io_pipe_phv_out_data_144; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_145 = mau_3_io_pipe_phv_out_data_145; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_146 = mau_3_io_pipe_phv_out_data_146; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_147 = mau_3_io_pipe_phv_out_data_147; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_148 = mau_3_io_pipe_phv_out_data_148; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_149 = mau_3_io_pipe_phv_out_data_149; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_150 = mau_3_io_pipe_phv_out_data_150; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_151 = mau_3_io_pipe_phv_out_data_151; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_152 = mau_3_io_pipe_phv_out_data_152; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_153 = mau_3_io_pipe_phv_out_data_153; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_154 = mau_3_io_pipe_phv_out_data_154; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_155 = mau_3_io_pipe_phv_out_data_155; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_156 = mau_3_io_pipe_phv_out_data_156; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_157 = mau_3_io_pipe_phv_out_data_157; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_158 = mau_3_io_pipe_phv_out_data_158; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_159 = mau_3_io_pipe_phv_out_data_159; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_160 = mau_3_io_pipe_phv_out_data_160; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_161 = mau_3_io_pipe_phv_out_data_161; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_162 = mau_3_io_pipe_phv_out_data_162; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_163 = mau_3_io_pipe_phv_out_data_163; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_164 = mau_3_io_pipe_phv_out_data_164; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_165 = mau_3_io_pipe_phv_out_data_165; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_166 = mau_3_io_pipe_phv_out_data_166; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_167 = mau_3_io_pipe_phv_out_data_167; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_168 = mau_3_io_pipe_phv_out_data_168; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_169 = mau_3_io_pipe_phv_out_data_169; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_170 = mau_3_io_pipe_phv_out_data_170; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_171 = mau_3_io_pipe_phv_out_data_171; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_172 = mau_3_io_pipe_phv_out_data_172; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_173 = mau_3_io_pipe_phv_out_data_173; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_174 = mau_3_io_pipe_phv_out_data_174; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_175 = mau_3_io_pipe_phv_out_data_175; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_176 = mau_3_io_pipe_phv_out_data_176; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_177 = mau_3_io_pipe_phv_out_data_177; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_178 = mau_3_io_pipe_phv_out_data_178; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_179 = mau_3_io_pipe_phv_out_data_179; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_180 = mau_3_io_pipe_phv_out_data_180; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_181 = mau_3_io_pipe_phv_out_data_181; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_182 = mau_3_io_pipe_phv_out_data_182; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_183 = mau_3_io_pipe_phv_out_data_183; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_184 = mau_3_io_pipe_phv_out_data_184; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_185 = mau_3_io_pipe_phv_out_data_185; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_186 = mau_3_io_pipe_phv_out_data_186; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_187 = mau_3_io_pipe_phv_out_data_187; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_188 = mau_3_io_pipe_phv_out_data_188; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_189 = mau_3_io_pipe_phv_out_data_189; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_190 = mau_3_io_pipe_phv_out_data_190; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_191 = mau_3_io_pipe_phv_out_data_191; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_192 = mau_3_io_pipe_phv_out_data_192; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_193 = mau_3_io_pipe_phv_out_data_193; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_194 = mau_3_io_pipe_phv_out_data_194; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_195 = mau_3_io_pipe_phv_out_data_195; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_196 = mau_3_io_pipe_phv_out_data_196; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_197 = mau_3_io_pipe_phv_out_data_197; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_198 = mau_3_io_pipe_phv_out_data_198; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_199 = mau_3_io_pipe_phv_out_data_199; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_200 = mau_3_io_pipe_phv_out_data_200; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_201 = mau_3_io_pipe_phv_out_data_201; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_202 = mau_3_io_pipe_phv_out_data_202; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_203 = mau_3_io_pipe_phv_out_data_203; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_204 = mau_3_io_pipe_phv_out_data_204; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_205 = mau_3_io_pipe_phv_out_data_205; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_206 = mau_3_io_pipe_phv_out_data_206; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_207 = mau_3_io_pipe_phv_out_data_207; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_208 = mau_3_io_pipe_phv_out_data_208; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_209 = mau_3_io_pipe_phv_out_data_209; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_210 = mau_3_io_pipe_phv_out_data_210; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_211 = mau_3_io_pipe_phv_out_data_211; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_212 = mau_3_io_pipe_phv_out_data_212; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_213 = mau_3_io_pipe_phv_out_data_213; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_214 = mau_3_io_pipe_phv_out_data_214; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_215 = mau_3_io_pipe_phv_out_data_215; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_216 = mau_3_io_pipe_phv_out_data_216; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_217 = mau_3_io_pipe_phv_out_data_217; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_218 = mau_3_io_pipe_phv_out_data_218; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_219 = mau_3_io_pipe_phv_out_data_219; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_220 = mau_3_io_pipe_phv_out_data_220; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_221 = mau_3_io_pipe_phv_out_data_221; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_222 = mau_3_io_pipe_phv_out_data_222; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_223 = mau_3_io_pipe_phv_out_data_223; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_224 = mau_3_io_pipe_phv_out_data_224; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_225 = mau_3_io_pipe_phv_out_data_225; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_226 = mau_3_io_pipe_phv_out_data_226; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_227 = mau_3_io_pipe_phv_out_data_227; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_228 = mau_3_io_pipe_phv_out_data_228; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_229 = mau_3_io_pipe_phv_out_data_229; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_230 = mau_3_io_pipe_phv_out_data_230; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_231 = mau_3_io_pipe_phv_out_data_231; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_232 = mau_3_io_pipe_phv_out_data_232; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_233 = mau_3_io_pipe_phv_out_data_233; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_234 = mau_3_io_pipe_phv_out_data_234; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_235 = mau_3_io_pipe_phv_out_data_235; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_236 = mau_3_io_pipe_phv_out_data_236; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_237 = mau_3_io_pipe_phv_out_data_237; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_238 = mau_3_io_pipe_phv_out_data_238; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_239 = mau_3_io_pipe_phv_out_data_239; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_240 = mau_3_io_pipe_phv_out_data_240; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_241 = mau_3_io_pipe_phv_out_data_241; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_242 = mau_3_io_pipe_phv_out_data_242; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_243 = mau_3_io_pipe_phv_out_data_243; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_244 = mau_3_io_pipe_phv_out_data_244; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_245 = mau_3_io_pipe_phv_out_data_245; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_246 = mau_3_io_pipe_phv_out_data_246; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_247 = mau_3_io_pipe_phv_out_data_247; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_248 = mau_3_io_pipe_phv_out_data_248; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_249 = mau_3_io_pipe_phv_out_data_249; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_250 = mau_3_io_pipe_phv_out_data_250; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_251 = mau_3_io_pipe_phv_out_data_251; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_252 = mau_3_io_pipe_phv_out_data_252; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_253 = mau_3_io_pipe_phv_out_data_253; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_254 = mau_3_io_pipe_phv_out_data_254; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_255 = mau_3_io_pipe_phv_out_data_255; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_256 = mau_3_io_pipe_phv_out_data_256; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_257 = mau_3_io_pipe_phv_out_data_257; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_258 = mau_3_io_pipe_phv_out_data_258; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_259 = mau_3_io_pipe_phv_out_data_259; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_260 = mau_3_io_pipe_phv_out_data_260; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_261 = mau_3_io_pipe_phv_out_data_261; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_262 = mau_3_io_pipe_phv_out_data_262; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_263 = mau_3_io_pipe_phv_out_data_263; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_264 = mau_3_io_pipe_phv_out_data_264; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_265 = mau_3_io_pipe_phv_out_data_265; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_266 = mau_3_io_pipe_phv_out_data_266; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_267 = mau_3_io_pipe_phv_out_data_267; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_268 = mau_3_io_pipe_phv_out_data_268; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_269 = mau_3_io_pipe_phv_out_data_269; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_270 = mau_3_io_pipe_phv_out_data_270; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_271 = mau_3_io_pipe_phv_out_data_271; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_272 = mau_3_io_pipe_phv_out_data_272; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_273 = mau_3_io_pipe_phv_out_data_273; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_274 = mau_3_io_pipe_phv_out_data_274; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_275 = mau_3_io_pipe_phv_out_data_275; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_276 = mau_3_io_pipe_phv_out_data_276; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_277 = mau_3_io_pipe_phv_out_data_277; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_278 = mau_3_io_pipe_phv_out_data_278; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_279 = mau_3_io_pipe_phv_out_data_279; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_280 = mau_3_io_pipe_phv_out_data_280; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_281 = mau_3_io_pipe_phv_out_data_281; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_282 = mau_3_io_pipe_phv_out_data_282; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_283 = mau_3_io_pipe_phv_out_data_283; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_284 = mau_3_io_pipe_phv_out_data_284; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_285 = mau_3_io_pipe_phv_out_data_285; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_286 = mau_3_io_pipe_phv_out_data_286; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_287 = mau_3_io_pipe_phv_out_data_287; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_288 = mau_3_io_pipe_phv_out_data_288; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_289 = mau_3_io_pipe_phv_out_data_289; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_290 = mau_3_io_pipe_phv_out_data_290; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_291 = mau_3_io_pipe_phv_out_data_291; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_292 = mau_3_io_pipe_phv_out_data_292; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_293 = mau_3_io_pipe_phv_out_data_293; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_294 = mau_3_io_pipe_phv_out_data_294; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_295 = mau_3_io_pipe_phv_out_data_295; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_296 = mau_3_io_pipe_phv_out_data_296; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_297 = mau_3_io_pipe_phv_out_data_297; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_298 = mau_3_io_pipe_phv_out_data_298; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_299 = mau_3_io_pipe_phv_out_data_299; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_300 = mau_3_io_pipe_phv_out_data_300; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_301 = mau_3_io_pipe_phv_out_data_301; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_302 = mau_3_io_pipe_phv_out_data_302; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_303 = mau_3_io_pipe_phv_out_data_303; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_304 = mau_3_io_pipe_phv_out_data_304; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_305 = mau_3_io_pipe_phv_out_data_305; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_306 = mau_3_io_pipe_phv_out_data_306; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_307 = mau_3_io_pipe_phv_out_data_307; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_308 = mau_3_io_pipe_phv_out_data_308; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_309 = mau_3_io_pipe_phv_out_data_309; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_310 = mau_3_io_pipe_phv_out_data_310; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_311 = mau_3_io_pipe_phv_out_data_311; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_312 = mau_3_io_pipe_phv_out_data_312; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_313 = mau_3_io_pipe_phv_out_data_313; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_314 = mau_3_io_pipe_phv_out_data_314; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_315 = mau_3_io_pipe_phv_out_data_315; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_316 = mau_3_io_pipe_phv_out_data_316; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_317 = mau_3_io_pipe_phv_out_data_317; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_318 = mau_3_io_pipe_phv_out_data_318; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_319 = mau_3_io_pipe_phv_out_data_319; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_320 = mau_3_io_pipe_phv_out_data_320; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_321 = mau_3_io_pipe_phv_out_data_321; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_322 = mau_3_io_pipe_phv_out_data_322; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_323 = mau_3_io_pipe_phv_out_data_323; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_324 = mau_3_io_pipe_phv_out_data_324; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_325 = mau_3_io_pipe_phv_out_data_325; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_326 = mau_3_io_pipe_phv_out_data_326; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_327 = mau_3_io_pipe_phv_out_data_327; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_328 = mau_3_io_pipe_phv_out_data_328; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_329 = mau_3_io_pipe_phv_out_data_329; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_330 = mau_3_io_pipe_phv_out_data_330; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_331 = mau_3_io_pipe_phv_out_data_331; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_332 = mau_3_io_pipe_phv_out_data_332; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_333 = mau_3_io_pipe_phv_out_data_333; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_334 = mau_3_io_pipe_phv_out_data_334; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_335 = mau_3_io_pipe_phv_out_data_335; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_336 = mau_3_io_pipe_phv_out_data_336; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_337 = mau_3_io_pipe_phv_out_data_337; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_338 = mau_3_io_pipe_phv_out_data_338; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_339 = mau_3_io_pipe_phv_out_data_339; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_340 = mau_3_io_pipe_phv_out_data_340; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_341 = mau_3_io_pipe_phv_out_data_341; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_342 = mau_3_io_pipe_phv_out_data_342; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_343 = mau_3_io_pipe_phv_out_data_343; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_344 = mau_3_io_pipe_phv_out_data_344; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_345 = mau_3_io_pipe_phv_out_data_345; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_346 = mau_3_io_pipe_phv_out_data_346; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_347 = mau_3_io_pipe_phv_out_data_347; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_348 = mau_3_io_pipe_phv_out_data_348; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_349 = mau_3_io_pipe_phv_out_data_349; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_350 = mau_3_io_pipe_phv_out_data_350; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_351 = mau_3_io_pipe_phv_out_data_351; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_352 = mau_3_io_pipe_phv_out_data_352; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_353 = mau_3_io_pipe_phv_out_data_353; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_354 = mau_3_io_pipe_phv_out_data_354; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_355 = mau_3_io_pipe_phv_out_data_355; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_356 = mau_3_io_pipe_phv_out_data_356; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_357 = mau_3_io_pipe_phv_out_data_357; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_358 = mau_3_io_pipe_phv_out_data_358; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_359 = mau_3_io_pipe_phv_out_data_359; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_360 = mau_3_io_pipe_phv_out_data_360; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_361 = mau_3_io_pipe_phv_out_data_361; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_362 = mau_3_io_pipe_phv_out_data_362; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_363 = mau_3_io_pipe_phv_out_data_363; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_364 = mau_3_io_pipe_phv_out_data_364; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_365 = mau_3_io_pipe_phv_out_data_365; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_366 = mau_3_io_pipe_phv_out_data_366; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_367 = mau_3_io_pipe_phv_out_data_367; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_368 = mau_3_io_pipe_phv_out_data_368; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_369 = mau_3_io_pipe_phv_out_data_369; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_370 = mau_3_io_pipe_phv_out_data_370; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_371 = mau_3_io_pipe_phv_out_data_371; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_372 = mau_3_io_pipe_phv_out_data_372; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_373 = mau_3_io_pipe_phv_out_data_373; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_374 = mau_3_io_pipe_phv_out_data_374; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_375 = mau_3_io_pipe_phv_out_data_375; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_376 = mau_3_io_pipe_phv_out_data_376; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_377 = mau_3_io_pipe_phv_out_data_377; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_378 = mau_3_io_pipe_phv_out_data_378; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_379 = mau_3_io_pipe_phv_out_data_379; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_380 = mau_3_io_pipe_phv_out_data_380; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_381 = mau_3_io_pipe_phv_out_data_381; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_382 = mau_3_io_pipe_phv_out_data_382; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_383 = mau_3_io_pipe_phv_out_data_383; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_384 = mau_3_io_pipe_phv_out_data_384; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_385 = mau_3_io_pipe_phv_out_data_385; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_386 = mau_3_io_pipe_phv_out_data_386; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_387 = mau_3_io_pipe_phv_out_data_387; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_388 = mau_3_io_pipe_phv_out_data_388; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_389 = mau_3_io_pipe_phv_out_data_389; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_390 = mau_3_io_pipe_phv_out_data_390; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_391 = mau_3_io_pipe_phv_out_data_391; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_392 = mau_3_io_pipe_phv_out_data_392; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_393 = mau_3_io_pipe_phv_out_data_393; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_394 = mau_3_io_pipe_phv_out_data_394; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_395 = mau_3_io_pipe_phv_out_data_395; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_396 = mau_3_io_pipe_phv_out_data_396; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_397 = mau_3_io_pipe_phv_out_data_397; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_398 = mau_3_io_pipe_phv_out_data_398; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_399 = mau_3_io_pipe_phv_out_data_399; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_400 = mau_3_io_pipe_phv_out_data_400; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_401 = mau_3_io_pipe_phv_out_data_401; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_402 = mau_3_io_pipe_phv_out_data_402; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_403 = mau_3_io_pipe_phv_out_data_403; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_404 = mau_3_io_pipe_phv_out_data_404; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_405 = mau_3_io_pipe_phv_out_data_405; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_406 = mau_3_io_pipe_phv_out_data_406; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_407 = mau_3_io_pipe_phv_out_data_407; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_408 = mau_3_io_pipe_phv_out_data_408; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_409 = mau_3_io_pipe_phv_out_data_409; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_410 = mau_3_io_pipe_phv_out_data_410; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_411 = mau_3_io_pipe_phv_out_data_411; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_412 = mau_3_io_pipe_phv_out_data_412; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_413 = mau_3_io_pipe_phv_out_data_413; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_414 = mau_3_io_pipe_phv_out_data_414; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_415 = mau_3_io_pipe_phv_out_data_415; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_416 = mau_3_io_pipe_phv_out_data_416; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_417 = mau_3_io_pipe_phv_out_data_417; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_418 = mau_3_io_pipe_phv_out_data_418; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_419 = mau_3_io_pipe_phv_out_data_419; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_420 = mau_3_io_pipe_phv_out_data_420; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_421 = mau_3_io_pipe_phv_out_data_421; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_422 = mau_3_io_pipe_phv_out_data_422; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_423 = mau_3_io_pipe_phv_out_data_423; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_424 = mau_3_io_pipe_phv_out_data_424; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_425 = mau_3_io_pipe_phv_out_data_425; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_426 = mau_3_io_pipe_phv_out_data_426; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_427 = mau_3_io_pipe_phv_out_data_427; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_428 = mau_3_io_pipe_phv_out_data_428; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_429 = mau_3_io_pipe_phv_out_data_429; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_430 = mau_3_io_pipe_phv_out_data_430; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_431 = mau_3_io_pipe_phv_out_data_431; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_432 = mau_3_io_pipe_phv_out_data_432; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_433 = mau_3_io_pipe_phv_out_data_433; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_434 = mau_3_io_pipe_phv_out_data_434; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_435 = mau_3_io_pipe_phv_out_data_435; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_436 = mau_3_io_pipe_phv_out_data_436; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_437 = mau_3_io_pipe_phv_out_data_437; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_438 = mau_3_io_pipe_phv_out_data_438; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_439 = mau_3_io_pipe_phv_out_data_439; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_440 = mau_3_io_pipe_phv_out_data_440; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_441 = mau_3_io_pipe_phv_out_data_441; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_442 = mau_3_io_pipe_phv_out_data_442; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_443 = mau_3_io_pipe_phv_out_data_443; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_444 = mau_3_io_pipe_phv_out_data_444; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_445 = mau_3_io_pipe_phv_out_data_445; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_446 = mau_3_io_pipe_phv_out_data_446; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_447 = mau_3_io_pipe_phv_out_data_447; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_448 = mau_3_io_pipe_phv_out_data_448; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_449 = mau_3_io_pipe_phv_out_data_449; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_450 = mau_3_io_pipe_phv_out_data_450; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_451 = mau_3_io_pipe_phv_out_data_451; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_452 = mau_3_io_pipe_phv_out_data_452; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_453 = mau_3_io_pipe_phv_out_data_453; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_454 = mau_3_io_pipe_phv_out_data_454; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_455 = mau_3_io_pipe_phv_out_data_455; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_456 = mau_3_io_pipe_phv_out_data_456; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_457 = mau_3_io_pipe_phv_out_data_457; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_458 = mau_3_io_pipe_phv_out_data_458; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_459 = mau_3_io_pipe_phv_out_data_459; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_460 = mau_3_io_pipe_phv_out_data_460; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_461 = mau_3_io_pipe_phv_out_data_461; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_462 = mau_3_io_pipe_phv_out_data_462; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_463 = mau_3_io_pipe_phv_out_data_463; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_464 = mau_3_io_pipe_phv_out_data_464; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_465 = mau_3_io_pipe_phv_out_data_465; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_466 = mau_3_io_pipe_phv_out_data_466; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_467 = mau_3_io_pipe_phv_out_data_467; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_468 = mau_3_io_pipe_phv_out_data_468; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_469 = mau_3_io_pipe_phv_out_data_469; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_470 = mau_3_io_pipe_phv_out_data_470; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_471 = mau_3_io_pipe_phv_out_data_471; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_472 = mau_3_io_pipe_phv_out_data_472; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_473 = mau_3_io_pipe_phv_out_data_473; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_474 = mau_3_io_pipe_phv_out_data_474; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_475 = mau_3_io_pipe_phv_out_data_475; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_476 = mau_3_io_pipe_phv_out_data_476; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_477 = mau_3_io_pipe_phv_out_data_477; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_478 = mau_3_io_pipe_phv_out_data_478; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_479 = mau_3_io_pipe_phv_out_data_479; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_480 = mau_3_io_pipe_phv_out_data_480; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_481 = mau_3_io_pipe_phv_out_data_481; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_482 = mau_3_io_pipe_phv_out_data_482; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_483 = mau_3_io_pipe_phv_out_data_483; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_484 = mau_3_io_pipe_phv_out_data_484; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_485 = mau_3_io_pipe_phv_out_data_485; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_486 = mau_3_io_pipe_phv_out_data_486; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_487 = mau_3_io_pipe_phv_out_data_487; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_488 = mau_3_io_pipe_phv_out_data_488; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_489 = mau_3_io_pipe_phv_out_data_489; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_490 = mau_3_io_pipe_phv_out_data_490; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_491 = mau_3_io_pipe_phv_out_data_491; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_492 = mau_3_io_pipe_phv_out_data_492; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_493 = mau_3_io_pipe_phv_out_data_493; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_494 = mau_3_io_pipe_phv_out_data_494; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_495 = mau_3_io_pipe_phv_out_data_495; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_496 = mau_3_io_pipe_phv_out_data_496; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_497 = mau_3_io_pipe_phv_out_data_497; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_498 = mau_3_io_pipe_phv_out_data_498; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_499 = mau_3_io_pipe_phv_out_data_499; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_500 = mau_3_io_pipe_phv_out_data_500; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_501 = mau_3_io_pipe_phv_out_data_501; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_502 = mau_3_io_pipe_phv_out_data_502; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_503 = mau_3_io_pipe_phv_out_data_503; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_504 = mau_3_io_pipe_phv_out_data_504; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_505 = mau_3_io_pipe_phv_out_data_505; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_506 = mau_3_io_pipe_phv_out_data_506; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_507 = mau_3_io_pipe_phv_out_data_507; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_508 = mau_3_io_pipe_phv_out_data_508; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_509 = mau_3_io_pipe_phv_out_data_509; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_510 = mau_3_io_pipe_phv_out_data_510; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_511 = mau_3_io_pipe_phv_out_data_511; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_header_0 = mau_3_io_pipe_phv_out_header_0; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_header_1 = mau_3_io_pipe_phv_out_header_1; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_header_2 = mau_3_io_pipe_phv_out_header_2; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_header_3 = mau_3_io_pipe_phv_out_header_3; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_header_4 = mau_3_io_pipe_phv_out_header_4; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_header_5 = mau_3_io_pipe_phv_out_header_5; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_header_6 = mau_3_io_pipe_phv_out_header_6; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_header_7 = mau_3_io_pipe_phv_out_header_7; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_header_8 = mau_3_io_pipe_phv_out_header_8; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_header_9 = mau_3_io_pipe_phv_out_header_9; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_header_10 = mau_3_io_pipe_phv_out_header_10; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_header_11 = mau_3_io_pipe_phv_out_header_11; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_header_12 = mau_3_io_pipe_phv_out_header_12; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_header_13 = mau_3_io_pipe_phv_out_header_13; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_header_14 = mau_3_io_pipe_phv_out_header_14; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_header_15 = mau_3_io_pipe_phv_out_header_15; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_parse_current_state = mau_3_io_pipe_phv_out_parse_current_state; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_parse_current_offset = mau_3_io_pipe_phv_out_parse_current_offset; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_parse_transition_field = mau_3_io_pipe_phv_out_parse_transition_field; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_next_processor_id = mau_3_io_pipe_phv_out_next_processor_id; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_next_config_id = mau_3_io_pipe_phv_out_next_config_id; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_is_valid_processor = mau_3_io_pipe_phv_out_is_valid_processor; // @[parser_pisa.scala 42:35]
  assign mau_4_io_mod_state_id_mod = io_mod_en ? io_mod_module_mod_state_id_mod & mod_j_4 :
    io_mod_module_mod_state_id_mod; // @[parser_pisa.scala 51:22 parser_pisa.scala 58:40 parser_pisa.scala 47:23]
  assign mau_4_io_mod_state_id = io_mod_module_mod_state_id; // @[parser_pisa.scala 47:23]
  assign mau_4_io_mod_sram_w_cs = io_mod_module_mod_sram_w_cs; // @[parser_pisa.scala 47:23]
  assign mau_4_io_mod_sram_w_en = io_mod_en ? io_mod_module_mod_sram_w_en & mod_j_4 : io_mod_module_mod_sram_w_en; // @[parser_pisa.scala 51:22 parser_pisa.scala 57:40 parser_pisa.scala 47:23]
  assign mau_4_io_mod_sram_w_addr = io_mod_module_mod_sram_w_addr; // @[parser_pisa.scala 47:23]
  assign mau_4_io_mod_sram_w_data = io_mod_module_mod_sram_w_data; // @[parser_pisa.scala 47:23]
  assign mau_5_clock = clock;
  assign mau_5_io_pipe_phv_in_data_0 = mau_4_io_pipe_phv_out_data_0; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_1 = mau_4_io_pipe_phv_out_data_1; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_2 = mau_4_io_pipe_phv_out_data_2; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_3 = mau_4_io_pipe_phv_out_data_3; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_4 = mau_4_io_pipe_phv_out_data_4; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_5 = mau_4_io_pipe_phv_out_data_5; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_6 = mau_4_io_pipe_phv_out_data_6; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_7 = mau_4_io_pipe_phv_out_data_7; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_8 = mau_4_io_pipe_phv_out_data_8; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_9 = mau_4_io_pipe_phv_out_data_9; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_10 = mau_4_io_pipe_phv_out_data_10; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_11 = mau_4_io_pipe_phv_out_data_11; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_12 = mau_4_io_pipe_phv_out_data_12; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_13 = mau_4_io_pipe_phv_out_data_13; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_14 = mau_4_io_pipe_phv_out_data_14; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_15 = mau_4_io_pipe_phv_out_data_15; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_16 = mau_4_io_pipe_phv_out_data_16; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_17 = mau_4_io_pipe_phv_out_data_17; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_18 = mau_4_io_pipe_phv_out_data_18; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_19 = mau_4_io_pipe_phv_out_data_19; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_20 = mau_4_io_pipe_phv_out_data_20; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_21 = mau_4_io_pipe_phv_out_data_21; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_22 = mau_4_io_pipe_phv_out_data_22; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_23 = mau_4_io_pipe_phv_out_data_23; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_24 = mau_4_io_pipe_phv_out_data_24; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_25 = mau_4_io_pipe_phv_out_data_25; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_26 = mau_4_io_pipe_phv_out_data_26; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_27 = mau_4_io_pipe_phv_out_data_27; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_28 = mau_4_io_pipe_phv_out_data_28; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_29 = mau_4_io_pipe_phv_out_data_29; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_30 = mau_4_io_pipe_phv_out_data_30; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_31 = mau_4_io_pipe_phv_out_data_31; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_32 = mau_4_io_pipe_phv_out_data_32; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_33 = mau_4_io_pipe_phv_out_data_33; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_34 = mau_4_io_pipe_phv_out_data_34; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_35 = mau_4_io_pipe_phv_out_data_35; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_36 = mau_4_io_pipe_phv_out_data_36; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_37 = mau_4_io_pipe_phv_out_data_37; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_38 = mau_4_io_pipe_phv_out_data_38; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_39 = mau_4_io_pipe_phv_out_data_39; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_40 = mau_4_io_pipe_phv_out_data_40; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_41 = mau_4_io_pipe_phv_out_data_41; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_42 = mau_4_io_pipe_phv_out_data_42; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_43 = mau_4_io_pipe_phv_out_data_43; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_44 = mau_4_io_pipe_phv_out_data_44; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_45 = mau_4_io_pipe_phv_out_data_45; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_46 = mau_4_io_pipe_phv_out_data_46; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_47 = mau_4_io_pipe_phv_out_data_47; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_48 = mau_4_io_pipe_phv_out_data_48; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_49 = mau_4_io_pipe_phv_out_data_49; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_50 = mau_4_io_pipe_phv_out_data_50; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_51 = mau_4_io_pipe_phv_out_data_51; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_52 = mau_4_io_pipe_phv_out_data_52; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_53 = mau_4_io_pipe_phv_out_data_53; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_54 = mau_4_io_pipe_phv_out_data_54; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_55 = mau_4_io_pipe_phv_out_data_55; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_56 = mau_4_io_pipe_phv_out_data_56; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_57 = mau_4_io_pipe_phv_out_data_57; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_58 = mau_4_io_pipe_phv_out_data_58; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_59 = mau_4_io_pipe_phv_out_data_59; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_60 = mau_4_io_pipe_phv_out_data_60; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_61 = mau_4_io_pipe_phv_out_data_61; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_62 = mau_4_io_pipe_phv_out_data_62; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_63 = mau_4_io_pipe_phv_out_data_63; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_64 = mau_4_io_pipe_phv_out_data_64; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_65 = mau_4_io_pipe_phv_out_data_65; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_66 = mau_4_io_pipe_phv_out_data_66; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_67 = mau_4_io_pipe_phv_out_data_67; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_68 = mau_4_io_pipe_phv_out_data_68; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_69 = mau_4_io_pipe_phv_out_data_69; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_70 = mau_4_io_pipe_phv_out_data_70; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_71 = mau_4_io_pipe_phv_out_data_71; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_72 = mau_4_io_pipe_phv_out_data_72; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_73 = mau_4_io_pipe_phv_out_data_73; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_74 = mau_4_io_pipe_phv_out_data_74; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_75 = mau_4_io_pipe_phv_out_data_75; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_76 = mau_4_io_pipe_phv_out_data_76; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_77 = mau_4_io_pipe_phv_out_data_77; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_78 = mau_4_io_pipe_phv_out_data_78; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_79 = mau_4_io_pipe_phv_out_data_79; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_80 = mau_4_io_pipe_phv_out_data_80; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_81 = mau_4_io_pipe_phv_out_data_81; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_82 = mau_4_io_pipe_phv_out_data_82; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_83 = mau_4_io_pipe_phv_out_data_83; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_84 = mau_4_io_pipe_phv_out_data_84; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_85 = mau_4_io_pipe_phv_out_data_85; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_86 = mau_4_io_pipe_phv_out_data_86; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_87 = mau_4_io_pipe_phv_out_data_87; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_88 = mau_4_io_pipe_phv_out_data_88; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_89 = mau_4_io_pipe_phv_out_data_89; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_90 = mau_4_io_pipe_phv_out_data_90; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_91 = mau_4_io_pipe_phv_out_data_91; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_92 = mau_4_io_pipe_phv_out_data_92; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_93 = mau_4_io_pipe_phv_out_data_93; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_94 = mau_4_io_pipe_phv_out_data_94; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_95 = mau_4_io_pipe_phv_out_data_95; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_96 = mau_4_io_pipe_phv_out_data_96; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_97 = mau_4_io_pipe_phv_out_data_97; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_98 = mau_4_io_pipe_phv_out_data_98; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_99 = mau_4_io_pipe_phv_out_data_99; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_100 = mau_4_io_pipe_phv_out_data_100; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_101 = mau_4_io_pipe_phv_out_data_101; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_102 = mau_4_io_pipe_phv_out_data_102; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_103 = mau_4_io_pipe_phv_out_data_103; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_104 = mau_4_io_pipe_phv_out_data_104; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_105 = mau_4_io_pipe_phv_out_data_105; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_106 = mau_4_io_pipe_phv_out_data_106; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_107 = mau_4_io_pipe_phv_out_data_107; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_108 = mau_4_io_pipe_phv_out_data_108; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_109 = mau_4_io_pipe_phv_out_data_109; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_110 = mau_4_io_pipe_phv_out_data_110; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_111 = mau_4_io_pipe_phv_out_data_111; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_112 = mau_4_io_pipe_phv_out_data_112; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_113 = mau_4_io_pipe_phv_out_data_113; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_114 = mau_4_io_pipe_phv_out_data_114; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_115 = mau_4_io_pipe_phv_out_data_115; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_116 = mau_4_io_pipe_phv_out_data_116; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_117 = mau_4_io_pipe_phv_out_data_117; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_118 = mau_4_io_pipe_phv_out_data_118; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_119 = mau_4_io_pipe_phv_out_data_119; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_120 = mau_4_io_pipe_phv_out_data_120; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_121 = mau_4_io_pipe_phv_out_data_121; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_122 = mau_4_io_pipe_phv_out_data_122; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_123 = mau_4_io_pipe_phv_out_data_123; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_124 = mau_4_io_pipe_phv_out_data_124; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_125 = mau_4_io_pipe_phv_out_data_125; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_126 = mau_4_io_pipe_phv_out_data_126; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_127 = mau_4_io_pipe_phv_out_data_127; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_128 = mau_4_io_pipe_phv_out_data_128; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_129 = mau_4_io_pipe_phv_out_data_129; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_130 = mau_4_io_pipe_phv_out_data_130; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_131 = mau_4_io_pipe_phv_out_data_131; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_132 = mau_4_io_pipe_phv_out_data_132; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_133 = mau_4_io_pipe_phv_out_data_133; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_134 = mau_4_io_pipe_phv_out_data_134; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_135 = mau_4_io_pipe_phv_out_data_135; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_136 = mau_4_io_pipe_phv_out_data_136; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_137 = mau_4_io_pipe_phv_out_data_137; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_138 = mau_4_io_pipe_phv_out_data_138; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_139 = mau_4_io_pipe_phv_out_data_139; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_140 = mau_4_io_pipe_phv_out_data_140; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_141 = mau_4_io_pipe_phv_out_data_141; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_142 = mau_4_io_pipe_phv_out_data_142; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_143 = mau_4_io_pipe_phv_out_data_143; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_144 = mau_4_io_pipe_phv_out_data_144; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_145 = mau_4_io_pipe_phv_out_data_145; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_146 = mau_4_io_pipe_phv_out_data_146; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_147 = mau_4_io_pipe_phv_out_data_147; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_148 = mau_4_io_pipe_phv_out_data_148; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_149 = mau_4_io_pipe_phv_out_data_149; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_150 = mau_4_io_pipe_phv_out_data_150; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_151 = mau_4_io_pipe_phv_out_data_151; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_152 = mau_4_io_pipe_phv_out_data_152; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_153 = mau_4_io_pipe_phv_out_data_153; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_154 = mau_4_io_pipe_phv_out_data_154; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_155 = mau_4_io_pipe_phv_out_data_155; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_156 = mau_4_io_pipe_phv_out_data_156; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_157 = mau_4_io_pipe_phv_out_data_157; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_158 = mau_4_io_pipe_phv_out_data_158; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_159 = mau_4_io_pipe_phv_out_data_159; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_160 = mau_4_io_pipe_phv_out_data_160; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_161 = mau_4_io_pipe_phv_out_data_161; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_162 = mau_4_io_pipe_phv_out_data_162; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_163 = mau_4_io_pipe_phv_out_data_163; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_164 = mau_4_io_pipe_phv_out_data_164; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_165 = mau_4_io_pipe_phv_out_data_165; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_166 = mau_4_io_pipe_phv_out_data_166; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_167 = mau_4_io_pipe_phv_out_data_167; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_168 = mau_4_io_pipe_phv_out_data_168; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_169 = mau_4_io_pipe_phv_out_data_169; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_170 = mau_4_io_pipe_phv_out_data_170; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_171 = mau_4_io_pipe_phv_out_data_171; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_172 = mau_4_io_pipe_phv_out_data_172; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_173 = mau_4_io_pipe_phv_out_data_173; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_174 = mau_4_io_pipe_phv_out_data_174; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_175 = mau_4_io_pipe_phv_out_data_175; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_176 = mau_4_io_pipe_phv_out_data_176; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_177 = mau_4_io_pipe_phv_out_data_177; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_178 = mau_4_io_pipe_phv_out_data_178; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_179 = mau_4_io_pipe_phv_out_data_179; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_180 = mau_4_io_pipe_phv_out_data_180; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_181 = mau_4_io_pipe_phv_out_data_181; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_182 = mau_4_io_pipe_phv_out_data_182; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_183 = mau_4_io_pipe_phv_out_data_183; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_184 = mau_4_io_pipe_phv_out_data_184; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_185 = mau_4_io_pipe_phv_out_data_185; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_186 = mau_4_io_pipe_phv_out_data_186; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_187 = mau_4_io_pipe_phv_out_data_187; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_188 = mau_4_io_pipe_phv_out_data_188; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_189 = mau_4_io_pipe_phv_out_data_189; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_190 = mau_4_io_pipe_phv_out_data_190; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_191 = mau_4_io_pipe_phv_out_data_191; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_192 = mau_4_io_pipe_phv_out_data_192; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_193 = mau_4_io_pipe_phv_out_data_193; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_194 = mau_4_io_pipe_phv_out_data_194; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_195 = mau_4_io_pipe_phv_out_data_195; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_196 = mau_4_io_pipe_phv_out_data_196; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_197 = mau_4_io_pipe_phv_out_data_197; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_198 = mau_4_io_pipe_phv_out_data_198; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_199 = mau_4_io_pipe_phv_out_data_199; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_200 = mau_4_io_pipe_phv_out_data_200; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_201 = mau_4_io_pipe_phv_out_data_201; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_202 = mau_4_io_pipe_phv_out_data_202; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_203 = mau_4_io_pipe_phv_out_data_203; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_204 = mau_4_io_pipe_phv_out_data_204; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_205 = mau_4_io_pipe_phv_out_data_205; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_206 = mau_4_io_pipe_phv_out_data_206; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_207 = mau_4_io_pipe_phv_out_data_207; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_208 = mau_4_io_pipe_phv_out_data_208; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_209 = mau_4_io_pipe_phv_out_data_209; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_210 = mau_4_io_pipe_phv_out_data_210; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_211 = mau_4_io_pipe_phv_out_data_211; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_212 = mau_4_io_pipe_phv_out_data_212; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_213 = mau_4_io_pipe_phv_out_data_213; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_214 = mau_4_io_pipe_phv_out_data_214; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_215 = mau_4_io_pipe_phv_out_data_215; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_216 = mau_4_io_pipe_phv_out_data_216; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_217 = mau_4_io_pipe_phv_out_data_217; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_218 = mau_4_io_pipe_phv_out_data_218; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_219 = mau_4_io_pipe_phv_out_data_219; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_220 = mau_4_io_pipe_phv_out_data_220; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_221 = mau_4_io_pipe_phv_out_data_221; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_222 = mau_4_io_pipe_phv_out_data_222; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_223 = mau_4_io_pipe_phv_out_data_223; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_224 = mau_4_io_pipe_phv_out_data_224; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_225 = mau_4_io_pipe_phv_out_data_225; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_226 = mau_4_io_pipe_phv_out_data_226; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_227 = mau_4_io_pipe_phv_out_data_227; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_228 = mau_4_io_pipe_phv_out_data_228; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_229 = mau_4_io_pipe_phv_out_data_229; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_230 = mau_4_io_pipe_phv_out_data_230; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_231 = mau_4_io_pipe_phv_out_data_231; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_232 = mau_4_io_pipe_phv_out_data_232; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_233 = mau_4_io_pipe_phv_out_data_233; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_234 = mau_4_io_pipe_phv_out_data_234; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_235 = mau_4_io_pipe_phv_out_data_235; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_236 = mau_4_io_pipe_phv_out_data_236; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_237 = mau_4_io_pipe_phv_out_data_237; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_238 = mau_4_io_pipe_phv_out_data_238; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_239 = mau_4_io_pipe_phv_out_data_239; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_240 = mau_4_io_pipe_phv_out_data_240; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_241 = mau_4_io_pipe_phv_out_data_241; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_242 = mau_4_io_pipe_phv_out_data_242; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_243 = mau_4_io_pipe_phv_out_data_243; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_244 = mau_4_io_pipe_phv_out_data_244; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_245 = mau_4_io_pipe_phv_out_data_245; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_246 = mau_4_io_pipe_phv_out_data_246; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_247 = mau_4_io_pipe_phv_out_data_247; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_248 = mau_4_io_pipe_phv_out_data_248; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_249 = mau_4_io_pipe_phv_out_data_249; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_250 = mau_4_io_pipe_phv_out_data_250; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_251 = mau_4_io_pipe_phv_out_data_251; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_252 = mau_4_io_pipe_phv_out_data_252; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_253 = mau_4_io_pipe_phv_out_data_253; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_254 = mau_4_io_pipe_phv_out_data_254; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_255 = mau_4_io_pipe_phv_out_data_255; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_256 = mau_4_io_pipe_phv_out_data_256; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_257 = mau_4_io_pipe_phv_out_data_257; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_258 = mau_4_io_pipe_phv_out_data_258; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_259 = mau_4_io_pipe_phv_out_data_259; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_260 = mau_4_io_pipe_phv_out_data_260; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_261 = mau_4_io_pipe_phv_out_data_261; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_262 = mau_4_io_pipe_phv_out_data_262; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_263 = mau_4_io_pipe_phv_out_data_263; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_264 = mau_4_io_pipe_phv_out_data_264; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_265 = mau_4_io_pipe_phv_out_data_265; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_266 = mau_4_io_pipe_phv_out_data_266; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_267 = mau_4_io_pipe_phv_out_data_267; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_268 = mau_4_io_pipe_phv_out_data_268; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_269 = mau_4_io_pipe_phv_out_data_269; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_270 = mau_4_io_pipe_phv_out_data_270; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_271 = mau_4_io_pipe_phv_out_data_271; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_272 = mau_4_io_pipe_phv_out_data_272; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_273 = mau_4_io_pipe_phv_out_data_273; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_274 = mau_4_io_pipe_phv_out_data_274; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_275 = mau_4_io_pipe_phv_out_data_275; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_276 = mau_4_io_pipe_phv_out_data_276; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_277 = mau_4_io_pipe_phv_out_data_277; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_278 = mau_4_io_pipe_phv_out_data_278; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_279 = mau_4_io_pipe_phv_out_data_279; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_280 = mau_4_io_pipe_phv_out_data_280; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_281 = mau_4_io_pipe_phv_out_data_281; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_282 = mau_4_io_pipe_phv_out_data_282; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_283 = mau_4_io_pipe_phv_out_data_283; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_284 = mau_4_io_pipe_phv_out_data_284; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_285 = mau_4_io_pipe_phv_out_data_285; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_286 = mau_4_io_pipe_phv_out_data_286; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_287 = mau_4_io_pipe_phv_out_data_287; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_288 = mau_4_io_pipe_phv_out_data_288; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_289 = mau_4_io_pipe_phv_out_data_289; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_290 = mau_4_io_pipe_phv_out_data_290; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_291 = mau_4_io_pipe_phv_out_data_291; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_292 = mau_4_io_pipe_phv_out_data_292; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_293 = mau_4_io_pipe_phv_out_data_293; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_294 = mau_4_io_pipe_phv_out_data_294; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_295 = mau_4_io_pipe_phv_out_data_295; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_296 = mau_4_io_pipe_phv_out_data_296; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_297 = mau_4_io_pipe_phv_out_data_297; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_298 = mau_4_io_pipe_phv_out_data_298; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_299 = mau_4_io_pipe_phv_out_data_299; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_300 = mau_4_io_pipe_phv_out_data_300; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_301 = mau_4_io_pipe_phv_out_data_301; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_302 = mau_4_io_pipe_phv_out_data_302; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_303 = mau_4_io_pipe_phv_out_data_303; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_304 = mau_4_io_pipe_phv_out_data_304; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_305 = mau_4_io_pipe_phv_out_data_305; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_306 = mau_4_io_pipe_phv_out_data_306; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_307 = mau_4_io_pipe_phv_out_data_307; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_308 = mau_4_io_pipe_phv_out_data_308; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_309 = mau_4_io_pipe_phv_out_data_309; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_310 = mau_4_io_pipe_phv_out_data_310; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_311 = mau_4_io_pipe_phv_out_data_311; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_312 = mau_4_io_pipe_phv_out_data_312; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_313 = mau_4_io_pipe_phv_out_data_313; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_314 = mau_4_io_pipe_phv_out_data_314; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_315 = mau_4_io_pipe_phv_out_data_315; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_316 = mau_4_io_pipe_phv_out_data_316; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_317 = mau_4_io_pipe_phv_out_data_317; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_318 = mau_4_io_pipe_phv_out_data_318; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_319 = mau_4_io_pipe_phv_out_data_319; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_320 = mau_4_io_pipe_phv_out_data_320; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_321 = mau_4_io_pipe_phv_out_data_321; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_322 = mau_4_io_pipe_phv_out_data_322; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_323 = mau_4_io_pipe_phv_out_data_323; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_324 = mau_4_io_pipe_phv_out_data_324; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_325 = mau_4_io_pipe_phv_out_data_325; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_326 = mau_4_io_pipe_phv_out_data_326; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_327 = mau_4_io_pipe_phv_out_data_327; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_328 = mau_4_io_pipe_phv_out_data_328; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_329 = mau_4_io_pipe_phv_out_data_329; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_330 = mau_4_io_pipe_phv_out_data_330; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_331 = mau_4_io_pipe_phv_out_data_331; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_332 = mau_4_io_pipe_phv_out_data_332; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_333 = mau_4_io_pipe_phv_out_data_333; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_334 = mau_4_io_pipe_phv_out_data_334; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_335 = mau_4_io_pipe_phv_out_data_335; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_336 = mau_4_io_pipe_phv_out_data_336; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_337 = mau_4_io_pipe_phv_out_data_337; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_338 = mau_4_io_pipe_phv_out_data_338; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_339 = mau_4_io_pipe_phv_out_data_339; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_340 = mau_4_io_pipe_phv_out_data_340; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_341 = mau_4_io_pipe_phv_out_data_341; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_342 = mau_4_io_pipe_phv_out_data_342; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_343 = mau_4_io_pipe_phv_out_data_343; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_344 = mau_4_io_pipe_phv_out_data_344; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_345 = mau_4_io_pipe_phv_out_data_345; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_346 = mau_4_io_pipe_phv_out_data_346; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_347 = mau_4_io_pipe_phv_out_data_347; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_348 = mau_4_io_pipe_phv_out_data_348; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_349 = mau_4_io_pipe_phv_out_data_349; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_350 = mau_4_io_pipe_phv_out_data_350; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_351 = mau_4_io_pipe_phv_out_data_351; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_352 = mau_4_io_pipe_phv_out_data_352; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_353 = mau_4_io_pipe_phv_out_data_353; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_354 = mau_4_io_pipe_phv_out_data_354; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_355 = mau_4_io_pipe_phv_out_data_355; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_356 = mau_4_io_pipe_phv_out_data_356; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_357 = mau_4_io_pipe_phv_out_data_357; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_358 = mau_4_io_pipe_phv_out_data_358; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_359 = mau_4_io_pipe_phv_out_data_359; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_360 = mau_4_io_pipe_phv_out_data_360; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_361 = mau_4_io_pipe_phv_out_data_361; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_362 = mau_4_io_pipe_phv_out_data_362; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_363 = mau_4_io_pipe_phv_out_data_363; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_364 = mau_4_io_pipe_phv_out_data_364; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_365 = mau_4_io_pipe_phv_out_data_365; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_366 = mau_4_io_pipe_phv_out_data_366; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_367 = mau_4_io_pipe_phv_out_data_367; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_368 = mau_4_io_pipe_phv_out_data_368; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_369 = mau_4_io_pipe_phv_out_data_369; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_370 = mau_4_io_pipe_phv_out_data_370; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_371 = mau_4_io_pipe_phv_out_data_371; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_372 = mau_4_io_pipe_phv_out_data_372; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_373 = mau_4_io_pipe_phv_out_data_373; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_374 = mau_4_io_pipe_phv_out_data_374; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_375 = mau_4_io_pipe_phv_out_data_375; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_376 = mau_4_io_pipe_phv_out_data_376; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_377 = mau_4_io_pipe_phv_out_data_377; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_378 = mau_4_io_pipe_phv_out_data_378; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_379 = mau_4_io_pipe_phv_out_data_379; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_380 = mau_4_io_pipe_phv_out_data_380; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_381 = mau_4_io_pipe_phv_out_data_381; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_382 = mau_4_io_pipe_phv_out_data_382; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_383 = mau_4_io_pipe_phv_out_data_383; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_384 = mau_4_io_pipe_phv_out_data_384; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_385 = mau_4_io_pipe_phv_out_data_385; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_386 = mau_4_io_pipe_phv_out_data_386; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_387 = mau_4_io_pipe_phv_out_data_387; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_388 = mau_4_io_pipe_phv_out_data_388; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_389 = mau_4_io_pipe_phv_out_data_389; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_390 = mau_4_io_pipe_phv_out_data_390; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_391 = mau_4_io_pipe_phv_out_data_391; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_392 = mau_4_io_pipe_phv_out_data_392; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_393 = mau_4_io_pipe_phv_out_data_393; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_394 = mau_4_io_pipe_phv_out_data_394; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_395 = mau_4_io_pipe_phv_out_data_395; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_396 = mau_4_io_pipe_phv_out_data_396; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_397 = mau_4_io_pipe_phv_out_data_397; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_398 = mau_4_io_pipe_phv_out_data_398; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_399 = mau_4_io_pipe_phv_out_data_399; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_400 = mau_4_io_pipe_phv_out_data_400; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_401 = mau_4_io_pipe_phv_out_data_401; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_402 = mau_4_io_pipe_phv_out_data_402; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_403 = mau_4_io_pipe_phv_out_data_403; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_404 = mau_4_io_pipe_phv_out_data_404; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_405 = mau_4_io_pipe_phv_out_data_405; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_406 = mau_4_io_pipe_phv_out_data_406; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_407 = mau_4_io_pipe_phv_out_data_407; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_408 = mau_4_io_pipe_phv_out_data_408; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_409 = mau_4_io_pipe_phv_out_data_409; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_410 = mau_4_io_pipe_phv_out_data_410; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_411 = mau_4_io_pipe_phv_out_data_411; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_412 = mau_4_io_pipe_phv_out_data_412; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_413 = mau_4_io_pipe_phv_out_data_413; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_414 = mau_4_io_pipe_phv_out_data_414; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_415 = mau_4_io_pipe_phv_out_data_415; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_416 = mau_4_io_pipe_phv_out_data_416; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_417 = mau_4_io_pipe_phv_out_data_417; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_418 = mau_4_io_pipe_phv_out_data_418; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_419 = mau_4_io_pipe_phv_out_data_419; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_420 = mau_4_io_pipe_phv_out_data_420; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_421 = mau_4_io_pipe_phv_out_data_421; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_422 = mau_4_io_pipe_phv_out_data_422; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_423 = mau_4_io_pipe_phv_out_data_423; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_424 = mau_4_io_pipe_phv_out_data_424; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_425 = mau_4_io_pipe_phv_out_data_425; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_426 = mau_4_io_pipe_phv_out_data_426; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_427 = mau_4_io_pipe_phv_out_data_427; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_428 = mau_4_io_pipe_phv_out_data_428; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_429 = mau_4_io_pipe_phv_out_data_429; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_430 = mau_4_io_pipe_phv_out_data_430; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_431 = mau_4_io_pipe_phv_out_data_431; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_432 = mau_4_io_pipe_phv_out_data_432; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_433 = mau_4_io_pipe_phv_out_data_433; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_434 = mau_4_io_pipe_phv_out_data_434; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_435 = mau_4_io_pipe_phv_out_data_435; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_436 = mau_4_io_pipe_phv_out_data_436; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_437 = mau_4_io_pipe_phv_out_data_437; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_438 = mau_4_io_pipe_phv_out_data_438; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_439 = mau_4_io_pipe_phv_out_data_439; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_440 = mau_4_io_pipe_phv_out_data_440; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_441 = mau_4_io_pipe_phv_out_data_441; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_442 = mau_4_io_pipe_phv_out_data_442; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_443 = mau_4_io_pipe_phv_out_data_443; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_444 = mau_4_io_pipe_phv_out_data_444; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_445 = mau_4_io_pipe_phv_out_data_445; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_446 = mau_4_io_pipe_phv_out_data_446; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_447 = mau_4_io_pipe_phv_out_data_447; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_448 = mau_4_io_pipe_phv_out_data_448; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_449 = mau_4_io_pipe_phv_out_data_449; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_450 = mau_4_io_pipe_phv_out_data_450; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_451 = mau_4_io_pipe_phv_out_data_451; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_452 = mau_4_io_pipe_phv_out_data_452; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_453 = mau_4_io_pipe_phv_out_data_453; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_454 = mau_4_io_pipe_phv_out_data_454; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_455 = mau_4_io_pipe_phv_out_data_455; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_456 = mau_4_io_pipe_phv_out_data_456; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_457 = mau_4_io_pipe_phv_out_data_457; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_458 = mau_4_io_pipe_phv_out_data_458; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_459 = mau_4_io_pipe_phv_out_data_459; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_460 = mau_4_io_pipe_phv_out_data_460; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_461 = mau_4_io_pipe_phv_out_data_461; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_462 = mau_4_io_pipe_phv_out_data_462; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_463 = mau_4_io_pipe_phv_out_data_463; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_464 = mau_4_io_pipe_phv_out_data_464; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_465 = mau_4_io_pipe_phv_out_data_465; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_466 = mau_4_io_pipe_phv_out_data_466; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_467 = mau_4_io_pipe_phv_out_data_467; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_468 = mau_4_io_pipe_phv_out_data_468; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_469 = mau_4_io_pipe_phv_out_data_469; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_470 = mau_4_io_pipe_phv_out_data_470; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_471 = mau_4_io_pipe_phv_out_data_471; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_472 = mau_4_io_pipe_phv_out_data_472; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_473 = mau_4_io_pipe_phv_out_data_473; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_474 = mau_4_io_pipe_phv_out_data_474; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_475 = mau_4_io_pipe_phv_out_data_475; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_476 = mau_4_io_pipe_phv_out_data_476; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_477 = mau_4_io_pipe_phv_out_data_477; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_478 = mau_4_io_pipe_phv_out_data_478; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_479 = mau_4_io_pipe_phv_out_data_479; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_480 = mau_4_io_pipe_phv_out_data_480; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_481 = mau_4_io_pipe_phv_out_data_481; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_482 = mau_4_io_pipe_phv_out_data_482; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_483 = mau_4_io_pipe_phv_out_data_483; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_484 = mau_4_io_pipe_phv_out_data_484; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_485 = mau_4_io_pipe_phv_out_data_485; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_486 = mau_4_io_pipe_phv_out_data_486; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_487 = mau_4_io_pipe_phv_out_data_487; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_488 = mau_4_io_pipe_phv_out_data_488; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_489 = mau_4_io_pipe_phv_out_data_489; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_490 = mau_4_io_pipe_phv_out_data_490; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_491 = mau_4_io_pipe_phv_out_data_491; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_492 = mau_4_io_pipe_phv_out_data_492; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_493 = mau_4_io_pipe_phv_out_data_493; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_494 = mau_4_io_pipe_phv_out_data_494; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_495 = mau_4_io_pipe_phv_out_data_495; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_496 = mau_4_io_pipe_phv_out_data_496; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_497 = mau_4_io_pipe_phv_out_data_497; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_498 = mau_4_io_pipe_phv_out_data_498; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_499 = mau_4_io_pipe_phv_out_data_499; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_500 = mau_4_io_pipe_phv_out_data_500; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_501 = mau_4_io_pipe_phv_out_data_501; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_502 = mau_4_io_pipe_phv_out_data_502; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_503 = mau_4_io_pipe_phv_out_data_503; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_504 = mau_4_io_pipe_phv_out_data_504; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_505 = mau_4_io_pipe_phv_out_data_505; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_506 = mau_4_io_pipe_phv_out_data_506; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_507 = mau_4_io_pipe_phv_out_data_507; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_508 = mau_4_io_pipe_phv_out_data_508; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_509 = mau_4_io_pipe_phv_out_data_509; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_510 = mau_4_io_pipe_phv_out_data_510; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_511 = mau_4_io_pipe_phv_out_data_511; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_header_0 = mau_4_io_pipe_phv_out_header_0; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_header_1 = mau_4_io_pipe_phv_out_header_1; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_header_2 = mau_4_io_pipe_phv_out_header_2; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_header_3 = mau_4_io_pipe_phv_out_header_3; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_header_4 = mau_4_io_pipe_phv_out_header_4; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_header_5 = mau_4_io_pipe_phv_out_header_5; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_header_6 = mau_4_io_pipe_phv_out_header_6; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_header_7 = mau_4_io_pipe_phv_out_header_7; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_header_8 = mau_4_io_pipe_phv_out_header_8; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_header_9 = mau_4_io_pipe_phv_out_header_9; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_header_10 = mau_4_io_pipe_phv_out_header_10; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_header_11 = mau_4_io_pipe_phv_out_header_11; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_header_12 = mau_4_io_pipe_phv_out_header_12; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_header_13 = mau_4_io_pipe_phv_out_header_13; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_header_14 = mau_4_io_pipe_phv_out_header_14; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_header_15 = mau_4_io_pipe_phv_out_header_15; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_parse_current_state = mau_4_io_pipe_phv_out_parse_current_state; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_parse_current_offset = mau_4_io_pipe_phv_out_parse_current_offset; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_parse_transition_field = mau_4_io_pipe_phv_out_parse_transition_field; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_next_processor_id = mau_4_io_pipe_phv_out_next_processor_id; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_next_config_id = mau_4_io_pipe_phv_out_next_config_id; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_is_valid_processor = mau_4_io_pipe_phv_out_is_valid_processor; // @[parser_pisa.scala 42:35]
  assign mau_5_io_mod_state_id_mod = io_mod_en ? io_mod_module_mod_state_id_mod & mod_j_5 :
    io_mod_module_mod_state_id_mod; // @[parser_pisa.scala 51:22 parser_pisa.scala 58:40 parser_pisa.scala 47:23]
  assign mau_5_io_mod_state_id = io_mod_module_mod_state_id; // @[parser_pisa.scala 47:23]
  assign mau_5_io_mod_sram_w_cs = io_mod_module_mod_sram_w_cs; // @[parser_pisa.scala 47:23]
  assign mau_5_io_mod_sram_w_en = io_mod_en ? io_mod_module_mod_sram_w_en & mod_j_5 : io_mod_module_mod_sram_w_en; // @[parser_pisa.scala 51:22 parser_pisa.scala 57:40 parser_pisa.scala 47:23]
  assign mau_5_io_mod_sram_w_addr = io_mod_module_mod_sram_w_addr; // @[parser_pisa.scala 47:23]
  assign mau_5_io_mod_sram_w_data = io_mod_module_mod_sram_w_data; // @[parser_pisa.scala 47:23]
  assign mau_6_clock = clock;
  assign mau_6_io_pipe_phv_in_data_0 = mau_5_io_pipe_phv_out_data_0; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_1 = mau_5_io_pipe_phv_out_data_1; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_2 = mau_5_io_pipe_phv_out_data_2; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_3 = mau_5_io_pipe_phv_out_data_3; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_4 = mau_5_io_pipe_phv_out_data_4; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_5 = mau_5_io_pipe_phv_out_data_5; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_6 = mau_5_io_pipe_phv_out_data_6; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_7 = mau_5_io_pipe_phv_out_data_7; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_8 = mau_5_io_pipe_phv_out_data_8; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_9 = mau_5_io_pipe_phv_out_data_9; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_10 = mau_5_io_pipe_phv_out_data_10; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_11 = mau_5_io_pipe_phv_out_data_11; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_12 = mau_5_io_pipe_phv_out_data_12; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_13 = mau_5_io_pipe_phv_out_data_13; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_14 = mau_5_io_pipe_phv_out_data_14; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_15 = mau_5_io_pipe_phv_out_data_15; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_16 = mau_5_io_pipe_phv_out_data_16; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_17 = mau_5_io_pipe_phv_out_data_17; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_18 = mau_5_io_pipe_phv_out_data_18; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_19 = mau_5_io_pipe_phv_out_data_19; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_20 = mau_5_io_pipe_phv_out_data_20; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_21 = mau_5_io_pipe_phv_out_data_21; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_22 = mau_5_io_pipe_phv_out_data_22; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_23 = mau_5_io_pipe_phv_out_data_23; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_24 = mau_5_io_pipe_phv_out_data_24; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_25 = mau_5_io_pipe_phv_out_data_25; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_26 = mau_5_io_pipe_phv_out_data_26; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_27 = mau_5_io_pipe_phv_out_data_27; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_28 = mau_5_io_pipe_phv_out_data_28; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_29 = mau_5_io_pipe_phv_out_data_29; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_30 = mau_5_io_pipe_phv_out_data_30; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_31 = mau_5_io_pipe_phv_out_data_31; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_32 = mau_5_io_pipe_phv_out_data_32; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_33 = mau_5_io_pipe_phv_out_data_33; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_34 = mau_5_io_pipe_phv_out_data_34; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_35 = mau_5_io_pipe_phv_out_data_35; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_36 = mau_5_io_pipe_phv_out_data_36; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_37 = mau_5_io_pipe_phv_out_data_37; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_38 = mau_5_io_pipe_phv_out_data_38; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_39 = mau_5_io_pipe_phv_out_data_39; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_40 = mau_5_io_pipe_phv_out_data_40; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_41 = mau_5_io_pipe_phv_out_data_41; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_42 = mau_5_io_pipe_phv_out_data_42; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_43 = mau_5_io_pipe_phv_out_data_43; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_44 = mau_5_io_pipe_phv_out_data_44; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_45 = mau_5_io_pipe_phv_out_data_45; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_46 = mau_5_io_pipe_phv_out_data_46; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_47 = mau_5_io_pipe_phv_out_data_47; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_48 = mau_5_io_pipe_phv_out_data_48; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_49 = mau_5_io_pipe_phv_out_data_49; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_50 = mau_5_io_pipe_phv_out_data_50; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_51 = mau_5_io_pipe_phv_out_data_51; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_52 = mau_5_io_pipe_phv_out_data_52; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_53 = mau_5_io_pipe_phv_out_data_53; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_54 = mau_5_io_pipe_phv_out_data_54; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_55 = mau_5_io_pipe_phv_out_data_55; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_56 = mau_5_io_pipe_phv_out_data_56; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_57 = mau_5_io_pipe_phv_out_data_57; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_58 = mau_5_io_pipe_phv_out_data_58; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_59 = mau_5_io_pipe_phv_out_data_59; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_60 = mau_5_io_pipe_phv_out_data_60; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_61 = mau_5_io_pipe_phv_out_data_61; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_62 = mau_5_io_pipe_phv_out_data_62; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_63 = mau_5_io_pipe_phv_out_data_63; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_64 = mau_5_io_pipe_phv_out_data_64; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_65 = mau_5_io_pipe_phv_out_data_65; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_66 = mau_5_io_pipe_phv_out_data_66; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_67 = mau_5_io_pipe_phv_out_data_67; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_68 = mau_5_io_pipe_phv_out_data_68; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_69 = mau_5_io_pipe_phv_out_data_69; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_70 = mau_5_io_pipe_phv_out_data_70; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_71 = mau_5_io_pipe_phv_out_data_71; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_72 = mau_5_io_pipe_phv_out_data_72; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_73 = mau_5_io_pipe_phv_out_data_73; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_74 = mau_5_io_pipe_phv_out_data_74; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_75 = mau_5_io_pipe_phv_out_data_75; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_76 = mau_5_io_pipe_phv_out_data_76; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_77 = mau_5_io_pipe_phv_out_data_77; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_78 = mau_5_io_pipe_phv_out_data_78; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_79 = mau_5_io_pipe_phv_out_data_79; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_80 = mau_5_io_pipe_phv_out_data_80; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_81 = mau_5_io_pipe_phv_out_data_81; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_82 = mau_5_io_pipe_phv_out_data_82; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_83 = mau_5_io_pipe_phv_out_data_83; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_84 = mau_5_io_pipe_phv_out_data_84; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_85 = mau_5_io_pipe_phv_out_data_85; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_86 = mau_5_io_pipe_phv_out_data_86; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_87 = mau_5_io_pipe_phv_out_data_87; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_88 = mau_5_io_pipe_phv_out_data_88; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_89 = mau_5_io_pipe_phv_out_data_89; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_90 = mau_5_io_pipe_phv_out_data_90; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_91 = mau_5_io_pipe_phv_out_data_91; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_92 = mau_5_io_pipe_phv_out_data_92; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_93 = mau_5_io_pipe_phv_out_data_93; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_94 = mau_5_io_pipe_phv_out_data_94; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_95 = mau_5_io_pipe_phv_out_data_95; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_96 = mau_5_io_pipe_phv_out_data_96; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_97 = mau_5_io_pipe_phv_out_data_97; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_98 = mau_5_io_pipe_phv_out_data_98; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_99 = mau_5_io_pipe_phv_out_data_99; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_100 = mau_5_io_pipe_phv_out_data_100; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_101 = mau_5_io_pipe_phv_out_data_101; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_102 = mau_5_io_pipe_phv_out_data_102; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_103 = mau_5_io_pipe_phv_out_data_103; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_104 = mau_5_io_pipe_phv_out_data_104; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_105 = mau_5_io_pipe_phv_out_data_105; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_106 = mau_5_io_pipe_phv_out_data_106; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_107 = mau_5_io_pipe_phv_out_data_107; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_108 = mau_5_io_pipe_phv_out_data_108; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_109 = mau_5_io_pipe_phv_out_data_109; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_110 = mau_5_io_pipe_phv_out_data_110; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_111 = mau_5_io_pipe_phv_out_data_111; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_112 = mau_5_io_pipe_phv_out_data_112; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_113 = mau_5_io_pipe_phv_out_data_113; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_114 = mau_5_io_pipe_phv_out_data_114; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_115 = mau_5_io_pipe_phv_out_data_115; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_116 = mau_5_io_pipe_phv_out_data_116; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_117 = mau_5_io_pipe_phv_out_data_117; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_118 = mau_5_io_pipe_phv_out_data_118; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_119 = mau_5_io_pipe_phv_out_data_119; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_120 = mau_5_io_pipe_phv_out_data_120; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_121 = mau_5_io_pipe_phv_out_data_121; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_122 = mau_5_io_pipe_phv_out_data_122; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_123 = mau_5_io_pipe_phv_out_data_123; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_124 = mau_5_io_pipe_phv_out_data_124; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_125 = mau_5_io_pipe_phv_out_data_125; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_126 = mau_5_io_pipe_phv_out_data_126; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_127 = mau_5_io_pipe_phv_out_data_127; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_128 = mau_5_io_pipe_phv_out_data_128; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_129 = mau_5_io_pipe_phv_out_data_129; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_130 = mau_5_io_pipe_phv_out_data_130; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_131 = mau_5_io_pipe_phv_out_data_131; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_132 = mau_5_io_pipe_phv_out_data_132; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_133 = mau_5_io_pipe_phv_out_data_133; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_134 = mau_5_io_pipe_phv_out_data_134; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_135 = mau_5_io_pipe_phv_out_data_135; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_136 = mau_5_io_pipe_phv_out_data_136; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_137 = mau_5_io_pipe_phv_out_data_137; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_138 = mau_5_io_pipe_phv_out_data_138; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_139 = mau_5_io_pipe_phv_out_data_139; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_140 = mau_5_io_pipe_phv_out_data_140; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_141 = mau_5_io_pipe_phv_out_data_141; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_142 = mau_5_io_pipe_phv_out_data_142; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_143 = mau_5_io_pipe_phv_out_data_143; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_144 = mau_5_io_pipe_phv_out_data_144; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_145 = mau_5_io_pipe_phv_out_data_145; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_146 = mau_5_io_pipe_phv_out_data_146; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_147 = mau_5_io_pipe_phv_out_data_147; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_148 = mau_5_io_pipe_phv_out_data_148; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_149 = mau_5_io_pipe_phv_out_data_149; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_150 = mau_5_io_pipe_phv_out_data_150; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_151 = mau_5_io_pipe_phv_out_data_151; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_152 = mau_5_io_pipe_phv_out_data_152; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_153 = mau_5_io_pipe_phv_out_data_153; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_154 = mau_5_io_pipe_phv_out_data_154; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_155 = mau_5_io_pipe_phv_out_data_155; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_156 = mau_5_io_pipe_phv_out_data_156; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_157 = mau_5_io_pipe_phv_out_data_157; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_158 = mau_5_io_pipe_phv_out_data_158; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_159 = mau_5_io_pipe_phv_out_data_159; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_160 = mau_5_io_pipe_phv_out_data_160; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_161 = mau_5_io_pipe_phv_out_data_161; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_162 = mau_5_io_pipe_phv_out_data_162; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_163 = mau_5_io_pipe_phv_out_data_163; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_164 = mau_5_io_pipe_phv_out_data_164; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_165 = mau_5_io_pipe_phv_out_data_165; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_166 = mau_5_io_pipe_phv_out_data_166; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_167 = mau_5_io_pipe_phv_out_data_167; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_168 = mau_5_io_pipe_phv_out_data_168; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_169 = mau_5_io_pipe_phv_out_data_169; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_170 = mau_5_io_pipe_phv_out_data_170; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_171 = mau_5_io_pipe_phv_out_data_171; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_172 = mau_5_io_pipe_phv_out_data_172; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_173 = mau_5_io_pipe_phv_out_data_173; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_174 = mau_5_io_pipe_phv_out_data_174; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_175 = mau_5_io_pipe_phv_out_data_175; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_176 = mau_5_io_pipe_phv_out_data_176; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_177 = mau_5_io_pipe_phv_out_data_177; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_178 = mau_5_io_pipe_phv_out_data_178; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_179 = mau_5_io_pipe_phv_out_data_179; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_180 = mau_5_io_pipe_phv_out_data_180; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_181 = mau_5_io_pipe_phv_out_data_181; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_182 = mau_5_io_pipe_phv_out_data_182; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_183 = mau_5_io_pipe_phv_out_data_183; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_184 = mau_5_io_pipe_phv_out_data_184; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_185 = mau_5_io_pipe_phv_out_data_185; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_186 = mau_5_io_pipe_phv_out_data_186; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_187 = mau_5_io_pipe_phv_out_data_187; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_188 = mau_5_io_pipe_phv_out_data_188; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_189 = mau_5_io_pipe_phv_out_data_189; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_190 = mau_5_io_pipe_phv_out_data_190; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_191 = mau_5_io_pipe_phv_out_data_191; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_192 = mau_5_io_pipe_phv_out_data_192; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_193 = mau_5_io_pipe_phv_out_data_193; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_194 = mau_5_io_pipe_phv_out_data_194; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_195 = mau_5_io_pipe_phv_out_data_195; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_196 = mau_5_io_pipe_phv_out_data_196; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_197 = mau_5_io_pipe_phv_out_data_197; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_198 = mau_5_io_pipe_phv_out_data_198; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_199 = mau_5_io_pipe_phv_out_data_199; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_200 = mau_5_io_pipe_phv_out_data_200; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_201 = mau_5_io_pipe_phv_out_data_201; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_202 = mau_5_io_pipe_phv_out_data_202; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_203 = mau_5_io_pipe_phv_out_data_203; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_204 = mau_5_io_pipe_phv_out_data_204; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_205 = mau_5_io_pipe_phv_out_data_205; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_206 = mau_5_io_pipe_phv_out_data_206; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_207 = mau_5_io_pipe_phv_out_data_207; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_208 = mau_5_io_pipe_phv_out_data_208; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_209 = mau_5_io_pipe_phv_out_data_209; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_210 = mau_5_io_pipe_phv_out_data_210; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_211 = mau_5_io_pipe_phv_out_data_211; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_212 = mau_5_io_pipe_phv_out_data_212; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_213 = mau_5_io_pipe_phv_out_data_213; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_214 = mau_5_io_pipe_phv_out_data_214; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_215 = mau_5_io_pipe_phv_out_data_215; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_216 = mau_5_io_pipe_phv_out_data_216; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_217 = mau_5_io_pipe_phv_out_data_217; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_218 = mau_5_io_pipe_phv_out_data_218; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_219 = mau_5_io_pipe_phv_out_data_219; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_220 = mau_5_io_pipe_phv_out_data_220; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_221 = mau_5_io_pipe_phv_out_data_221; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_222 = mau_5_io_pipe_phv_out_data_222; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_223 = mau_5_io_pipe_phv_out_data_223; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_224 = mau_5_io_pipe_phv_out_data_224; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_225 = mau_5_io_pipe_phv_out_data_225; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_226 = mau_5_io_pipe_phv_out_data_226; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_227 = mau_5_io_pipe_phv_out_data_227; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_228 = mau_5_io_pipe_phv_out_data_228; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_229 = mau_5_io_pipe_phv_out_data_229; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_230 = mau_5_io_pipe_phv_out_data_230; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_231 = mau_5_io_pipe_phv_out_data_231; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_232 = mau_5_io_pipe_phv_out_data_232; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_233 = mau_5_io_pipe_phv_out_data_233; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_234 = mau_5_io_pipe_phv_out_data_234; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_235 = mau_5_io_pipe_phv_out_data_235; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_236 = mau_5_io_pipe_phv_out_data_236; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_237 = mau_5_io_pipe_phv_out_data_237; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_238 = mau_5_io_pipe_phv_out_data_238; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_239 = mau_5_io_pipe_phv_out_data_239; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_240 = mau_5_io_pipe_phv_out_data_240; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_241 = mau_5_io_pipe_phv_out_data_241; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_242 = mau_5_io_pipe_phv_out_data_242; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_243 = mau_5_io_pipe_phv_out_data_243; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_244 = mau_5_io_pipe_phv_out_data_244; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_245 = mau_5_io_pipe_phv_out_data_245; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_246 = mau_5_io_pipe_phv_out_data_246; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_247 = mau_5_io_pipe_phv_out_data_247; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_248 = mau_5_io_pipe_phv_out_data_248; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_249 = mau_5_io_pipe_phv_out_data_249; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_250 = mau_5_io_pipe_phv_out_data_250; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_251 = mau_5_io_pipe_phv_out_data_251; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_252 = mau_5_io_pipe_phv_out_data_252; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_253 = mau_5_io_pipe_phv_out_data_253; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_254 = mau_5_io_pipe_phv_out_data_254; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_255 = mau_5_io_pipe_phv_out_data_255; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_256 = mau_5_io_pipe_phv_out_data_256; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_257 = mau_5_io_pipe_phv_out_data_257; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_258 = mau_5_io_pipe_phv_out_data_258; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_259 = mau_5_io_pipe_phv_out_data_259; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_260 = mau_5_io_pipe_phv_out_data_260; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_261 = mau_5_io_pipe_phv_out_data_261; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_262 = mau_5_io_pipe_phv_out_data_262; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_263 = mau_5_io_pipe_phv_out_data_263; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_264 = mau_5_io_pipe_phv_out_data_264; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_265 = mau_5_io_pipe_phv_out_data_265; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_266 = mau_5_io_pipe_phv_out_data_266; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_267 = mau_5_io_pipe_phv_out_data_267; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_268 = mau_5_io_pipe_phv_out_data_268; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_269 = mau_5_io_pipe_phv_out_data_269; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_270 = mau_5_io_pipe_phv_out_data_270; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_271 = mau_5_io_pipe_phv_out_data_271; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_272 = mau_5_io_pipe_phv_out_data_272; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_273 = mau_5_io_pipe_phv_out_data_273; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_274 = mau_5_io_pipe_phv_out_data_274; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_275 = mau_5_io_pipe_phv_out_data_275; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_276 = mau_5_io_pipe_phv_out_data_276; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_277 = mau_5_io_pipe_phv_out_data_277; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_278 = mau_5_io_pipe_phv_out_data_278; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_279 = mau_5_io_pipe_phv_out_data_279; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_280 = mau_5_io_pipe_phv_out_data_280; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_281 = mau_5_io_pipe_phv_out_data_281; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_282 = mau_5_io_pipe_phv_out_data_282; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_283 = mau_5_io_pipe_phv_out_data_283; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_284 = mau_5_io_pipe_phv_out_data_284; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_285 = mau_5_io_pipe_phv_out_data_285; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_286 = mau_5_io_pipe_phv_out_data_286; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_287 = mau_5_io_pipe_phv_out_data_287; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_288 = mau_5_io_pipe_phv_out_data_288; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_289 = mau_5_io_pipe_phv_out_data_289; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_290 = mau_5_io_pipe_phv_out_data_290; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_291 = mau_5_io_pipe_phv_out_data_291; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_292 = mau_5_io_pipe_phv_out_data_292; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_293 = mau_5_io_pipe_phv_out_data_293; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_294 = mau_5_io_pipe_phv_out_data_294; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_295 = mau_5_io_pipe_phv_out_data_295; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_296 = mau_5_io_pipe_phv_out_data_296; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_297 = mau_5_io_pipe_phv_out_data_297; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_298 = mau_5_io_pipe_phv_out_data_298; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_299 = mau_5_io_pipe_phv_out_data_299; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_300 = mau_5_io_pipe_phv_out_data_300; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_301 = mau_5_io_pipe_phv_out_data_301; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_302 = mau_5_io_pipe_phv_out_data_302; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_303 = mau_5_io_pipe_phv_out_data_303; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_304 = mau_5_io_pipe_phv_out_data_304; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_305 = mau_5_io_pipe_phv_out_data_305; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_306 = mau_5_io_pipe_phv_out_data_306; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_307 = mau_5_io_pipe_phv_out_data_307; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_308 = mau_5_io_pipe_phv_out_data_308; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_309 = mau_5_io_pipe_phv_out_data_309; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_310 = mau_5_io_pipe_phv_out_data_310; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_311 = mau_5_io_pipe_phv_out_data_311; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_312 = mau_5_io_pipe_phv_out_data_312; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_313 = mau_5_io_pipe_phv_out_data_313; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_314 = mau_5_io_pipe_phv_out_data_314; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_315 = mau_5_io_pipe_phv_out_data_315; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_316 = mau_5_io_pipe_phv_out_data_316; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_317 = mau_5_io_pipe_phv_out_data_317; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_318 = mau_5_io_pipe_phv_out_data_318; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_319 = mau_5_io_pipe_phv_out_data_319; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_320 = mau_5_io_pipe_phv_out_data_320; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_321 = mau_5_io_pipe_phv_out_data_321; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_322 = mau_5_io_pipe_phv_out_data_322; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_323 = mau_5_io_pipe_phv_out_data_323; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_324 = mau_5_io_pipe_phv_out_data_324; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_325 = mau_5_io_pipe_phv_out_data_325; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_326 = mau_5_io_pipe_phv_out_data_326; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_327 = mau_5_io_pipe_phv_out_data_327; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_328 = mau_5_io_pipe_phv_out_data_328; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_329 = mau_5_io_pipe_phv_out_data_329; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_330 = mau_5_io_pipe_phv_out_data_330; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_331 = mau_5_io_pipe_phv_out_data_331; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_332 = mau_5_io_pipe_phv_out_data_332; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_333 = mau_5_io_pipe_phv_out_data_333; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_334 = mau_5_io_pipe_phv_out_data_334; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_335 = mau_5_io_pipe_phv_out_data_335; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_336 = mau_5_io_pipe_phv_out_data_336; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_337 = mau_5_io_pipe_phv_out_data_337; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_338 = mau_5_io_pipe_phv_out_data_338; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_339 = mau_5_io_pipe_phv_out_data_339; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_340 = mau_5_io_pipe_phv_out_data_340; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_341 = mau_5_io_pipe_phv_out_data_341; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_342 = mau_5_io_pipe_phv_out_data_342; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_343 = mau_5_io_pipe_phv_out_data_343; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_344 = mau_5_io_pipe_phv_out_data_344; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_345 = mau_5_io_pipe_phv_out_data_345; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_346 = mau_5_io_pipe_phv_out_data_346; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_347 = mau_5_io_pipe_phv_out_data_347; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_348 = mau_5_io_pipe_phv_out_data_348; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_349 = mau_5_io_pipe_phv_out_data_349; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_350 = mau_5_io_pipe_phv_out_data_350; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_351 = mau_5_io_pipe_phv_out_data_351; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_352 = mau_5_io_pipe_phv_out_data_352; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_353 = mau_5_io_pipe_phv_out_data_353; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_354 = mau_5_io_pipe_phv_out_data_354; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_355 = mau_5_io_pipe_phv_out_data_355; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_356 = mau_5_io_pipe_phv_out_data_356; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_357 = mau_5_io_pipe_phv_out_data_357; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_358 = mau_5_io_pipe_phv_out_data_358; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_359 = mau_5_io_pipe_phv_out_data_359; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_360 = mau_5_io_pipe_phv_out_data_360; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_361 = mau_5_io_pipe_phv_out_data_361; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_362 = mau_5_io_pipe_phv_out_data_362; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_363 = mau_5_io_pipe_phv_out_data_363; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_364 = mau_5_io_pipe_phv_out_data_364; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_365 = mau_5_io_pipe_phv_out_data_365; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_366 = mau_5_io_pipe_phv_out_data_366; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_367 = mau_5_io_pipe_phv_out_data_367; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_368 = mau_5_io_pipe_phv_out_data_368; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_369 = mau_5_io_pipe_phv_out_data_369; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_370 = mau_5_io_pipe_phv_out_data_370; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_371 = mau_5_io_pipe_phv_out_data_371; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_372 = mau_5_io_pipe_phv_out_data_372; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_373 = mau_5_io_pipe_phv_out_data_373; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_374 = mau_5_io_pipe_phv_out_data_374; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_375 = mau_5_io_pipe_phv_out_data_375; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_376 = mau_5_io_pipe_phv_out_data_376; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_377 = mau_5_io_pipe_phv_out_data_377; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_378 = mau_5_io_pipe_phv_out_data_378; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_379 = mau_5_io_pipe_phv_out_data_379; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_380 = mau_5_io_pipe_phv_out_data_380; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_381 = mau_5_io_pipe_phv_out_data_381; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_382 = mau_5_io_pipe_phv_out_data_382; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_383 = mau_5_io_pipe_phv_out_data_383; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_384 = mau_5_io_pipe_phv_out_data_384; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_385 = mau_5_io_pipe_phv_out_data_385; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_386 = mau_5_io_pipe_phv_out_data_386; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_387 = mau_5_io_pipe_phv_out_data_387; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_388 = mau_5_io_pipe_phv_out_data_388; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_389 = mau_5_io_pipe_phv_out_data_389; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_390 = mau_5_io_pipe_phv_out_data_390; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_391 = mau_5_io_pipe_phv_out_data_391; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_392 = mau_5_io_pipe_phv_out_data_392; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_393 = mau_5_io_pipe_phv_out_data_393; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_394 = mau_5_io_pipe_phv_out_data_394; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_395 = mau_5_io_pipe_phv_out_data_395; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_396 = mau_5_io_pipe_phv_out_data_396; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_397 = mau_5_io_pipe_phv_out_data_397; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_398 = mau_5_io_pipe_phv_out_data_398; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_399 = mau_5_io_pipe_phv_out_data_399; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_400 = mau_5_io_pipe_phv_out_data_400; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_401 = mau_5_io_pipe_phv_out_data_401; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_402 = mau_5_io_pipe_phv_out_data_402; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_403 = mau_5_io_pipe_phv_out_data_403; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_404 = mau_5_io_pipe_phv_out_data_404; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_405 = mau_5_io_pipe_phv_out_data_405; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_406 = mau_5_io_pipe_phv_out_data_406; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_407 = mau_5_io_pipe_phv_out_data_407; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_408 = mau_5_io_pipe_phv_out_data_408; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_409 = mau_5_io_pipe_phv_out_data_409; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_410 = mau_5_io_pipe_phv_out_data_410; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_411 = mau_5_io_pipe_phv_out_data_411; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_412 = mau_5_io_pipe_phv_out_data_412; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_413 = mau_5_io_pipe_phv_out_data_413; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_414 = mau_5_io_pipe_phv_out_data_414; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_415 = mau_5_io_pipe_phv_out_data_415; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_416 = mau_5_io_pipe_phv_out_data_416; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_417 = mau_5_io_pipe_phv_out_data_417; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_418 = mau_5_io_pipe_phv_out_data_418; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_419 = mau_5_io_pipe_phv_out_data_419; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_420 = mau_5_io_pipe_phv_out_data_420; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_421 = mau_5_io_pipe_phv_out_data_421; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_422 = mau_5_io_pipe_phv_out_data_422; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_423 = mau_5_io_pipe_phv_out_data_423; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_424 = mau_5_io_pipe_phv_out_data_424; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_425 = mau_5_io_pipe_phv_out_data_425; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_426 = mau_5_io_pipe_phv_out_data_426; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_427 = mau_5_io_pipe_phv_out_data_427; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_428 = mau_5_io_pipe_phv_out_data_428; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_429 = mau_5_io_pipe_phv_out_data_429; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_430 = mau_5_io_pipe_phv_out_data_430; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_431 = mau_5_io_pipe_phv_out_data_431; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_432 = mau_5_io_pipe_phv_out_data_432; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_433 = mau_5_io_pipe_phv_out_data_433; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_434 = mau_5_io_pipe_phv_out_data_434; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_435 = mau_5_io_pipe_phv_out_data_435; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_436 = mau_5_io_pipe_phv_out_data_436; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_437 = mau_5_io_pipe_phv_out_data_437; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_438 = mau_5_io_pipe_phv_out_data_438; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_439 = mau_5_io_pipe_phv_out_data_439; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_440 = mau_5_io_pipe_phv_out_data_440; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_441 = mau_5_io_pipe_phv_out_data_441; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_442 = mau_5_io_pipe_phv_out_data_442; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_443 = mau_5_io_pipe_phv_out_data_443; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_444 = mau_5_io_pipe_phv_out_data_444; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_445 = mau_5_io_pipe_phv_out_data_445; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_446 = mau_5_io_pipe_phv_out_data_446; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_447 = mau_5_io_pipe_phv_out_data_447; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_448 = mau_5_io_pipe_phv_out_data_448; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_449 = mau_5_io_pipe_phv_out_data_449; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_450 = mau_5_io_pipe_phv_out_data_450; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_451 = mau_5_io_pipe_phv_out_data_451; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_452 = mau_5_io_pipe_phv_out_data_452; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_453 = mau_5_io_pipe_phv_out_data_453; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_454 = mau_5_io_pipe_phv_out_data_454; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_455 = mau_5_io_pipe_phv_out_data_455; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_456 = mau_5_io_pipe_phv_out_data_456; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_457 = mau_5_io_pipe_phv_out_data_457; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_458 = mau_5_io_pipe_phv_out_data_458; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_459 = mau_5_io_pipe_phv_out_data_459; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_460 = mau_5_io_pipe_phv_out_data_460; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_461 = mau_5_io_pipe_phv_out_data_461; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_462 = mau_5_io_pipe_phv_out_data_462; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_463 = mau_5_io_pipe_phv_out_data_463; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_464 = mau_5_io_pipe_phv_out_data_464; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_465 = mau_5_io_pipe_phv_out_data_465; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_466 = mau_5_io_pipe_phv_out_data_466; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_467 = mau_5_io_pipe_phv_out_data_467; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_468 = mau_5_io_pipe_phv_out_data_468; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_469 = mau_5_io_pipe_phv_out_data_469; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_470 = mau_5_io_pipe_phv_out_data_470; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_471 = mau_5_io_pipe_phv_out_data_471; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_472 = mau_5_io_pipe_phv_out_data_472; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_473 = mau_5_io_pipe_phv_out_data_473; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_474 = mau_5_io_pipe_phv_out_data_474; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_475 = mau_5_io_pipe_phv_out_data_475; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_476 = mau_5_io_pipe_phv_out_data_476; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_477 = mau_5_io_pipe_phv_out_data_477; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_478 = mau_5_io_pipe_phv_out_data_478; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_479 = mau_5_io_pipe_phv_out_data_479; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_480 = mau_5_io_pipe_phv_out_data_480; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_481 = mau_5_io_pipe_phv_out_data_481; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_482 = mau_5_io_pipe_phv_out_data_482; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_483 = mau_5_io_pipe_phv_out_data_483; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_484 = mau_5_io_pipe_phv_out_data_484; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_485 = mau_5_io_pipe_phv_out_data_485; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_486 = mau_5_io_pipe_phv_out_data_486; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_487 = mau_5_io_pipe_phv_out_data_487; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_488 = mau_5_io_pipe_phv_out_data_488; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_489 = mau_5_io_pipe_phv_out_data_489; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_490 = mau_5_io_pipe_phv_out_data_490; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_491 = mau_5_io_pipe_phv_out_data_491; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_492 = mau_5_io_pipe_phv_out_data_492; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_493 = mau_5_io_pipe_phv_out_data_493; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_494 = mau_5_io_pipe_phv_out_data_494; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_495 = mau_5_io_pipe_phv_out_data_495; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_496 = mau_5_io_pipe_phv_out_data_496; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_497 = mau_5_io_pipe_phv_out_data_497; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_498 = mau_5_io_pipe_phv_out_data_498; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_499 = mau_5_io_pipe_phv_out_data_499; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_500 = mau_5_io_pipe_phv_out_data_500; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_501 = mau_5_io_pipe_phv_out_data_501; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_502 = mau_5_io_pipe_phv_out_data_502; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_503 = mau_5_io_pipe_phv_out_data_503; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_504 = mau_5_io_pipe_phv_out_data_504; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_505 = mau_5_io_pipe_phv_out_data_505; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_506 = mau_5_io_pipe_phv_out_data_506; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_507 = mau_5_io_pipe_phv_out_data_507; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_508 = mau_5_io_pipe_phv_out_data_508; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_509 = mau_5_io_pipe_phv_out_data_509; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_510 = mau_5_io_pipe_phv_out_data_510; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_511 = mau_5_io_pipe_phv_out_data_511; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_header_0 = mau_5_io_pipe_phv_out_header_0; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_header_1 = mau_5_io_pipe_phv_out_header_1; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_header_2 = mau_5_io_pipe_phv_out_header_2; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_header_3 = mau_5_io_pipe_phv_out_header_3; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_header_4 = mau_5_io_pipe_phv_out_header_4; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_header_5 = mau_5_io_pipe_phv_out_header_5; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_header_6 = mau_5_io_pipe_phv_out_header_6; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_header_7 = mau_5_io_pipe_phv_out_header_7; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_header_8 = mau_5_io_pipe_phv_out_header_8; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_header_9 = mau_5_io_pipe_phv_out_header_9; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_header_10 = mau_5_io_pipe_phv_out_header_10; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_header_11 = mau_5_io_pipe_phv_out_header_11; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_header_12 = mau_5_io_pipe_phv_out_header_12; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_header_13 = mau_5_io_pipe_phv_out_header_13; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_header_14 = mau_5_io_pipe_phv_out_header_14; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_header_15 = mau_5_io_pipe_phv_out_header_15; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_parse_current_state = mau_5_io_pipe_phv_out_parse_current_state; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_parse_current_offset = mau_5_io_pipe_phv_out_parse_current_offset; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_parse_transition_field = mau_5_io_pipe_phv_out_parse_transition_field; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_next_processor_id = mau_5_io_pipe_phv_out_next_processor_id; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_next_config_id = mau_5_io_pipe_phv_out_next_config_id; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_is_valid_processor = mau_5_io_pipe_phv_out_is_valid_processor; // @[parser_pisa.scala 42:35]
  assign mau_6_io_mod_state_id_mod = io_mod_en ? io_mod_module_mod_state_id_mod & mod_j_6 :
    io_mod_module_mod_state_id_mod; // @[parser_pisa.scala 51:22 parser_pisa.scala 58:40 parser_pisa.scala 47:23]
  assign mau_6_io_mod_state_id = io_mod_module_mod_state_id; // @[parser_pisa.scala 47:23]
  assign mau_6_io_mod_sram_w_cs = io_mod_module_mod_sram_w_cs; // @[parser_pisa.scala 47:23]
  assign mau_6_io_mod_sram_w_en = io_mod_en ? io_mod_module_mod_sram_w_en & mod_j_6 : io_mod_module_mod_sram_w_en; // @[parser_pisa.scala 51:22 parser_pisa.scala 57:40 parser_pisa.scala 47:23]
  assign mau_6_io_mod_sram_w_addr = io_mod_module_mod_sram_w_addr; // @[parser_pisa.scala 47:23]
  assign mau_6_io_mod_sram_w_data = io_mod_module_mod_sram_w_data; // @[parser_pisa.scala 47:23]
  assign mau_7_clock = clock;
  assign mau_7_io_pipe_phv_in_data_0 = mau_6_io_pipe_phv_out_data_0; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_1 = mau_6_io_pipe_phv_out_data_1; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_2 = mau_6_io_pipe_phv_out_data_2; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_3 = mau_6_io_pipe_phv_out_data_3; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_4 = mau_6_io_pipe_phv_out_data_4; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_5 = mau_6_io_pipe_phv_out_data_5; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_6 = mau_6_io_pipe_phv_out_data_6; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_7 = mau_6_io_pipe_phv_out_data_7; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_8 = mau_6_io_pipe_phv_out_data_8; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_9 = mau_6_io_pipe_phv_out_data_9; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_10 = mau_6_io_pipe_phv_out_data_10; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_11 = mau_6_io_pipe_phv_out_data_11; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_12 = mau_6_io_pipe_phv_out_data_12; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_13 = mau_6_io_pipe_phv_out_data_13; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_14 = mau_6_io_pipe_phv_out_data_14; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_15 = mau_6_io_pipe_phv_out_data_15; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_16 = mau_6_io_pipe_phv_out_data_16; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_17 = mau_6_io_pipe_phv_out_data_17; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_18 = mau_6_io_pipe_phv_out_data_18; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_19 = mau_6_io_pipe_phv_out_data_19; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_20 = mau_6_io_pipe_phv_out_data_20; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_21 = mau_6_io_pipe_phv_out_data_21; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_22 = mau_6_io_pipe_phv_out_data_22; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_23 = mau_6_io_pipe_phv_out_data_23; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_24 = mau_6_io_pipe_phv_out_data_24; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_25 = mau_6_io_pipe_phv_out_data_25; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_26 = mau_6_io_pipe_phv_out_data_26; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_27 = mau_6_io_pipe_phv_out_data_27; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_28 = mau_6_io_pipe_phv_out_data_28; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_29 = mau_6_io_pipe_phv_out_data_29; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_30 = mau_6_io_pipe_phv_out_data_30; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_31 = mau_6_io_pipe_phv_out_data_31; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_32 = mau_6_io_pipe_phv_out_data_32; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_33 = mau_6_io_pipe_phv_out_data_33; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_34 = mau_6_io_pipe_phv_out_data_34; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_35 = mau_6_io_pipe_phv_out_data_35; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_36 = mau_6_io_pipe_phv_out_data_36; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_37 = mau_6_io_pipe_phv_out_data_37; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_38 = mau_6_io_pipe_phv_out_data_38; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_39 = mau_6_io_pipe_phv_out_data_39; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_40 = mau_6_io_pipe_phv_out_data_40; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_41 = mau_6_io_pipe_phv_out_data_41; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_42 = mau_6_io_pipe_phv_out_data_42; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_43 = mau_6_io_pipe_phv_out_data_43; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_44 = mau_6_io_pipe_phv_out_data_44; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_45 = mau_6_io_pipe_phv_out_data_45; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_46 = mau_6_io_pipe_phv_out_data_46; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_47 = mau_6_io_pipe_phv_out_data_47; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_48 = mau_6_io_pipe_phv_out_data_48; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_49 = mau_6_io_pipe_phv_out_data_49; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_50 = mau_6_io_pipe_phv_out_data_50; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_51 = mau_6_io_pipe_phv_out_data_51; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_52 = mau_6_io_pipe_phv_out_data_52; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_53 = mau_6_io_pipe_phv_out_data_53; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_54 = mau_6_io_pipe_phv_out_data_54; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_55 = mau_6_io_pipe_phv_out_data_55; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_56 = mau_6_io_pipe_phv_out_data_56; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_57 = mau_6_io_pipe_phv_out_data_57; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_58 = mau_6_io_pipe_phv_out_data_58; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_59 = mau_6_io_pipe_phv_out_data_59; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_60 = mau_6_io_pipe_phv_out_data_60; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_61 = mau_6_io_pipe_phv_out_data_61; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_62 = mau_6_io_pipe_phv_out_data_62; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_63 = mau_6_io_pipe_phv_out_data_63; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_64 = mau_6_io_pipe_phv_out_data_64; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_65 = mau_6_io_pipe_phv_out_data_65; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_66 = mau_6_io_pipe_phv_out_data_66; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_67 = mau_6_io_pipe_phv_out_data_67; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_68 = mau_6_io_pipe_phv_out_data_68; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_69 = mau_6_io_pipe_phv_out_data_69; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_70 = mau_6_io_pipe_phv_out_data_70; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_71 = mau_6_io_pipe_phv_out_data_71; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_72 = mau_6_io_pipe_phv_out_data_72; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_73 = mau_6_io_pipe_phv_out_data_73; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_74 = mau_6_io_pipe_phv_out_data_74; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_75 = mau_6_io_pipe_phv_out_data_75; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_76 = mau_6_io_pipe_phv_out_data_76; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_77 = mau_6_io_pipe_phv_out_data_77; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_78 = mau_6_io_pipe_phv_out_data_78; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_79 = mau_6_io_pipe_phv_out_data_79; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_80 = mau_6_io_pipe_phv_out_data_80; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_81 = mau_6_io_pipe_phv_out_data_81; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_82 = mau_6_io_pipe_phv_out_data_82; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_83 = mau_6_io_pipe_phv_out_data_83; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_84 = mau_6_io_pipe_phv_out_data_84; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_85 = mau_6_io_pipe_phv_out_data_85; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_86 = mau_6_io_pipe_phv_out_data_86; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_87 = mau_6_io_pipe_phv_out_data_87; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_88 = mau_6_io_pipe_phv_out_data_88; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_89 = mau_6_io_pipe_phv_out_data_89; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_90 = mau_6_io_pipe_phv_out_data_90; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_91 = mau_6_io_pipe_phv_out_data_91; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_92 = mau_6_io_pipe_phv_out_data_92; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_93 = mau_6_io_pipe_phv_out_data_93; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_94 = mau_6_io_pipe_phv_out_data_94; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_95 = mau_6_io_pipe_phv_out_data_95; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_96 = mau_6_io_pipe_phv_out_data_96; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_97 = mau_6_io_pipe_phv_out_data_97; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_98 = mau_6_io_pipe_phv_out_data_98; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_99 = mau_6_io_pipe_phv_out_data_99; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_100 = mau_6_io_pipe_phv_out_data_100; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_101 = mau_6_io_pipe_phv_out_data_101; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_102 = mau_6_io_pipe_phv_out_data_102; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_103 = mau_6_io_pipe_phv_out_data_103; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_104 = mau_6_io_pipe_phv_out_data_104; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_105 = mau_6_io_pipe_phv_out_data_105; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_106 = mau_6_io_pipe_phv_out_data_106; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_107 = mau_6_io_pipe_phv_out_data_107; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_108 = mau_6_io_pipe_phv_out_data_108; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_109 = mau_6_io_pipe_phv_out_data_109; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_110 = mau_6_io_pipe_phv_out_data_110; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_111 = mau_6_io_pipe_phv_out_data_111; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_112 = mau_6_io_pipe_phv_out_data_112; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_113 = mau_6_io_pipe_phv_out_data_113; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_114 = mau_6_io_pipe_phv_out_data_114; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_115 = mau_6_io_pipe_phv_out_data_115; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_116 = mau_6_io_pipe_phv_out_data_116; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_117 = mau_6_io_pipe_phv_out_data_117; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_118 = mau_6_io_pipe_phv_out_data_118; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_119 = mau_6_io_pipe_phv_out_data_119; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_120 = mau_6_io_pipe_phv_out_data_120; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_121 = mau_6_io_pipe_phv_out_data_121; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_122 = mau_6_io_pipe_phv_out_data_122; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_123 = mau_6_io_pipe_phv_out_data_123; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_124 = mau_6_io_pipe_phv_out_data_124; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_125 = mau_6_io_pipe_phv_out_data_125; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_126 = mau_6_io_pipe_phv_out_data_126; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_127 = mau_6_io_pipe_phv_out_data_127; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_128 = mau_6_io_pipe_phv_out_data_128; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_129 = mau_6_io_pipe_phv_out_data_129; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_130 = mau_6_io_pipe_phv_out_data_130; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_131 = mau_6_io_pipe_phv_out_data_131; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_132 = mau_6_io_pipe_phv_out_data_132; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_133 = mau_6_io_pipe_phv_out_data_133; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_134 = mau_6_io_pipe_phv_out_data_134; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_135 = mau_6_io_pipe_phv_out_data_135; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_136 = mau_6_io_pipe_phv_out_data_136; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_137 = mau_6_io_pipe_phv_out_data_137; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_138 = mau_6_io_pipe_phv_out_data_138; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_139 = mau_6_io_pipe_phv_out_data_139; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_140 = mau_6_io_pipe_phv_out_data_140; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_141 = mau_6_io_pipe_phv_out_data_141; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_142 = mau_6_io_pipe_phv_out_data_142; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_143 = mau_6_io_pipe_phv_out_data_143; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_144 = mau_6_io_pipe_phv_out_data_144; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_145 = mau_6_io_pipe_phv_out_data_145; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_146 = mau_6_io_pipe_phv_out_data_146; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_147 = mau_6_io_pipe_phv_out_data_147; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_148 = mau_6_io_pipe_phv_out_data_148; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_149 = mau_6_io_pipe_phv_out_data_149; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_150 = mau_6_io_pipe_phv_out_data_150; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_151 = mau_6_io_pipe_phv_out_data_151; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_152 = mau_6_io_pipe_phv_out_data_152; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_153 = mau_6_io_pipe_phv_out_data_153; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_154 = mau_6_io_pipe_phv_out_data_154; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_155 = mau_6_io_pipe_phv_out_data_155; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_156 = mau_6_io_pipe_phv_out_data_156; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_157 = mau_6_io_pipe_phv_out_data_157; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_158 = mau_6_io_pipe_phv_out_data_158; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_159 = mau_6_io_pipe_phv_out_data_159; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_160 = mau_6_io_pipe_phv_out_data_160; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_161 = mau_6_io_pipe_phv_out_data_161; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_162 = mau_6_io_pipe_phv_out_data_162; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_163 = mau_6_io_pipe_phv_out_data_163; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_164 = mau_6_io_pipe_phv_out_data_164; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_165 = mau_6_io_pipe_phv_out_data_165; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_166 = mau_6_io_pipe_phv_out_data_166; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_167 = mau_6_io_pipe_phv_out_data_167; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_168 = mau_6_io_pipe_phv_out_data_168; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_169 = mau_6_io_pipe_phv_out_data_169; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_170 = mau_6_io_pipe_phv_out_data_170; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_171 = mau_6_io_pipe_phv_out_data_171; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_172 = mau_6_io_pipe_phv_out_data_172; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_173 = mau_6_io_pipe_phv_out_data_173; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_174 = mau_6_io_pipe_phv_out_data_174; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_175 = mau_6_io_pipe_phv_out_data_175; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_176 = mau_6_io_pipe_phv_out_data_176; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_177 = mau_6_io_pipe_phv_out_data_177; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_178 = mau_6_io_pipe_phv_out_data_178; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_179 = mau_6_io_pipe_phv_out_data_179; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_180 = mau_6_io_pipe_phv_out_data_180; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_181 = mau_6_io_pipe_phv_out_data_181; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_182 = mau_6_io_pipe_phv_out_data_182; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_183 = mau_6_io_pipe_phv_out_data_183; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_184 = mau_6_io_pipe_phv_out_data_184; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_185 = mau_6_io_pipe_phv_out_data_185; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_186 = mau_6_io_pipe_phv_out_data_186; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_187 = mau_6_io_pipe_phv_out_data_187; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_188 = mau_6_io_pipe_phv_out_data_188; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_189 = mau_6_io_pipe_phv_out_data_189; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_190 = mau_6_io_pipe_phv_out_data_190; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_191 = mau_6_io_pipe_phv_out_data_191; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_192 = mau_6_io_pipe_phv_out_data_192; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_193 = mau_6_io_pipe_phv_out_data_193; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_194 = mau_6_io_pipe_phv_out_data_194; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_195 = mau_6_io_pipe_phv_out_data_195; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_196 = mau_6_io_pipe_phv_out_data_196; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_197 = mau_6_io_pipe_phv_out_data_197; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_198 = mau_6_io_pipe_phv_out_data_198; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_199 = mau_6_io_pipe_phv_out_data_199; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_200 = mau_6_io_pipe_phv_out_data_200; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_201 = mau_6_io_pipe_phv_out_data_201; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_202 = mau_6_io_pipe_phv_out_data_202; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_203 = mau_6_io_pipe_phv_out_data_203; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_204 = mau_6_io_pipe_phv_out_data_204; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_205 = mau_6_io_pipe_phv_out_data_205; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_206 = mau_6_io_pipe_phv_out_data_206; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_207 = mau_6_io_pipe_phv_out_data_207; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_208 = mau_6_io_pipe_phv_out_data_208; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_209 = mau_6_io_pipe_phv_out_data_209; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_210 = mau_6_io_pipe_phv_out_data_210; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_211 = mau_6_io_pipe_phv_out_data_211; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_212 = mau_6_io_pipe_phv_out_data_212; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_213 = mau_6_io_pipe_phv_out_data_213; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_214 = mau_6_io_pipe_phv_out_data_214; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_215 = mau_6_io_pipe_phv_out_data_215; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_216 = mau_6_io_pipe_phv_out_data_216; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_217 = mau_6_io_pipe_phv_out_data_217; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_218 = mau_6_io_pipe_phv_out_data_218; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_219 = mau_6_io_pipe_phv_out_data_219; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_220 = mau_6_io_pipe_phv_out_data_220; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_221 = mau_6_io_pipe_phv_out_data_221; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_222 = mau_6_io_pipe_phv_out_data_222; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_223 = mau_6_io_pipe_phv_out_data_223; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_224 = mau_6_io_pipe_phv_out_data_224; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_225 = mau_6_io_pipe_phv_out_data_225; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_226 = mau_6_io_pipe_phv_out_data_226; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_227 = mau_6_io_pipe_phv_out_data_227; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_228 = mau_6_io_pipe_phv_out_data_228; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_229 = mau_6_io_pipe_phv_out_data_229; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_230 = mau_6_io_pipe_phv_out_data_230; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_231 = mau_6_io_pipe_phv_out_data_231; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_232 = mau_6_io_pipe_phv_out_data_232; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_233 = mau_6_io_pipe_phv_out_data_233; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_234 = mau_6_io_pipe_phv_out_data_234; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_235 = mau_6_io_pipe_phv_out_data_235; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_236 = mau_6_io_pipe_phv_out_data_236; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_237 = mau_6_io_pipe_phv_out_data_237; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_238 = mau_6_io_pipe_phv_out_data_238; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_239 = mau_6_io_pipe_phv_out_data_239; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_240 = mau_6_io_pipe_phv_out_data_240; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_241 = mau_6_io_pipe_phv_out_data_241; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_242 = mau_6_io_pipe_phv_out_data_242; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_243 = mau_6_io_pipe_phv_out_data_243; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_244 = mau_6_io_pipe_phv_out_data_244; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_245 = mau_6_io_pipe_phv_out_data_245; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_246 = mau_6_io_pipe_phv_out_data_246; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_247 = mau_6_io_pipe_phv_out_data_247; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_248 = mau_6_io_pipe_phv_out_data_248; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_249 = mau_6_io_pipe_phv_out_data_249; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_250 = mau_6_io_pipe_phv_out_data_250; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_251 = mau_6_io_pipe_phv_out_data_251; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_252 = mau_6_io_pipe_phv_out_data_252; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_253 = mau_6_io_pipe_phv_out_data_253; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_254 = mau_6_io_pipe_phv_out_data_254; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_255 = mau_6_io_pipe_phv_out_data_255; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_256 = mau_6_io_pipe_phv_out_data_256; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_257 = mau_6_io_pipe_phv_out_data_257; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_258 = mau_6_io_pipe_phv_out_data_258; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_259 = mau_6_io_pipe_phv_out_data_259; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_260 = mau_6_io_pipe_phv_out_data_260; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_261 = mau_6_io_pipe_phv_out_data_261; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_262 = mau_6_io_pipe_phv_out_data_262; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_263 = mau_6_io_pipe_phv_out_data_263; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_264 = mau_6_io_pipe_phv_out_data_264; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_265 = mau_6_io_pipe_phv_out_data_265; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_266 = mau_6_io_pipe_phv_out_data_266; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_267 = mau_6_io_pipe_phv_out_data_267; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_268 = mau_6_io_pipe_phv_out_data_268; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_269 = mau_6_io_pipe_phv_out_data_269; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_270 = mau_6_io_pipe_phv_out_data_270; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_271 = mau_6_io_pipe_phv_out_data_271; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_272 = mau_6_io_pipe_phv_out_data_272; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_273 = mau_6_io_pipe_phv_out_data_273; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_274 = mau_6_io_pipe_phv_out_data_274; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_275 = mau_6_io_pipe_phv_out_data_275; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_276 = mau_6_io_pipe_phv_out_data_276; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_277 = mau_6_io_pipe_phv_out_data_277; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_278 = mau_6_io_pipe_phv_out_data_278; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_279 = mau_6_io_pipe_phv_out_data_279; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_280 = mau_6_io_pipe_phv_out_data_280; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_281 = mau_6_io_pipe_phv_out_data_281; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_282 = mau_6_io_pipe_phv_out_data_282; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_283 = mau_6_io_pipe_phv_out_data_283; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_284 = mau_6_io_pipe_phv_out_data_284; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_285 = mau_6_io_pipe_phv_out_data_285; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_286 = mau_6_io_pipe_phv_out_data_286; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_287 = mau_6_io_pipe_phv_out_data_287; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_288 = mau_6_io_pipe_phv_out_data_288; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_289 = mau_6_io_pipe_phv_out_data_289; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_290 = mau_6_io_pipe_phv_out_data_290; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_291 = mau_6_io_pipe_phv_out_data_291; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_292 = mau_6_io_pipe_phv_out_data_292; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_293 = mau_6_io_pipe_phv_out_data_293; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_294 = mau_6_io_pipe_phv_out_data_294; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_295 = mau_6_io_pipe_phv_out_data_295; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_296 = mau_6_io_pipe_phv_out_data_296; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_297 = mau_6_io_pipe_phv_out_data_297; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_298 = mau_6_io_pipe_phv_out_data_298; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_299 = mau_6_io_pipe_phv_out_data_299; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_300 = mau_6_io_pipe_phv_out_data_300; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_301 = mau_6_io_pipe_phv_out_data_301; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_302 = mau_6_io_pipe_phv_out_data_302; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_303 = mau_6_io_pipe_phv_out_data_303; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_304 = mau_6_io_pipe_phv_out_data_304; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_305 = mau_6_io_pipe_phv_out_data_305; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_306 = mau_6_io_pipe_phv_out_data_306; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_307 = mau_6_io_pipe_phv_out_data_307; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_308 = mau_6_io_pipe_phv_out_data_308; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_309 = mau_6_io_pipe_phv_out_data_309; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_310 = mau_6_io_pipe_phv_out_data_310; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_311 = mau_6_io_pipe_phv_out_data_311; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_312 = mau_6_io_pipe_phv_out_data_312; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_313 = mau_6_io_pipe_phv_out_data_313; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_314 = mau_6_io_pipe_phv_out_data_314; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_315 = mau_6_io_pipe_phv_out_data_315; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_316 = mau_6_io_pipe_phv_out_data_316; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_317 = mau_6_io_pipe_phv_out_data_317; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_318 = mau_6_io_pipe_phv_out_data_318; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_319 = mau_6_io_pipe_phv_out_data_319; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_320 = mau_6_io_pipe_phv_out_data_320; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_321 = mau_6_io_pipe_phv_out_data_321; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_322 = mau_6_io_pipe_phv_out_data_322; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_323 = mau_6_io_pipe_phv_out_data_323; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_324 = mau_6_io_pipe_phv_out_data_324; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_325 = mau_6_io_pipe_phv_out_data_325; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_326 = mau_6_io_pipe_phv_out_data_326; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_327 = mau_6_io_pipe_phv_out_data_327; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_328 = mau_6_io_pipe_phv_out_data_328; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_329 = mau_6_io_pipe_phv_out_data_329; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_330 = mau_6_io_pipe_phv_out_data_330; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_331 = mau_6_io_pipe_phv_out_data_331; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_332 = mau_6_io_pipe_phv_out_data_332; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_333 = mau_6_io_pipe_phv_out_data_333; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_334 = mau_6_io_pipe_phv_out_data_334; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_335 = mau_6_io_pipe_phv_out_data_335; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_336 = mau_6_io_pipe_phv_out_data_336; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_337 = mau_6_io_pipe_phv_out_data_337; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_338 = mau_6_io_pipe_phv_out_data_338; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_339 = mau_6_io_pipe_phv_out_data_339; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_340 = mau_6_io_pipe_phv_out_data_340; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_341 = mau_6_io_pipe_phv_out_data_341; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_342 = mau_6_io_pipe_phv_out_data_342; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_343 = mau_6_io_pipe_phv_out_data_343; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_344 = mau_6_io_pipe_phv_out_data_344; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_345 = mau_6_io_pipe_phv_out_data_345; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_346 = mau_6_io_pipe_phv_out_data_346; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_347 = mau_6_io_pipe_phv_out_data_347; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_348 = mau_6_io_pipe_phv_out_data_348; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_349 = mau_6_io_pipe_phv_out_data_349; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_350 = mau_6_io_pipe_phv_out_data_350; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_351 = mau_6_io_pipe_phv_out_data_351; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_352 = mau_6_io_pipe_phv_out_data_352; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_353 = mau_6_io_pipe_phv_out_data_353; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_354 = mau_6_io_pipe_phv_out_data_354; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_355 = mau_6_io_pipe_phv_out_data_355; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_356 = mau_6_io_pipe_phv_out_data_356; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_357 = mau_6_io_pipe_phv_out_data_357; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_358 = mau_6_io_pipe_phv_out_data_358; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_359 = mau_6_io_pipe_phv_out_data_359; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_360 = mau_6_io_pipe_phv_out_data_360; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_361 = mau_6_io_pipe_phv_out_data_361; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_362 = mau_6_io_pipe_phv_out_data_362; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_363 = mau_6_io_pipe_phv_out_data_363; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_364 = mau_6_io_pipe_phv_out_data_364; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_365 = mau_6_io_pipe_phv_out_data_365; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_366 = mau_6_io_pipe_phv_out_data_366; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_367 = mau_6_io_pipe_phv_out_data_367; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_368 = mau_6_io_pipe_phv_out_data_368; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_369 = mau_6_io_pipe_phv_out_data_369; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_370 = mau_6_io_pipe_phv_out_data_370; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_371 = mau_6_io_pipe_phv_out_data_371; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_372 = mau_6_io_pipe_phv_out_data_372; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_373 = mau_6_io_pipe_phv_out_data_373; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_374 = mau_6_io_pipe_phv_out_data_374; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_375 = mau_6_io_pipe_phv_out_data_375; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_376 = mau_6_io_pipe_phv_out_data_376; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_377 = mau_6_io_pipe_phv_out_data_377; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_378 = mau_6_io_pipe_phv_out_data_378; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_379 = mau_6_io_pipe_phv_out_data_379; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_380 = mau_6_io_pipe_phv_out_data_380; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_381 = mau_6_io_pipe_phv_out_data_381; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_382 = mau_6_io_pipe_phv_out_data_382; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_383 = mau_6_io_pipe_phv_out_data_383; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_384 = mau_6_io_pipe_phv_out_data_384; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_385 = mau_6_io_pipe_phv_out_data_385; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_386 = mau_6_io_pipe_phv_out_data_386; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_387 = mau_6_io_pipe_phv_out_data_387; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_388 = mau_6_io_pipe_phv_out_data_388; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_389 = mau_6_io_pipe_phv_out_data_389; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_390 = mau_6_io_pipe_phv_out_data_390; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_391 = mau_6_io_pipe_phv_out_data_391; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_392 = mau_6_io_pipe_phv_out_data_392; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_393 = mau_6_io_pipe_phv_out_data_393; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_394 = mau_6_io_pipe_phv_out_data_394; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_395 = mau_6_io_pipe_phv_out_data_395; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_396 = mau_6_io_pipe_phv_out_data_396; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_397 = mau_6_io_pipe_phv_out_data_397; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_398 = mau_6_io_pipe_phv_out_data_398; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_399 = mau_6_io_pipe_phv_out_data_399; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_400 = mau_6_io_pipe_phv_out_data_400; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_401 = mau_6_io_pipe_phv_out_data_401; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_402 = mau_6_io_pipe_phv_out_data_402; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_403 = mau_6_io_pipe_phv_out_data_403; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_404 = mau_6_io_pipe_phv_out_data_404; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_405 = mau_6_io_pipe_phv_out_data_405; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_406 = mau_6_io_pipe_phv_out_data_406; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_407 = mau_6_io_pipe_phv_out_data_407; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_408 = mau_6_io_pipe_phv_out_data_408; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_409 = mau_6_io_pipe_phv_out_data_409; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_410 = mau_6_io_pipe_phv_out_data_410; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_411 = mau_6_io_pipe_phv_out_data_411; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_412 = mau_6_io_pipe_phv_out_data_412; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_413 = mau_6_io_pipe_phv_out_data_413; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_414 = mau_6_io_pipe_phv_out_data_414; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_415 = mau_6_io_pipe_phv_out_data_415; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_416 = mau_6_io_pipe_phv_out_data_416; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_417 = mau_6_io_pipe_phv_out_data_417; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_418 = mau_6_io_pipe_phv_out_data_418; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_419 = mau_6_io_pipe_phv_out_data_419; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_420 = mau_6_io_pipe_phv_out_data_420; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_421 = mau_6_io_pipe_phv_out_data_421; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_422 = mau_6_io_pipe_phv_out_data_422; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_423 = mau_6_io_pipe_phv_out_data_423; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_424 = mau_6_io_pipe_phv_out_data_424; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_425 = mau_6_io_pipe_phv_out_data_425; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_426 = mau_6_io_pipe_phv_out_data_426; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_427 = mau_6_io_pipe_phv_out_data_427; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_428 = mau_6_io_pipe_phv_out_data_428; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_429 = mau_6_io_pipe_phv_out_data_429; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_430 = mau_6_io_pipe_phv_out_data_430; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_431 = mau_6_io_pipe_phv_out_data_431; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_432 = mau_6_io_pipe_phv_out_data_432; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_433 = mau_6_io_pipe_phv_out_data_433; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_434 = mau_6_io_pipe_phv_out_data_434; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_435 = mau_6_io_pipe_phv_out_data_435; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_436 = mau_6_io_pipe_phv_out_data_436; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_437 = mau_6_io_pipe_phv_out_data_437; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_438 = mau_6_io_pipe_phv_out_data_438; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_439 = mau_6_io_pipe_phv_out_data_439; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_440 = mau_6_io_pipe_phv_out_data_440; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_441 = mau_6_io_pipe_phv_out_data_441; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_442 = mau_6_io_pipe_phv_out_data_442; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_443 = mau_6_io_pipe_phv_out_data_443; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_444 = mau_6_io_pipe_phv_out_data_444; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_445 = mau_6_io_pipe_phv_out_data_445; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_446 = mau_6_io_pipe_phv_out_data_446; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_447 = mau_6_io_pipe_phv_out_data_447; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_448 = mau_6_io_pipe_phv_out_data_448; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_449 = mau_6_io_pipe_phv_out_data_449; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_450 = mau_6_io_pipe_phv_out_data_450; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_451 = mau_6_io_pipe_phv_out_data_451; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_452 = mau_6_io_pipe_phv_out_data_452; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_453 = mau_6_io_pipe_phv_out_data_453; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_454 = mau_6_io_pipe_phv_out_data_454; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_455 = mau_6_io_pipe_phv_out_data_455; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_456 = mau_6_io_pipe_phv_out_data_456; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_457 = mau_6_io_pipe_phv_out_data_457; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_458 = mau_6_io_pipe_phv_out_data_458; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_459 = mau_6_io_pipe_phv_out_data_459; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_460 = mau_6_io_pipe_phv_out_data_460; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_461 = mau_6_io_pipe_phv_out_data_461; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_462 = mau_6_io_pipe_phv_out_data_462; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_463 = mau_6_io_pipe_phv_out_data_463; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_464 = mau_6_io_pipe_phv_out_data_464; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_465 = mau_6_io_pipe_phv_out_data_465; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_466 = mau_6_io_pipe_phv_out_data_466; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_467 = mau_6_io_pipe_phv_out_data_467; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_468 = mau_6_io_pipe_phv_out_data_468; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_469 = mau_6_io_pipe_phv_out_data_469; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_470 = mau_6_io_pipe_phv_out_data_470; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_471 = mau_6_io_pipe_phv_out_data_471; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_472 = mau_6_io_pipe_phv_out_data_472; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_473 = mau_6_io_pipe_phv_out_data_473; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_474 = mau_6_io_pipe_phv_out_data_474; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_475 = mau_6_io_pipe_phv_out_data_475; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_476 = mau_6_io_pipe_phv_out_data_476; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_477 = mau_6_io_pipe_phv_out_data_477; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_478 = mau_6_io_pipe_phv_out_data_478; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_479 = mau_6_io_pipe_phv_out_data_479; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_480 = mau_6_io_pipe_phv_out_data_480; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_481 = mau_6_io_pipe_phv_out_data_481; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_482 = mau_6_io_pipe_phv_out_data_482; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_483 = mau_6_io_pipe_phv_out_data_483; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_484 = mau_6_io_pipe_phv_out_data_484; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_485 = mau_6_io_pipe_phv_out_data_485; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_486 = mau_6_io_pipe_phv_out_data_486; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_487 = mau_6_io_pipe_phv_out_data_487; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_488 = mau_6_io_pipe_phv_out_data_488; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_489 = mau_6_io_pipe_phv_out_data_489; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_490 = mau_6_io_pipe_phv_out_data_490; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_491 = mau_6_io_pipe_phv_out_data_491; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_492 = mau_6_io_pipe_phv_out_data_492; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_493 = mau_6_io_pipe_phv_out_data_493; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_494 = mau_6_io_pipe_phv_out_data_494; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_495 = mau_6_io_pipe_phv_out_data_495; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_496 = mau_6_io_pipe_phv_out_data_496; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_497 = mau_6_io_pipe_phv_out_data_497; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_498 = mau_6_io_pipe_phv_out_data_498; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_499 = mau_6_io_pipe_phv_out_data_499; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_500 = mau_6_io_pipe_phv_out_data_500; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_501 = mau_6_io_pipe_phv_out_data_501; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_502 = mau_6_io_pipe_phv_out_data_502; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_503 = mau_6_io_pipe_phv_out_data_503; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_504 = mau_6_io_pipe_phv_out_data_504; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_505 = mau_6_io_pipe_phv_out_data_505; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_506 = mau_6_io_pipe_phv_out_data_506; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_507 = mau_6_io_pipe_phv_out_data_507; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_508 = mau_6_io_pipe_phv_out_data_508; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_509 = mau_6_io_pipe_phv_out_data_509; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_510 = mau_6_io_pipe_phv_out_data_510; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_511 = mau_6_io_pipe_phv_out_data_511; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_header_0 = mau_6_io_pipe_phv_out_header_0; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_header_1 = mau_6_io_pipe_phv_out_header_1; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_header_2 = mau_6_io_pipe_phv_out_header_2; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_header_3 = mau_6_io_pipe_phv_out_header_3; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_header_4 = mau_6_io_pipe_phv_out_header_4; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_header_5 = mau_6_io_pipe_phv_out_header_5; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_header_6 = mau_6_io_pipe_phv_out_header_6; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_header_7 = mau_6_io_pipe_phv_out_header_7; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_header_8 = mau_6_io_pipe_phv_out_header_8; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_header_9 = mau_6_io_pipe_phv_out_header_9; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_header_10 = mau_6_io_pipe_phv_out_header_10; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_header_11 = mau_6_io_pipe_phv_out_header_11; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_header_12 = mau_6_io_pipe_phv_out_header_12; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_header_13 = mau_6_io_pipe_phv_out_header_13; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_header_14 = mau_6_io_pipe_phv_out_header_14; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_header_15 = mau_6_io_pipe_phv_out_header_15; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_parse_current_state = mau_6_io_pipe_phv_out_parse_current_state; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_parse_current_offset = mau_6_io_pipe_phv_out_parse_current_offset; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_parse_transition_field = mau_6_io_pipe_phv_out_parse_transition_field; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_next_processor_id = mau_6_io_pipe_phv_out_next_processor_id; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_next_config_id = mau_6_io_pipe_phv_out_next_config_id; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_is_valid_processor = mau_6_io_pipe_phv_out_is_valid_processor; // @[parser_pisa.scala 42:35]
  assign mau_7_io_mod_state_id_mod = io_mod_en ? io_mod_module_mod_state_id_mod & mod_j_7 :
    io_mod_module_mod_state_id_mod; // @[parser_pisa.scala 51:22 parser_pisa.scala 58:40 parser_pisa.scala 47:23]
  assign mau_7_io_mod_state_id = io_mod_module_mod_state_id; // @[parser_pisa.scala 47:23]
  assign mau_7_io_mod_sram_w_cs = io_mod_module_mod_sram_w_cs; // @[parser_pisa.scala 47:23]
  assign mau_7_io_mod_sram_w_en = io_mod_en ? io_mod_module_mod_sram_w_en & mod_j_7 : io_mod_module_mod_sram_w_en; // @[parser_pisa.scala 51:22 parser_pisa.scala 57:40 parser_pisa.scala 47:23]
  assign mau_7_io_mod_sram_w_addr = io_mod_module_mod_sram_w_addr; // @[parser_pisa.scala 47:23]
  assign mau_7_io_mod_sram_w_data = io_mod_module_mod_sram_w_data; // @[parser_pisa.scala 47:23]
  always @(posedge clock) begin
    if (io_mod_en) begin // @[parser_pisa.scala 51:22]
      if (io_mod_last_mau_id_mod) begin // @[parser_pisa.scala 52:39]
        last_mau_id <= io_mod_last_mau_id; // @[parser_pisa.scala 53:25]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  last_mau_id = _RAND_0[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
