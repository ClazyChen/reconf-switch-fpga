module PrimitiveWriteBack(
  input         clock,
  input  [7:0]  io_pipe_phv_in_data_0,
  input  [7:0]  io_pipe_phv_in_data_1,
  input  [7:0]  io_pipe_phv_in_data_2,
  input  [7:0]  io_pipe_phv_in_data_3,
  input  [7:0]  io_pipe_phv_in_data_4,
  input  [7:0]  io_pipe_phv_in_data_5,
  input  [7:0]  io_pipe_phv_in_data_6,
  input  [7:0]  io_pipe_phv_in_data_7,
  input  [7:0]  io_pipe_phv_in_data_8,
  input  [7:0]  io_pipe_phv_in_data_9,
  input  [7:0]  io_pipe_phv_in_data_10,
  input  [7:0]  io_pipe_phv_in_data_11,
  input  [7:0]  io_pipe_phv_in_data_12,
  input  [7:0]  io_pipe_phv_in_data_13,
  input  [7:0]  io_pipe_phv_in_data_14,
  input  [7:0]  io_pipe_phv_in_data_15,
  input  [7:0]  io_pipe_phv_in_data_16,
  input  [7:0]  io_pipe_phv_in_data_17,
  input  [7:0]  io_pipe_phv_in_data_18,
  input  [7:0]  io_pipe_phv_in_data_19,
  input  [7:0]  io_pipe_phv_in_data_20,
  input  [7:0]  io_pipe_phv_in_data_21,
  input  [7:0]  io_pipe_phv_in_data_22,
  input  [7:0]  io_pipe_phv_in_data_23,
  input  [7:0]  io_pipe_phv_in_data_24,
  input  [7:0]  io_pipe_phv_in_data_25,
  input  [7:0]  io_pipe_phv_in_data_26,
  input  [7:0]  io_pipe_phv_in_data_27,
  input  [7:0]  io_pipe_phv_in_data_28,
  input  [7:0]  io_pipe_phv_in_data_29,
  input  [7:0]  io_pipe_phv_in_data_30,
  input  [7:0]  io_pipe_phv_in_data_31,
  input  [7:0]  io_pipe_phv_in_data_32,
  input  [7:0]  io_pipe_phv_in_data_33,
  input  [7:0]  io_pipe_phv_in_data_34,
  input  [7:0]  io_pipe_phv_in_data_35,
  input  [7:0]  io_pipe_phv_in_data_36,
  input  [7:0]  io_pipe_phv_in_data_37,
  input  [7:0]  io_pipe_phv_in_data_38,
  input  [7:0]  io_pipe_phv_in_data_39,
  input  [7:0]  io_pipe_phv_in_data_40,
  input  [7:0]  io_pipe_phv_in_data_41,
  input  [7:0]  io_pipe_phv_in_data_42,
  input  [7:0]  io_pipe_phv_in_data_43,
  input  [7:0]  io_pipe_phv_in_data_44,
  input  [7:0]  io_pipe_phv_in_data_45,
  input  [7:0]  io_pipe_phv_in_data_46,
  input  [7:0]  io_pipe_phv_in_data_47,
  input  [7:0]  io_pipe_phv_in_data_48,
  input  [7:0]  io_pipe_phv_in_data_49,
  input  [7:0]  io_pipe_phv_in_data_50,
  input  [7:0]  io_pipe_phv_in_data_51,
  input  [7:0]  io_pipe_phv_in_data_52,
  input  [7:0]  io_pipe_phv_in_data_53,
  input  [7:0]  io_pipe_phv_in_data_54,
  input  [7:0]  io_pipe_phv_in_data_55,
  input  [7:0]  io_pipe_phv_in_data_56,
  input  [7:0]  io_pipe_phv_in_data_57,
  input  [7:0]  io_pipe_phv_in_data_58,
  input  [7:0]  io_pipe_phv_in_data_59,
  input  [7:0]  io_pipe_phv_in_data_60,
  input  [7:0]  io_pipe_phv_in_data_61,
  input  [7:0]  io_pipe_phv_in_data_62,
  input  [7:0]  io_pipe_phv_in_data_63,
  input  [7:0]  io_pipe_phv_in_data_64,
  input  [7:0]  io_pipe_phv_in_data_65,
  input  [7:0]  io_pipe_phv_in_data_66,
  input  [7:0]  io_pipe_phv_in_data_67,
  input  [7:0]  io_pipe_phv_in_data_68,
  input  [7:0]  io_pipe_phv_in_data_69,
  input  [7:0]  io_pipe_phv_in_data_70,
  input  [7:0]  io_pipe_phv_in_data_71,
  input  [7:0]  io_pipe_phv_in_data_72,
  input  [7:0]  io_pipe_phv_in_data_73,
  input  [7:0]  io_pipe_phv_in_data_74,
  input  [7:0]  io_pipe_phv_in_data_75,
  input  [7:0]  io_pipe_phv_in_data_76,
  input  [7:0]  io_pipe_phv_in_data_77,
  input  [7:0]  io_pipe_phv_in_data_78,
  input  [7:0]  io_pipe_phv_in_data_79,
  input  [7:0]  io_pipe_phv_in_data_80,
  input  [7:0]  io_pipe_phv_in_data_81,
  input  [7:0]  io_pipe_phv_in_data_82,
  input  [7:0]  io_pipe_phv_in_data_83,
  input  [7:0]  io_pipe_phv_in_data_84,
  input  [7:0]  io_pipe_phv_in_data_85,
  input  [7:0]  io_pipe_phv_in_data_86,
  input  [7:0]  io_pipe_phv_in_data_87,
  input  [7:0]  io_pipe_phv_in_data_88,
  input  [7:0]  io_pipe_phv_in_data_89,
  input  [7:0]  io_pipe_phv_in_data_90,
  input  [7:0]  io_pipe_phv_in_data_91,
  input  [7:0]  io_pipe_phv_in_data_92,
  input  [7:0]  io_pipe_phv_in_data_93,
  input  [7:0]  io_pipe_phv_in_data_94,
  input  [7:0]  io_pipe_phv_in_data_95,
  input  [7:0]  io_pipe_phv_in_data_96,
  input  [7:0]  io_pipe_phv_in_data_97,
  input  [7:0]  io_pipe_phv_in_data_98,
  input  [7:0]  io_pipe_phv_in_data_99,
  input  [7:0]  io_pipe_phv_in_data_100,
  input  [7:0]  io_pipe_phv_in_data_101,
  input  [7:0]  io_pipe_phv_in_data_102,
  input  [7:0]  io_pipe_phv_in_data_103,
  input  [7:0]  io_pipe_phv_in_data_104,
  input  [7:0]  io_pipe_phv_in_data_105,
  input  [7:0]  io_pipe_phv_in_data_106,
  input  [7:0]  io_pipe_phv_in_data_107,
  input  [7:0]  io_pipe_phv_in_data_108,
  input  [7:0]  io_pipe_phv_in_data_109,
  input  [7:0]  io_pipe_phv_in_data_110,
  input  [7:0]  io_pipe_phv_in_data_111,
  input  [7:0]  io_pipe_phv_in_data_112,
  input  [7:0]  io_pipe_phv_in_data_113,
  input  [7:0]  io_pipe_phv_in_data_114,
  input  [7:0]  io_pipe_phv_in_data_115,
  input  [7:0]  io_pipe_phv_in_data_116,
  input  [7:0]  io_pipe_phv_in_data_117,
  input  [7:0]  io_pipe_phv_in_data_118,
  input  [7:0]  io_pipe_phv_in_data_119,
  input  [7:0]  io_pipe_phv_in_data_120,
  input  [7:0]  io_pipe_phv_in_data_121,
  input  [7:0]  io_pipe_phv_in_data_122,
  input  [7:0]  io_pipe_phv_in_data_123,
  input  [7:0]  io_pipe_phv_in_data_124,
  input  [7:0]  io_pipe_phv_in_data_125,
  input  [7:0]  io_pipe_phv_in_data_126,
  input  [7:0]  io_pipe_phv_in_data_127,
  input  [7:0]  io_pipe_phv_in_data_128,
  input  [7:0]  io_pipe_phv_in_data_129,
  input  [7:0]  io_pipe_phv_in_data_130,
  input  [7:0]  io_pipe_phv_in_data_131,
  input  [7:0]  io_pipe_phv_in_data_132,
  input  [7:0]  io_pipe_phv_in_data_133,
  input  [7:0]  io_pipe_phv_in_data_134,
  input  [7:0]  io_pipe_phv_in_data_135,
  input  [7:0]  io_pipe_phv_in_data_136,
  input  [7:0]  io_pipe_phv_in_data_137,
  input  [7:0]  io_pipe_phv_in_data_138,
  input  [7:0]  io_pipe_phv_in_data_139,
  input  [7:0]  io_pipe_phv_in_data_140,
  input  [7:0]  io_pipe_phv_in_data_141,
  input  [7:0]  io_pipe_phv_in_data_142,
  input  [7:0]  io_pipe_phv_in_data_143,
  input  [7:0]  io_pipe_phv_in_data_144,
  input  [7:0]  io_pipe_phv_in_data_145,
  input  [7:0]  io_pipe_phv_in_data_146,
  input  [7:0]  io_pipe_phv_in_data_147,
  input  [7:0]  io_pipe_phv_in_data_148,
  input  [7:0]  io_pipe_phv_in_data_149,
  input  [7:0]  io_pipe_phv_in_data_150,
  input  [7:0]  io_pipe_phv_in_data_151,
  input  [7:0]  io_pipe_phv_in_data_152,
  input  [7:0]  io_pipe_phv_in_data_153,
  input  [7:0]  io_pipe_phv_in_data_154,
  input  [7:0]  io_pipe_phv_in_data_155,
  input  [7:0]  io_pipe_phv_in_data_156,
  input  [7:0]  io_pipe_phv_in_data_157,
  input  [7:0]  io_pipe_phv_in_data_158,
  input  [7:0]  io_pipe_phv_in_data_159,
  input  [15:0] io_pipe_phv_in_header_0,
  input  [15:0] io_pipe_phv_in_header_1,
  input  [15:0] io_pipe_phv_in_header_2,
  input  [15:0] io_pipe_phv_in_header_3,
  input  [15:0] io_pipe_phv_in_header_4,
  input  [15:0] io_pipe_phv_in_header_5,
  input  [15:0] io_pipe_phv_in_header_6,
  input  [15:0] io_pipe_phv_in_header_7,
  input  [15:0] io_pipe_phv_in_header_8,
  input  [15:0] io_pipe_phv_in_header_9,
  input  [15:0] io_pipe_phv_in_header_10,
  input  [15:0] io_pipe_phv_in_header_11,
  input  [15:0] io_pipe_phv_in_header_12,
  input  [15:0] io_pipe_phv_in_header_13,
  input  [15:0] io_pipe_phv_in_header_14,
  input  [15:0] io_pipe_phv_in_header_15,
  input  [7:0]  io_pipe_phv_in_parse_current_state,
  input  [7:0]  io_pipe_phv_in_parse_current_offset,
  input  [15:0] io_pipe_phv_in_parse_transition_field,
  input  [3:0]  io_pipe_phv_in_next_processor_id,
  input         io_pipe_phv_in_next_config_id,
  input         io_pipe_phv_in_is_valid_processor,
  output [7:0]  io_pipe_phv_out_data_0,
  output [7:0]  io_pipe_phv_out_data_1,
  output [7:0]  io_pipe_phv_out_data_2,
  output [7:0]  io_pipe_phv_out_data_3,
  output [7:0]  io_pipe_phv_out_data_4,
  output [7:0]  io_pipe_phv_out_data_5,
  output [7:0]  io_pipe_phv_out_data_6,
  output [7:0]  io_pipe_phv_out_data_7,
  output [7:0]  io_pipe_phv_out_data_8,
  output [7:0]  io_pipe_phv_out_data_9,
  output [7:0]  io_pipe_phv_out_data_10,
  output [7:0]  io_pipe_phv_out_data_11,
  output [7:0]  io_pipe_phv_out_data_12,
  output [7:0]  io_pipe_phv_out_data_13,
  output [7:0]  io_pipe_phv_out_data_14,
  output [7:0]  io_pipe_phv_out_data_15,
  output [7:0]  io_pipe_phv_out_data_16,
  output [7:0]  io_pipe_phv_out_data_17,
  output [7:0]  io_pipe_phv_out_data_18,
  output [7:0]  io_pipe_phv_out_data_19,
  output [7:0]  io_pipe_phv_out_data_20,
  output [7:0]  io_pipe_phv_out_data_21,
  output [7:0]  io_pipe_phv_out_data_22,
  output [7:0]  io_pipe_phv_out_data_23,
  output [7:0]  io_pipe_phv_out_data_24,
  output [7:0]  io_pipe_phv_out_data_25,
  output [7:0]  io_pipe_phv_out_data_26,
  output [7:0]  io_pipe_phv_out_data_27,
  output [7:0]  io_pipe_phv_out_data_28,
  output [7:0]  io_pipe_phv_out_data_29,
  output [7:0]  io_pipe_phv_out_data_30,
  output [7:0]  io_pipe_phv_out_data_31,
  output [7:0]  io_pipe_phv_out_data_32,
  output [7:0]  io_pipe_phv_out_data_33,
  output [7:0]  io_pipe_phv_out_data_34,
  output [7:0]  io_pipe_phv_out_data_35,
  output [7:0]  io_pipe_phv_out_data_36,
  output [7:0]  io_pipe_phv_out_data_37,
  output [7:0]  io_pipe_phv_out_data_38,
  output [7:0]  io_pipe_phv_out_data_39,
  output [7:0]  io_pipe_phv_out_data_40,
  output [7:0]  io_pipe_phv_out_data_41,
  output [7:0]  io_pipe_phv_out_data_42,
  output [7:0]  io_pipe_phv_out_data_43,
  output [7:0]  io_pipe_phv_out_data_44,
  output [7:0]  io_pipe_phv_out_data_45,
  output [7:0]  io_pipe_phv_out_data_46,
  output [7:0]  io_pipe_phv_out_data_47,
  output [7:0]  io_pipe_phv_out_data_48,
  output [7:0]  io_pipe_phv_out_data_49,
  output [7:0]  io_pipe_phv_out_data_50,
  output [7:0]  io_pipe_phv_out_data_51,
  output [7:0]  io_pipe_phv_out_data_52,
  output [7:0]  io_pipe_phv_out_data_53,
  output [7:0]  io_pipe_phv_out_data_54,
  output [7:0]  io_pipe_phv_out_data_55,
  output [7:0]  io_pipe_phv_out_data_56,
  output [7:0]  io_pipe_phv_out_data_57,
  output [7:0]  io_pipe_phv_out_data_58,
  output [7:0]  io_pipe_phv_out_data_59,
  output [7:0]  io_pipe_phv_out_data_60,
  output [7:0]  io_pipe_phv_out_data_61,
  output [7:0]  io_pipe_phv_out_data_62,
  output [7:0]  io_pipe_phv_out_data_63,
  output [7:0]  io_pipe_phv_out_data_64,
  output [7:0]  io_pipe_phv_out_data_65,
  output [7:0]  io_pipe_phv_out_data_66,
  output [7:0]  io_pipe_phv_out_data_67,
  output [7:0]  io_pipe_phv_out_data_68,
  output [7:0]  io_pipe_phv_out_data_69,
  output [7:0]  io_pipe_phv_out_data_70,
  output [7:0]  io_pipe_phv_out_data_71,
  output [7:0]  io_pipe_phv_out_data_72,
  output [7:0]  io_pipe_phv_out_data_73,
  output [7:0]  io_pipe_phv_out_data_74,
  output [7:0]  io_pipe_phv_out_data_75,
  output [7:0]  io_pipe_phv_out_data_76,
  output [7:0]  io_pipe_phv_out_data_77,
  output [7:0]  io_pipe_phv_out_data_78,
  output [7:0]  io_pipe_phv_out_data_79,
  output [7:0]  io_pipe_phv_out_data_80,
  output [7:0]  io_pipe_phv_out_data_81,
  output [7:0]  io_pipe_phv_out_data_82,
  output [7:0]  io_pipe_phv_out_data_83,
  output [7:0]  io_pipe_phv_out_data_84,
  output [7:0]  io_pipe_phv_out_data_85,
  output [7:0]  io_pipe_phv_out_data_86,
  output [7:0]  io_pipe_phv_out_data_87,
  output [7:0]  io_pipe_phv_out_data_88,
  output [7:0]  io_pipe_phv_out_data_89,
  output [7:0]  io_pipe_phv_out_data_90,
  output [7:0]  io_pipe_phv_out_data_91,
  output [7:0]  io_pipe_phv_out_data_92,
  output [7:0]  io_pipe_phv_out_data_93,
  output [7:0]  io_pipe_phv_out_data_94,
  output [7:0]  io_pipe_phv_out_data_95,
  output [7:0]  io_pipe_phv_out_data_96,
  output [7:0]  io_pipe_phv_out_data_97,
  output [7:0]  io_pipe_phv_out_data_98,
  output [7:0]  io_pipe_phv_out_data_99,
  output [7:0]  io_pipe_phv_out_data_100,
  output [7:0]  io_pipe_phv_out_data_101,
  output [7:0]  io_pipe_phv_out_data_102,
  output [7:0]  io_pipe_phv_out_data_103,
  output [7:0]  io_pipe_phv_out_data_104,
  output [7:0]  io_pipe_phv_out_data_105,
  output [7:0]  io_pipe_phv_out_data_106,
  output [7:0]  io_pipe_phv_out_data_107,
  output [7:0]  io_pipe_phv_out_data_108,
  output [7:0]  io_pipe_phv_out_data_109,
  output [7:0]  io_pipe_phv_out_data_110,
  output [7:0]  io_pipe_phv_out_data_111,
  output [7:0]  io_pipe_phv_out_data_112,
  output [7:0]  io_pipe_phv_out_data_113,
  output [7:0]  io_pipe_phv_out_data_114,
  output [7:0]  io_pipe_phv_out_data_115,
  output [7:0]  io_pipe_phv_out_data_116,
  output [7:0]  io_pipe_phv_out_data_117,
  output [7:0]  io_pipe_phv_out_data_118,
  output [7:0]  io_pipe_phv_out_data_119,
  output [7:0]  io_pipe_phv_out_data_120,
  output [7:0]  io_pipe_phv_out_data_121,
  output [7:0]  io_pipe_phv_out_data_122,
  output [7:0]  io_pipe_phv_out_data_123,
  output [7:0]  io_pipe_phv_out_data_124,
  output [7:0]  io_pipe_phv_out_data_125,
  output [7:0]  io_pipe_phv_out_data_126,
  output [7:0]  io_pipe_phv_out_data_127,
  output [7:0]  io_pipe_phv_out_data_128,
  output [7:0]  io_pipe_phv_out_data_129,
  output [7:0]  io_pipe_phv_out_data_130,
  output [7:0]  io_pipe_phv_out_data_131,
  output [7:0]  io_pipe_phv_out_data_132,
  output [7:0]  io_pipe_phv_out_data_133,
  output [7:0]  io_pipe_phv_out_data_134,
  output [7:0]  io_pipe_phv_out_data_135,
  output [7:0]  io_pipe_phv_out_data_136,
  output [7:0]  io_pipe_phv_out_data_137,
  output [7:0]  io_pipe_phv_out_data_138,
  output [7:0]  io_pipe_phv_out_data_139,
  output [7:0]  io_pipe_phv_out_data_140,
  output [7:0]  io_pipe_phv_out_data_141,
  output [7:0]  io_pipe_phv_out_data_142,
  output [7:0]  io_pipe_phv_out_data_143,
  output [7:0]  io_pipe_phv_out_data_144,
  output [7:0]  io_pipe_phv_out_data_145,
  output [7:0]  io_pipe_phv_out_data_146,
  output [7:0]  io_pipe_phv_out_data_147,
  output [7:0]  io_pipe_phv_out_data_148,
  output [7:0]  io_pipe_phv_out_data_149,
  output [7:0]  io_pipe_phv_out_data_150,
  output [7:0]  io_pipe_phv_out_data_151,
  output [7:0]  io_pipe_phv_out_data_152,
  output [7:0]  io_pipe_phv_out_data_153,
  output [7:0]  io_pipe_phv_out_data_154,
  output [7:0]  io_pipe_phv_out_data_155,
  output [7:0]  io_pipe_phv_out_data_156,
  output [7:0]  io_pipe_phv_out_data_157,
  output [7:0]  io_pipe_phv_out_data_158,
  output [7:0]  io_pipe_phv_out_data_159,
  output [15:0] io_pipe_phv_out_header_0,
  output [15:0] io_pipe_phv_out_header_1,
  output [15:0] io_pipe_phv_out_header_2,
  output [15:0] io_pipe_phv_out_header_3,
  output [15:0] io_pipe_phv_out_header_4,
  output [15:0] io_pipe_phv_out_header_5,
  output [15:0] io_pipe_phv_out_header_6,
  output [15:0] io_pipe_phv_out_header_7,
  output [15:0] io_pipe_phv_out_header_8,
  output [15:0] io_pipe_phv_out_header_9,
  output [15:0] io_pipe_phv_out_header_10,
  output [15:0] io_pipe_phv_out_header_11,
  output [15:0] io_pipe_phv_out_header_12,
  output [15:0] io_pipe_phv_out_header_13,
  output [15:0] io_pipe_phv_out_header_14,
  output [15:0] io_pipe_phv_out_header_15,
  output [7:0]  io_pipe_phv_out_parse_current_state,
  output [7:0]  io_pipe_phv_out_parse_current_offset,
  output [15:0] io_pipe_phv_out_parse_transition_field,
  output [3:0]  io_pipe_phv_out_next_processor_id,
  output        io_pipe_phv_out_next_config_id,
  input  [7:0]  io_offset_in_0,
  input  [7:0]  io_offset_in_1,
  input  [7:0]  io_offset_in_2,
  input  [7:0]  io_offset_in_3,
  input  [7:0]  io_length_in_0,
  input  [7:0]  io_length_in_1,
  input  [7:0]  io_length_in_2,
  input  [7:0]  io_length_in_3,
  input  [63:0] io_field_in_0,
  input  [63:0] io_field_in_1,
  input  [63:0] io_field_in_2,
  input  [63:0] io_field_in_3
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [63:0] _RAND_190;
  reg [63:0] _RAND_191;
  reg [63:0] _RAND_192;
  reg [63:0] _RAND_193;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] phv_data_0; // @[executor.scala 284:22]
  reg [7:0] phv_data_1; // @[executor.scala 284:22]
  reg [7:0] phv_data_2; // @[executor.scala 284:22]
  reg [7:0] phv_data_3; // @[executor.scala 284:22]
  reg [7:0] phv_data_4; // @[executor.scala 284:22]
  reg [7:0] phv_data_5; // @[executor.scala 284:22]
  reg [7:0] phv_data_6; // @[executor.scala 284:22]
  reg [7:0] phv_data_7; // @[executor.scala 284:22]
  reg [7:0] phv_data_8; // @[executor.scala 284:22]
  reg [7:0] phv_data_9; // @[executor.scala 284:22]
  reg [7:0] phv_data_10; // @[executor.scala 284:22]
  reg [7:0] phv_data_11; // @[executor.scala 284:22]
  reg [7:0] phv_data_12; // @[executor.scala 284:22]
  reg [7:0] phv_data_13; // @[executor.scala 284:22]
  reg [7:0] phv_data_14; // @[executor.scala 284:22]
  reg [7:0] phv_data_15; // @[executor.scala 284:22]
  reg [7:0] phv_data_16; // @[executor.scala 284:22]
  reg [7:0] phv_data_17; // @[executor.scala 284:22]
  reg [7:0] phv_data_18; // @[executor.scala 284:22]
  reg [7:0] phv_data_19; // @[executor.scala 284:22]
  reg [7:0] phv_data_20; // @[executor.scala 284:22]
  reg [7:0] phv_data_21; // @[executor.scala 284:22]
  reg [7:0] phv_data_22; // @[executor.scala 284:22]
  reg [7:0] phv_data_23; // @[executor.scala 284:22]
  reg [7:0] phv_data_24; // @[executor.scala 284:22]
  reg [7:0] phv_data_25; // @[executor.scala 284:22]
  reg [7:0] phv_data_26; // @[executor.scala 284:22]
  reg [7:0] phv_data_27; // @[executor.scala 284:22]
  reg [7:0] phv_data_28; // @[executor.scala 284:22]
  reg [7:0] phv_data_29; // @[executor.scala 284:22]
  reg [7:0] phv_data_30; // @[executor.scala 284:22]
  reg [7:0] phv_data_31; // @[executor.scala 284:22]
  reg [7:0] phv_data_32; // @[executor.scala 284:22]
  reg [7:0] phv_data_33; // @[executor.scala 284:22]
  reg [7:0] phv_data_34; // @[executor.scala 284:22]
  reg [7:0] phv_data_35; // @[executor.scala 284:22]
  reg [7:0] phv_data_36; // @[executor.scala 284:22]
  reg [7:0] phv_data_37; // @[executor.scala 284:22]
  reg [7:0] phv_data_38; // @[executor.scala 284:22]
  reg [7:0] phv_data_39; // @[executor.scala 284:22]
  reg [7:0] phv_data_40; // @[executor.scala 284:22]
  reg [7:0] phv_data_41; // @[executor.scala 284:22]
  reg [7:0] phv_data_42; // @[executor.scala 284:22]
  reg [7:0] phv_data_43; // @[executor.scala 284:22]
  reg [7:0] phv_data_44; // @[executor.scala 284:22]
  reg [7:0] phv_data_45; // @[executor.scala 284:22]
  reg [7:0] phv_data_46; // @[executor.scala 284:22]
  reg [7:0] phv_data_47; // @[executor.scala 284:22]
  reg [7:0] phv_data_48; // @[executor.scala 284:22]
  reg [7:0] phv_data_49; // @[executor.scala 284:22]
  reg [7:0] phv_data_50; // @[executor.scala 284:22]
  reg [7:0] phv_data_51; // @[executor.scala 284:22]
  reg [7:0] phv_data_52; // @[executor.scala 284:22]
  reg [7:0] phv_data_53; // @[executor.scala 284:22]
  reg [7:0] phv_data_54; // @[executor.scala 284:22]
  reg [7:0] phv_data_55; // @[executor.scala 284:22]
  reg [7:0] phv_data_56; // @[executor.scala 284:22]
  reg [7:0] phv_data_57; // @[executor.scala 284:22]
  reg [7:0] phv_data_58; // @[executor.scala 284:22]
  reg [7:0] phv_data_59; // @[executor.scala 284:22]
  reg [7:0] phv_data_60; // @[executor.scala 284:22]
  reg [7:0] phv_data_61; // @[executor.scala 284:22]
  reg [7:0] phv_data_62; // @[executor.scala 284:22]
  reg [7:0] phv_data_63; // @[executor.scala 284:22]
  reg [7:0] phv_data_64; // @[executor.scala 284:22]
  reg [7:0] phv_data_65; // @[executor.scala 284:22]
  reg [7:0] phv_data_66; // @[executor.scala 284:22]
  reg [7:0] phv_data_67; // @[executor.scala 284:22]
  reg [7:0] phv_data_68; // @[executor.scala 284:22]
  reg [7:0] phv_data_69; // @[executor.scala 284:22]
  reg [7:0] phv_data_70; // @[executor.scala 284:22]
  reg [7:0] phv_data_71; // @[executor.scala 284:22]
  reg [7:0] phv_data_72; // @[executor.scala 284:22]
  reg [7:0] phv_data_73; // @[executor.scala 284:22]
  reg [7:0] phv_data_74; // @[executor.scala 284:22]
  reg [7:0] phv_data_75; // @[executor.scala 284:22]
  reg [7:0] phv_data_76; // @[executor.scala 284:22]
  reg [7:0] phv_data_77; // @[executor.scala 284:22]
  reg [7:0] phv_data_78; // @[executor.scala 284:22]
  reg [7:0] phv_data_79; // @[executor.scala 284:22]
  reg [7:0] phv_data_80; // @[executor.scala 284:22]
  reg [7:0] phv_data_81; // @[executor.scala 284:22]
  reg [7:0] phv_data_82; // @[executor.scala 284:22]
  reg [7:0] phv_data_83; // @[executor.scala 284:22]
  reg [7:0] phv_data_84; // @[executor.scala 284:22]
  reg [7:0] phv_data_85; // @[executor.scala 284:22]
  reg [7:0] phv_data_86; // @[executor.scala 284:22]
  reg [7:0] phv_data_87; // @[executor.scala 284:22]
  reg [7:0] phv_data_88; // @[executor.scala 284:22]
  reg [7:0] phv_data_89; // @[executor.scala 284:22]
  reg [7:0] phv_data_90; // @[executor.scala 284:22]
  reg [7:0] phv_data_91; // @[executor.scala 284:22]
  reg [7:0] phv_data_92; // @[executor.scala 284:22]
  reg [7:0] phv_data_93; // @[executor.scala 284:22]
  reg [7:0] phv_data_94; // @[executor.scala 284:22]
  reg [7:0] phv_data_95; // @[executor.scala 284:22]
  reg [7:0] phv_data_96; // @[executor.scala 284:22]
  reg [7:0] phv_data_97; // @[executor.scala 284:22]
  reg [7:0] phv_data_98; // @[executor.scala 284:22]
  reg [7:0] phv_data_99; // @[executor.scala 284:22]
  reg [7:0] phv_data_100; // @[executor.scala 284:22]
  reg [7:0] phv_data_101; // @[executor.scala 284:22]
  reg [7:0] phv_data_102; // @[executor.scala 284:22]
  reg [7:0] phv_data_103; // @[executor.scala 284:22]
  reg [7:0] phv_data_104; // @[executor.scala 284:22]
  reg [7:0] phv_data_105; // @[executor.scala 284:22]
  reg [7:0] phv_data_106; // @[executor.scala 284:22]
  reg [7:0] phv_data_107; // @[executor.scala 284:22]
  reg [7:0] phv_data_108; // @[executor.scala 284:22]
  reg [7:0] phv_data_109; // @[executor.scala 284:22]
  reg [7:0] phv_data_110; // @[executor.scala 284:22]
  reg [7:0] phv_data_111; // @[executor.scala 284:22]
  reg [7:0] phv_data_112; // @[executor.scala 284:22]
  reg [7:0] phv_data_113; // @[executor.scala 284:22]
  reg [7:0] phv_data_114; // @[executor.scala 284:22]
  reg [7:0] phv_data_115; // @[executor.scala 284:22]
  reg [7:0] phv_data_116; // @[executor.scala 284:22]
  reg [7:0] phv_data_117; // @[executor.scala 284:22]
  reg [7:0] phv_data_118; // @[executor.scala 284:22]
  reg [7:0] phv_data_119; // @[executor.scala 284:22]
  reg [7:0] phv_data_120; // @[executor.scala 284:22]
  reg [7:0] phv_data_121; // @[executor.scala 284:22]
  reg [7:0] phv_data_122; // @[executor.scala 284:22]
  reg [7:0] phv_data_123; // @[executor.scala 284:22]
  reg [7:0] phv_data_124; // @[executor.scala 284:22]
  reg [7:0] phv_data_125; // @[executor.scala 284:22]
  reg [7:0] phv_data_126; // @[executor.scala 284:22]
  reg [7:0] phv_data_127; // @[executor.scala 284:22]
  reg [7:0] phv_data_128; // @[executor.scala 284:22]
  reg [7:0] phv_data_129; // @[executor.scala 284:22]
  reg [7:0] phv_data_130; // @[executor.scala 284:22]
  reg [7:0] phv_data_131; // @[executor.scala 284:22]
  reg [7:0] phv_data_132; // @[executor.scala 284:22]
  reg [7:0] phv_data_133; // @[executor.scala 284:22]
  reg [7:0] phv_data_134; // @[executor.scala 284:22]
  reg [7:0] phv_data_135; // @[executor.scala 284:22]
  reg [7:0] phv_data_136; // @[executor.scala 284:22]
  reg [7:0] phv_data_137; // @[executor.scala 284:22]
  reg [7:0] phv_data_138; // @[executor.scala 284:22]
  reg [7:0] phv_data_139; // @[executor.scala 284:22]
  reg [7:0] phv_data_140; // @[executor.scala 284:22]
  reg [7:0] phv_data_141; // @[executor.scala 284:22]
  reg [7:0] phv_data_142; // @[executor.scala 284:22]
  reg [7:0] phv_data_143; // @[executor.scala 284:22]
  reg [7:0] phv_data_144; // @[executor.scala 284:22]
  reg [7:0] phv_data_145; // @[executor.scala 284:22]
  reg [7:0] phv_data_146; // @[executor.scala 284:22]
  reg [7:0] phv_data_147; // @[executor.scala 284:22]
  reg [7:0] phv_data_148; // @[executor.scala 284:22]
  reg [7:0] phv_data_149; // @[executor.scala 284:22]
  reg [7:0] phv_data_150; // @[executor.scala 284:22]
  reg [7:0] phv_data_151; // @[executor.scala 284:22]
  reg [7:0] phv_data_152; // @[executor.scala 284:22]
  reg [7:0] phv_data_153; // @[executor.scala 284:22]
  reg [7:0] phv_data_154; // @[executor.scala 284:22]
  reg [7:0] phv_data_155; // @[executor.scala 284:22]
  reg [7:0] phv_data_156; // @[executor.scala 284:22]
  reg [7:0] phv_data_157; // @[executor.scala 284:22]
  reg [7:0] phv_data_158; // @[executor.scala 284:22]
  reg [7:0] phv_data_159; // @[executor.scala 284:22]
  reg [15:0] phv_header_0; // @[executor.scala 284:22]
  reg [15:0] phv_header_1; // @[executor.scala 284:22]
  reg [15:0] phv_header_2; // @[executor.scala 284:22]
  reg [15:0] phv_header_3; // @[executor.scala 284:22]
  reg [15:0] phv_header_4; // @[executor.scala 284:22]
  reg [15:0] phv_header_5; // @[executor.scala 284:22]
  reg [15:0] phv_header_6; // @[executor.scala 284:22]
  reg [15:0] phv_header_7; // @[executor.scala 284:22]
  reg [15:0] phv_header_8; // @[executor.scala 284:22]
  reg [15:0] phv_header_9; // @[executor.scala 284:22]
  reg [15:0] phv_header_10; // @[executor.scala 284:22]
  reg [15:0] phv_header_11; // @[executor.scala 284:22]
  reg [15:0] phv_header_12; // @[executor.scala 284:22]
  reg [15:0] phv_header_13; // @[executor.scala 284:22]
  reg [15:0] phv_header_14; // @[executor.scala 284:22]
  reg [15:0] phv_header_15; // @[executor.scala 284:22]
  reg [7:0] phv_parse_current_state; // @[executor.scala 284:22]
  reg [7:0] phv_parse_current_offset; // @[executor.scala 284:22]
  reg [15:0] phv_parse_transition_field; // @[executor.scala 284:22]
  reg [3:0] phv_next_processor_id; // @[executor.scala 284:22]
  reg  phv_next_config_id; // @[executor.scala 284:22]
  reg  phv_is_valid_processor; // @[executor.scala 284:22]
  reg [7:0] offset_0; // @[executor.scala 288:25]
  reg [7:0] offset_1; // @[executor.scala 288:25]
  reg [7:0] offset_2; // @[executor.scala 288:25]
  reg [7:0] offset_3; // @[executor.scala 288:25]
  reg [7:0] length_0; // @[executor.scala 289:25]
  reg [7:0] length_1; // @[executor.scala 289:25]
  reg [7:0] length_2; // @[executor.scala 289:25]
  reg [7:0] length_3; // @[executor.scala 289:25]
  reg [63:0] field_0; // @[executor.scala 290:25]
  reg [63:0] field_1; // @[executor.scala 290:25]
  reg [63:0] field_2; // @[executor.scala 290:25]
  reg [63:0] field_3; // @[executor.scala 290:25]
  wire [7:0] field_byte = field_0[63:56]; // @[executor.scala 305:57]
  wire [8:0] _total_offset_T = {{1'd0}, offset_0}; // @[executor.scala 307:57]
  wire [7:0] total_offset = _total_offset_T[7:0]; // @[executor.scala 307:57]
  wire [7:0] _GEN_0 = 8'h0 == total_offset ? field_byte : phv_data_0; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_1 = 8'h1 == total_offset ? field_byte : phv_data_1; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_2 = 8'h2 == total_offset ? field_byte : phv_data_2; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_3 = 8'h3 == total_offset ? field_byte : phv_data_3; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_4 = 8'h4 == total_offset ? field_byte : phv_data_4; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_5 = 8'h5 == total_offset ? field_byte : phv_data_5; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_6 = 8'h6 == total_offset ? field_byte : phv_data_6; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_7 = 8'h7 == total_offset ? field_byte : phv_data_7; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_8 = 8'h8 == total_offset ? field_byte : phv_data_8; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_9 = 8'h9 == total_offset ? field_byte : phv_data_9; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_10 = 8'ha == total_offset ? field_byte : phv_data_10; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_11 = 8'hb == total_offset ? field_byte : phv_data_11; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_12 = 8'hc == total_offset ? field_byte : phv_data_12; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_13 = 8'hd == total_offset ? field_byte : phv_data_13; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_14 = 8'he == total_offset ? field_byte : phv_data_14; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_15 = 8'hf == total_offset ? field_byte : phv_data_15; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_16 = 8'h10 == total_offset ? field_byte : phv_data_16; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_17 = 8'h11 == total_offset ? field_byte : phv_data_17; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_18 = 8'h12 == total_offset ? field_byte : phv_data_18; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_19 = 8'h13 == total_offset ? field_byte : phv_data_19; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_20 = 8'h14 == total_offset ? field_byte : phv_data_20; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_21 = 8'h15 == total_offset ? field_byte : phv_data_21; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_22 = 8'h16 == total_offset ? field_byte : phv_data_22; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_23 = 8'h17 == total_offset ? field_byte : phv_data_23; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_24 = 8'h18 == total_offset ? field_byte : phv_data_24; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_25 = 8'h19 == total_offset ? field_byte : phv_data_25; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_26 = 8'h1a == total_offset ? field_byte : phv_data_26; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_27 = 8'h1b == total_offset ? field_byte : phv_data_27; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_28 = 8'h1c == total_offset ? field_byte : phv_data_28; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_29 = 8'h1d == total_offset ? field_byte : phv_data_29; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_30 = 8'h1e == total_offset ? field_byte : phv_data_30; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_31 = 8'h1f == total_offset ? field_byte : phv_data_31; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_32 = 8'h20 == total_offset ? field_byte : phv_data_32; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_33 = 8'h21 == total_offset ? field_byte : phv_data_33; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_34 = 8'h22 == total_offset ? field_byte : phv_data_34; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_35 = 8'h23 == total_offset ? field_byte : phv_data_35; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_36 = 8'h24 == total_offset ? field_byte : phv_data_36; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_37 = 8'h25 == total_offset ? field_byte : phv_data_37; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_38 = 8'h26 == total_offset ? field_byte : phv_data_38; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_39 = 8'h27 == total_offset ? field_byte : phv_data_39; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_40 = 8'h28 == total_offset ? field_byte : phv_data_40; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_41 = 8'h29 == total_offset ? field_byte : phv_data_41; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_42 = 8'h2a == total_offset ? field_byte : phv_data_42; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_43 = 8'h2b == total_offset ? field_byte : phv_data_43; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_44 = 8'h2c == total_offset ? field_byte : phv_data_44; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_45 = 8'h2d == total_offset ? field_byte : phv_data_45; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_46 = 8'h2e == total_offset ? field_byte : phv_data_46; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_47 = 8'h2f == total_offset ? field_byte : phv_data_47; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_48 = 8'h30 == total_offset ? field_byte : phv_data_48; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_49 = 8'h31 == total_offset ? field_byte : phv_data_49; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_50 = 8'h32 == total_offset ? field_byte : phv_data_50; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_51 = 8'h33 == total_offset ? field_byte : phv_data_51; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_52 = 8'h34 == total_offset ? field_byte : phv_data_52; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_53 = 8'h35 == total_offset ? field_byte : phv_data_53; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_54 = 8'h36 == total_offset ? field_byte : phv_data_54; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_55 = 8'h37 == total_offset ? field_byte : phv_data_55; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_56 = 8'h38 == total_offset ? field_byte : phv_data_56; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_57 = 8'h39 == total_offset ? field_byte : phv_data_57; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_58 = 8'h3a == total_offset ? field_byte : phv_data_58; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_59 = 8'h3b == total_offset ? field_byte : phv_data_59; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_60 = 8'h3c == total_offset ? field_byte : phv_data_60; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_61 = 8'h3d == total_offset ? field_byte : phv_data_61; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_62 = 8'h3e == total_offset ? field_byte : phv_data_62; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_63 = 8'h3f == total_offset ? field_byte : phv_data_63; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_64 = 8'h40 == total_offset ? field_byte : phv_data_64; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_65 = 8'h41 == total_offset ? field_byte : phv_data_65; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_66 = 8'h42 == total_offset ? field_byte : phv_data_66; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_67 = 8'h43 == total_offset ? field_byte : phv_data_67; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_68 = 8'h44 == total_offset ? field_byte : phv_data_68; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_69 = 8'h45 == total_offset ? field_byte : phv_data_69; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_70 = 8'h46 == total_offset ? field_byte : phv_data_70; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_71 = 8'h47 == total_offset ? field_byte : phv_data_71; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_72 = 8'h48 == total_offset ? field_byte : phv_data_72; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_73 = 8'h49 == total_offset ? field_byte : phv_data_73; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_74 = 8'h4a == total_offset ? field_byte : phv_data_74; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_75 = 8'h4b == total_offset ? field_byte : phv_data_75; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_76 = 8'h4c == total_offset ? field_byte : phv_data_76; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_77 = 8'h4d == total_offset ? field_byte : phv_data_77; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_78 = 8'h4e == total_offset ? field_byte : phv_data_78; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_79 = 8'h4f == total_offset ? field_byte : phv_data_79; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_80 = 8'h50 == total_offset ? field_byte : phv_data_80; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_81 = 8'h51 == total_offset ? field_byte : phv_data_81; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_82 = 8'h52 == total_offset ? field_byte : phv_data_82; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_83 = 8'h53 == total_offset ? field_byte : phv_data_83; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_84 = 8'h54 == total_offset ? field_byte : phv_data_84; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_85 = 8'h55 == total_offset ? field_byte : phv_data_85; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_86 = 8'h56 == total_offset ? field_byte : phv_data_86; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_87 = 8'h57 == total_offset ? field_byte : phv_data_87; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_88 = 8'h58 == total_offset ? field_byte : phv_data_88; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_89 = 8'h59 == total_offset ? field_byte : phv_data_89; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_90 = 8'h5a == total_offset ? field_byte : phv_data_90; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_91 = 8'h5b == total_offset ? field_byte : phv_data_91; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_92 = 8'h5c == total_offset ? field_byte : phv_data_92; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_93 = 8'h5d == total_offset ? field_byte : phv_data_93; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_94 = 8'h5e == total_offset ? field_byte : phv_data_94; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_95 = 8'h5f == total_offset ? field_byte : phv_data_95; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_96 = 8'h60 == total_offset ? field_byte : phv_data_96; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_97 = 8'h61 == total_offset ? field_byte : phv_data_97; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_98 = 8'h62 == total_offset ? field_byte : phv_data_98; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_99 = 8'h63 == total_offset ? field_byte : phv_data_99; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_100 = 8'h64 == total_offset ? field_byte : phv_data_100; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_101 = 8'h65 == total_offset ? field_byte : phv_data_101; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_102 = 8'h66 == total_offset ? field_byte : phv_data_102; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_103 = 8'h67 == total_offset ? field_byte : phv_data_103; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_104 = 8'h68 == total_offset ? field_byte : phv_data_104; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_105 = 8'h69 == total_offset ? field_byte : phv_data_105; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_106 = 8'h6a == total_offset ? field_byte : phv_data_106; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_107 = 8'h6b == total_offset ? field_byte : phv_data_107; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_108 = 8'h6c == total_offset ? field_byte : phv_data_108; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_109 = 8'h6d == total_offset ? field_byte : phv_data_109; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_110 = 8'h6e == total_offset ? field_byte : phv_data_110; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_111 = 8'h6f == total_offset ? field_byte : phv_data_111; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_112 = 8'h70 == total_offset ? field_byte : phv_data_112; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_113 = 8'h71 == total_offset ? field_byte : phv_data_113; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_114 = 8'h72 == total_offset ? field_byte : phv_data_114; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_115 = 8'h73 == total_offset ? field_byte : phv_data_115; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_116 = 8'h74 == total_offset ? field_byte : phv_data_116; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_117 = 8'h75 == total_offset ? field_byte : phv_data_117; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_118 = 8'h76 == total_offset ? field_byte : phv_data_118; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_119 = 8'h77 == total_offset ? field_byte : phv_data_119; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_120 = 8'h78 == total_offset ? field_byte : phv_data_120; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_121 = 8'h79 == total_offset ? field_byte : phv_data_121; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_122 = 8'h7a == total_offset ? field_byte : phv_data_122; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_123 = 8'h7b == total_offset ? field_byte : phv_data_123; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_124 = 8'h7c == total_offset ? field_byte : phv_data_124; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_125 = 8'h7d == total_offset ? field_byte : phv_data_125; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_126 = 8'h7e == total_offset ? field_byte : phv_data_126; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_127 = 8'h7f == total_offset ? field_byte : phv_data_127; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_128 = 8'h80 == total_offset ? field_byte : phv_data_128; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_129 = 8'h81 == total_offset ? field_byte : phv_data_129; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_130 = 8'h82 == total_offset ? field_byte : phv_data_130; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_131 = 8'h83 == total_offset ? field_byte : phv_data_131; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_132 = 8'h84 == total_offset ? field_byte : phv_data_132; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_133 = 8'h85 == total_offset ? field_byte : phv_data_133; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_134 = 8'h86 == total_offset ? field_byte : phv_data_134; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_135 = 8'h87 == total_offset ? field_byte : phv_data_135; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_136 = 8'h88 == total_offset ? field_byte : phv_data_136; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_137 = 8'h89 == total_offset ? field_byte : phv_data_137; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_138 = 8'h8a == total_offset ? field_byte : phv_data_138; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_139 = 8'h8b == total_offset ? field_byte : phv_data_139; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_140 = 8'h8c == total_offset ? field_byte : phv_data_140; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_141 = 8'h8d == total_offset ? field_byte : phv_data_141; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_142 = 8'h8e == total_offset ? field_byte : phv_data_142; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_143 = 8'h8f == total_offset ? field_byte : phv_data_143; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_144 = 8'h90 == total_offset ? field_byte : phv_data_144; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_145 = 8'h91 == total_offset ? field_byte : phv_data_145; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_146 = 8'h92 == total_offset ? field_byte : phv_data_146; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_147 = 8'h93 == total_offset ? field_byte : phv_data_147; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_148 = 8'h94 == total_offset ? field_byte : phv_data_148; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_149 = 8'h95 == total_offset ? field_byte : phv_data_149; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_150 = 8'h96 == total_offset ? field_byte : phv_data_150; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_151 = 8'h97 == total_offset ? field_byte : phv_data_151; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_152 = 8'h98 == total_offset ? field_byte : phv_data_152; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_153 = 8'h99 == total_offset ? field_byte : phv_data_153; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_154 = 8'h9a == total_offset ? field_byte : phv_data_154; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_155 = 8'h9b == total_offset ? field_byte : phv_data_155; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_156 = 8'h9c == total_offset ? field_byte : phv_data_156; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_157 = 8'h9d == total_offset ? field_byte : phv_data_157; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_158 = 8'h9e == total_offset ? field_byte : phv_data_158; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_159 = 8'h9f == total_offset ? field_byte : phv_data_159; // @[executor.scala 309:64 executor.scala 309:64 executor.scala 286:25]
  wire [7:0] _GEN_160 = 8'h0 < length_0 ? _GEN_0 : phv_data_0; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_161 = 8'h0 < length_0 ? _GEN_1 : phv_data_1; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_162 = 8'h0 < length_0 ? _GEN_2 : phv_data_2; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_163 = 8'h0 < length_0 ? _GEN_3 : phv_data_3; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_164 = 8'h0 < length_0 ? _GEN_4 : phv_data_4; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_165 = 8'h0 < length_0 ? _GEN_5 : phv_data_5; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_166 = 8'h0 < length_0 ? _GEN_6 : phv_data_6; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_167 = 8'h0 < length_0 ? _GEN_7 : phv_data_7; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_168 = 8'h0 < length_0 ? _GEN_8 : phv_data_8; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_169 = 8'h0 < length_0 ? _GEN_9 : phv_data_9; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_170 = 8'h0 < length_0 ? _GEN_10 : phv_data_10; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_171 = 8'h0 < length_0 ? _GEN_11 : phv_data_11; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_172 = 8'h0 < length_0 ? _GEN_12 : phv_data_12; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_173 = 8'h0 < length_0 ? _GEN_13 : phv_data_13; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_174 = 8'h0 < length_0 ? _GEN_14 : phv_data_14; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_175 = 8'h0 < length_0 ? _GEN_15 : phv_data_15; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_176 = 8'h0 < length_0 ? _GEN_16 : phv_data_16; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_177 = 8'h0 < length_0 ? _GEN_17 : phv_data_17; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_178 = 8'h0 < length_0 ? _GEN_18 : phv_data_18; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_179 = 8'h0 < length_0 ? _GEN_19 : phv_data_19; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_180 = 8'h0 < length_0 ? _GEN_20 : phv_data_20; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_181 = 8'h0 < length_0 ? _GEN_21 : phv_data_21; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_182 = 8'h0 < length_0 ? _GEN_22 : phv_data_22; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_183 = 8'h0 < length_0 ? _GEN_23 : phv_data_23; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_184 = 8'h0 < length_0 ? _GEN_24 : phv_data_24; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_185 = 8'h0 < length_0 ? _GEN_25 : phv_data_25; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_186 = 8'h0 < length_0 ? _GEN_26 : phv_data_26; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_187 = 8'h0 < length_0 ? _GEN_27 : phv_data_27; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_188 = 8'h0 < length_0 ? _GEN_28 : phv_data_28; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_189 = 8'h0 < length_0 ? _GEN_29 : phv_data_29; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_190 = 8'h0 < length_0 ? _GEN_30 : phv_data_30; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_191 = 8'h0 < length_0 ? _GEN_31 : phv_data_31; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_192 = 8'h0 < length_0 ? _GEN_32 : phv_data_32; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_193 = 8'h0 < length_0 ? _GEN_33 : phv_data_33; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_194 = 8'h0 < length_0 ? _GEN_34 : phv_data_34; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_195 = 8'h0 < length_0 ? _GEN_35 : phv_data_35; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_196 = 8'h0 < length_0 ? _GEN_36 : phv_data_36; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_197 = 8'h0 < length_0 ? _GEN_37 : phv_data_37; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_198 = 8'h0 < length_0 ? _GEN_38 : phv_data_38; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_199 = 8'h0 < length_0 ? _GEN_39 : phv_data_39; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_200 = 8'h0 < length_0 ? _GEN_40 : phv_data_40; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_201 = 8'h0 < length_0 ? _GEN_41 : phv_data_41; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_202 = 8'h0 < length_0 ? _GEN_42 : phv_data_42; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_203 = 8'h0 < length_0 ? _GEN_43 : phv_data_43; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_204 = 8'h0 < length_0 ? _GEN_44 : phv_data_44; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_205 = 8'h0 < length_0 ? _GEN_45 : phv_data_45; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_206 = 8'h0 < length_0 ? _GEN_46 : phv_data_46; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_207 = 8'h0 < length_0 ? _GEN_47 : phv_data_47; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_208 = 8'h0 < length_0 ? _GEN_48 : phv_data_48; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_209 = 8'h0 < length_0 ? _GEN_49 : phv_data_49; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_210 = 8'h0 < length_0 ? _GEN_50 : phv_data_50; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_211 = 8'h0 < length_0 ? _GEN_51 : phv_data_51; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_212 = 8'h0 < length_0 ? _GEN_52 : phv_data_52; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_213 = 8'h0 < length_0 ? _GEN_53 : phv_data_53; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_214 = 8'h0 < length_0 ? _GEN_54 : phv_data_54; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_215 = 8'h0 < length_0 ? _GEN_55 : phv_data_55; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_216 = 8'h0 < length_0 ? _GEN_56 : phv_data_56; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_217 = 8'h0 < length_0 ? _GEN_57 : phv_data_57; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_218 = 8'h0 < length_0 ? _GEN_58 : phv_data_58; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_219 = 8'h0 < length_0 ? _GEN_59 : phv_data_59; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_220 = 8'h0 < length_0 ? _GEN_60 : phv_data_60; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_221 = 8'h0 < length_0 ? _GEN_61 : phv_data_61; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_222 = 8'h0 < length_0 ? _GEN_62 : phv_data_62; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_223 = 8'h0 < length_0 ? _GEN_63 : phv_data_63; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_224 = 8'h0 < length_0 ? _GEN_64 : phv_data_64; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_225 = 8'h0 < length_0 ? _GEN_65 : phv_data_65; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_226 = 8'h0 < length_0 ? _GEN_66 : phv_data_66; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_227 = 8'h0 < length_0 ? _GEN_67 : phv_data_67; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_228 = 8'h0 < length_0 ? _GEN_68 : phv_data_68; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_229 = 8'h0 < length_0 ? _GEN_69 : phv_data_69; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_230 = 8'h0 < length_0 ? _GEN_70 : phv_data_70; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_231 = 8'h0 < length_0 ? _GEN_71 : phv_data_71; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_232 = 8'h0 < length_0 ? _GEN_72 : phv_data_72; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_233 = 8'h0 < length_0 ? _GEN_73 : phv_data_73; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_234 = 8'h0 < length_0 ? _GEN_74 : phv_data_74; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_235 = 8'h0 < length_0 ? _GEN_75 : phv_data_75; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_236 = 8'h0 < length_0 ? _GEN_76 : phv_data_76; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_237 = 8'h0 < length_0 ? _GEN_77 : phv_data_77; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_238 = 8'h0 < length_0 ? _GEN_78 : phv_data_78; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_239 = 8'h0 < length_0 ? _GEN_79 : phv_data_79; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_240 = 8'h0 < length_0 ? _GEN_80 : phv_data_80; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_241 = 8'h0 < length_0 ? _GEN_81 : phv_data_81; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_242 = 8'h0 < length_0 ? _GEN_82 : phv_data_82; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_243 = 8'h0 < length_0 ? _GEN_83 : phv_data_83; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_244 = 8'h0 < length_0 ? _GEN_84 : phv_data_84; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_245 = 8'h0 < length_0 ? _GEN_85 : phv_data_85; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_246 = 8'h0 < length_0 ? _GEN_86 : phv_data_86; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_247 = 8'h0 < length_0 ? _GEN_87 : phv_data_87; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_248 = 8'h0 < length_0 ? _GEN_88 : phv_data_88; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_249 = 8'h0 < length_0 ? _GEN_89 : phv_data_89; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_250 = 8'h0 < length_0 ? _GEN_90 : phv_data_90; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_251 = 8'h0 < length_0 ? _GEN_91 : phv_data_91; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_252 = 8'h0 < length_0 ? _GEN_92 : phv_data_92; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_253 = 8'h0 < length_0 ? _GEN_93 : phv_data_93; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_254 = 8'h0 < length_0 ? _GEN_94 : phv_data_94; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_255 = 8'h0 < length_0 ? _GEN_95 : phv_data_95; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_256 = 8'h0 < length_0 ? _GEN_96 : phv_data_96; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_257 = 8'h0 < length_0 ? _GEN_97 : phv_data_97; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_258 = 8'h0 < length_0 ? _GEN_98 : phv_data_98; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_259 = 8'h0 < length_0 ? _GEN_99 : phv_data_99; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_260 = 8'h0 < length_0 ? _GEN_100 : phv_data_100; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_261 = 8'h0 < length_0 ? _GEN_101 : phv_data_101; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_262 = 8'h0 < length_0 ? _GEN_102 : phv_data_102; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_263 = 8'h0 < length_0 ? _GEN_103 : phv_data_103; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_264 = 8'h0 < length_0 ? _GEN_104 : phv_data_104; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_265 = 8'h0 < length_0 ? _GEN_105 : phv_data_105; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_266 = 8'h0 < length_0 ? _GEN_106 : phv_data_106; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_267 = 8'h0 < length_0 ? _GEN_107 : phv_data_107; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_268 = 8'h0 < length_0 ? _GEN_108 : phv_data_108; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_269 = 8'h0 < length_0 ? _GEN_109 : phv_data_109; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_270 = 8'h0 < length_0 ? _GEN_110 : phv_data_110; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_271 = 8'h0 < length_0 ? _GEN_111 : phv_data_111; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_272 = 8'h0 < length_0 ? _GEN_112 : phv_data_112; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_273 = 8'h0 < length_0 ? _GEN_113 : phv_data_113; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_274 = 8'h0 < length_0 ? _GEN_114 : phv_data_114; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_275 = 8'h0 < length_0 ? _GEN_115 : phv_data_115; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_276 = 8'h0 < length_0 ? _GEN_116 : phv_data_116; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_277 = 8'h0 < length_0 ? _GEN_117 : phv_data_117; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_278 = 8'h0 < length_0 ? _GEN_118 : phv_data_118; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_279 = 8'h0 < length_0 ? _GEN_119 : phv_data_119; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_280 = 8'h0 < length_0 ? _GEN_120 : phv_data_120; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_281 = 8'h0 < length_0 ? _GEN_121 : phv_data_121; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_282 = 8'h0 < length_0 ? _GEN_122 : phv_data_122; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_283 = 8'h0 < length_0 ? _GEN_123 : phv_data_123; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_284 = 8'h0 < length_0 ? _GEN_124 : phv_data_124; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_285 = 8'h0 < length_0 ? _GEN_125 : phv_data_125; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_286 = 8'h0 < length_0 ? _GEN_126 : phv_data_126; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_287 = 8'h0 < length_0 ? _GEN_127 : phv_data_127; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_288 = 8'h0 < length_0 ? _GEN_128 : phv_data_128; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_289 = 8'h0 < length_0 ? _GEN_129 : phv_data_129; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_290 = 8'h0 < length_0 ? _GEN_130 : phv_data_130; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_291 = 8'h0 < length_0 ? _GEN_131 : phv_data_131; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_292 = 8'h0 < length_0 ? _GEN_132 : phv_data_132; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_293 = 8'h0 < length_0 ? _GEN_133 : phv_data_133; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_294 = 8'h0 < length_0 ? _GEN_134 : phv_data_134; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_295 = 8'h0 < length_0 ? _GEN_135 : phv_data_135; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_296 = 8'h0 < length_0 ? _GEN_136 : phv_data_136; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_297 = 8'h0 < length_0 ? _GEN_137 : phv_data_137; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_298 = 8'h0 < length_0 ? _GEN_138 : phv_data_138; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_299 = 8'h0 < length_0 ? _GEN_139 : phv_data_139; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_300 = 8'h0 < length_0 ? _GEN_140 : phv_data_140; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_301 = 8'h0 < length_0 ? _GEN_141 : phv_data_141; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_302 = 8'h0 < length_0 ? _GEN_142 : phv_data_142; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_303 = 8'h0 < length_0 ? _GEN_143 : phv_data_143; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_304 = 8'h0 < length_0 ? _GEN_144 : phv_data_144; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_305 = 8'h0 < length_0 ? _GEN_145 : phv_data_145; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_306 = 8'h0 < length_0 ? _GEN_146 : phv_data_146; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_307 = 8'h0 < length_0 ? _GEN_147 : phv_data_147; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_308 = 8'h0 < length_0 ? _GEN_148 : phv_data_148; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_309 = 8'h0 < length_0 ? _GEN_149 : phv_data_149; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_310 = 8'h0 < length_0 ? _GEN_150 : phv_data_150; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_311 = 8'h0 < length_0 ? _GEN_151 : phv_data_151; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_312 = 8'h0 < length_0 ? _GEN_152 : phv_data_152; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_313 = 8'h0 < length_0 ? _GEN_153 : phv_data_153; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_314 = 8'h0 < length_0 ? _GEN_154 : phv_data_154; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_315 = 8'h0 < length_0 ? _GEN_155 : phv_data_155; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_316 = 8'h0 < length_0 ? _GEN_156 : phv_data_156; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_317 = 8'h0 < length_0 ? _GEN_157 : phv_data_157; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_318 = 8'h0 < length_0 ? _GEN_158 : phv_data_158; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] _GEN_319 = 8'h0 < length_0 ? _GEN_159 : phv_data_159; // @[executor.scala 308:60 executor.scala 286:25]
  wire [7:0] field_byte_1 = field_0[55:48]; // @[executor.scala 305:57]
  wire [7:0] total_offset_1 = offset_0 + 8'h1; // @[executor.scala 307:57]
  wire [7:0] _GEN_320 = 8'h0 == total_offset_1 ? field_byte_1 : _GEN_160; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_321 = 8'h1 == total_offset_1 ? field_byte_1 : _GEN_161; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_322 = 8'h2 == total_offset_1 ? field_byte_1 : _GEN_162; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_323 = 8'h3 == total_offset_1 ? field_byte_1 : _GEN_163; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_324 = 8'h4 == total_offset_1 ? field_byte_1 : _GEN_164; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_325 = 8'h5 == total_offset_1 ? field_byte_1 : _GEN_165; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_326 = 8'h6 == total_offset_1 ? field_byte_1 : _GEN_166; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_327 = 8'h7 == total_offset_1 ? field_byte_1 : _GEN_167; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_328 = 8'h8 == total_offset_1 ? field_byte_1 : _GEN_168; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_329 = 8'h9 == total_offset_1 ? field_byte_1 : _GEN_169; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_330 = 8'ha == total_offset_1 ? field_byte_1 : _GEN_170; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_331 = 8'hb == total_offset_1 ? field_byte_1 : _GEN_171; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_332 = 8'hc == total_offset_1 ? field_byte_1 : _GEN_172; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_333 = 8'hd == total_offset_1 ? field_byte_1 : _GEN_173; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_334 = 8'he == total_offset_1 ? field_byte_1 : _GEN_174; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_335 = 8'hf == total_offset_1 ? field_byte_1 : _GEN_175; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_336 = 8'h10 == total_offset_1 ? field_byte_1 : _GEN_176; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_337 = 8'h11 == total_offset_1 ? field_byte_1 : _GEN_177; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_338 = 8'h12 == total_offset_1 ? field_byte_1 : _GEN_178; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_339 = 8'h13 == total_offset_1 ? field_byte_1 : _GEN_179; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_340 = 8'h14 == total_offset_1 ? field_byte_1 : _GEN_180; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_341 = 8'h15 == total_offset_1 ? field_byte_1 : _GEN_181; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_342 = 8'h16 == total_offset_1 ? field_byte_1 : _GEN_182; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_343 = 8'h17 == total_offset_1 ? field_byte_1 : _GEN_183; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_344 = 8'h18 == total_offset_1 ? field_byte_1 : _GEN_184; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_345 = 8'h19 == total_offset_1 ? field_byte_1 : _GEN_185; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_346 = 8'h1a == total_offset_1 ? field_byte_1 : _GEN_186; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_347 = 8'h1b == total_offset_1 ? field_byte_1 : _GEN_187; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_348 = 8'h1c == total_offset_1 ? field_byte_1 : _GEN_188; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_349 = 8'h1d == total_offset_1 ? field_byte_1 : _GEN_189; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_350 = 8'h1e == total_offset_1 ? field_byte_1 : _GEN_190; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_351 = 8'h1f == total_offset_1 ? field_byte_1 : _GEN_191; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_352 = 8'h20 == total_offset_1 ? field_byte_1 : _GEN_192; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_353 = 8'h21 == total_offset_1 ? field_byte_1 : _GEN_193; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_354 = 8'h22 == total_offset_1 ? field_byte_1 : _GEN_194; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_355 = 8'h23 == total_offset_1 ? field_byte_1 : _GEN_195; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_356 = 8'h24 == total_offset_1 ? field_byte_1 : _GEN_196; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_357 = 8'h25 == total_offset_1 ? field_byte_1 : _GEN_197; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_358 = 8'h26 == total_offset_1 ? field_byte_1 : _GEN_198; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_359 = 8'h27 == total_offset_1 ? field_byte_1 : _GEN_199; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_360 = 8'h28 == total_offset_1 ? field_byte_1 : _GEN_200; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_361 = 8'h29 == total_offset_1 ? field_byte_1 : _GEN_201; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_362 = 8'h2a == total_offset_1 ? field_byte_1 : _GEN_202; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_363 = 8'h2b == total_offset_1 ? field_byte_1 : _GEN_203; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_364 = 8'h2c == total_offset_1 ? field_byte_1 : _GEN_204; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_365 = 8'h2d == total_offset_1 ? field_byte_1 : _GEN_205; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_366 = 8'h2e == total_offset_1 ? field_byte_1 : _GEN_206; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_367 = 8'h2f == total_offset_1 ? field_byte_1 : _GEN_207; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_368 = 8'h30 == total_offset_1 ? field_byte_1 : _GEN_208; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_369 = 8'h31 == total_offset_1 ? field_byte_1 : _GEN_209; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_370 = 8'h32 == total_offset_1 ? field_byte_1 : _GEN_210; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_371 = 8'h33 == total_offset_1 ? field_byte_1 : _GEN_211; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_372 = 8'h34 == total_offset_1 ? field_byte_1 : _GEN_212; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_373 = 8'h35 == total_offset_1 ? field_byte_1 : _GEN_213; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_374 = 8'h36 == total_offset_1 ? field_byte_1 : _GEN_214; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_375 = 8'h37 == total_offset_1 ? field_byte_1 : _GEN_215; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_376 = 8'h38 == total_offset_1 ? field_byte_1 : _GEN_216; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_377 = 8'h39 == total_offset_1 ? field_byte_1 : _GEN_217; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_378 = 8'h3a == total_offset_1 ? field_byte_1 : _GEN_218; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_379 = 8'h3b == total_offset_1 ? field_byte_1 : _GEN_219; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_380 = 8'h3c == total_offset_1 ? field_byte_1 : _GEN_220; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_381 = 8'h3d == total_offset_1 ? field_byte_1 : _GEN_221; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_382 = 8'h3e == total_offset_1 ? field_byte_1 : _GEN_222; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_383 = 8'h3f == total_offset_1 ? field_byte_1 : _GEN_223; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_384 = 8'h40 == total_offset_1 ? field_byte_1 : _GEN_224; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_385 = 8'h41 == total_offset_1 ? field_byte_1 : _GEN_225; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_386 = 8'h42 == total_offset_1 ? field_byte_1 : _GEN_226; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_387 = 8'h43 == total_offset_1 ? field_byte_1 : _GEN_227; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_388 = 8'h44 == total_offset_1 ? field_byte_1 : _GEN_228; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_389 = 8'h45 == total_offset_1 ? field_byte_1 : _GEN_229; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_390 = 8'h46 == total_offset_1 ? field_byte_1 : _GEN_230; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_391 = 8'h47 == total_offset_1 ? field_byte_1 : _GEN_231; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_392 = 8'h48 == total_offset_1 ? field_byte_1 : _GEN_232; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_393 = 8'h49 == total_offset_1 ? field_byte_1 : _GEN_233; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_394 = 8'h4a == total_offset_1 ? field_byte_1 : _GEN_234; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_395 = 8'h4b == total_offset_1 ? field_byte_1 : _GEN_235; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_396 = 8'h4c == total_offset_1 ? field_byte_1 : _GEN_236; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_397 = 8'h4d == total_offset_1 ? field_byte_1 : _GEN_237; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_398 = 8'h4e == total_offset_1 ? field_byte_1 : _GEN_238; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_399 = 8'h4f == total_offset_1 ? field_byte_1 : _GEN_239; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_400 = 8'h50 == total_offset_1 ? field_byte_1 : _GEN_240; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_401 = 8'h51 == total_offset_1 ? field_byte_1 : _GEN_241; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_402 = 8'h52 == total_offset_1 ? field_byte_1 : _GEN_242; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_403 = 8'h53 == total_offset_1 ? field_byte_1 : _GEN_243; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_404 = 8'h54 == total_offset_1 ? field_byte_1 : _GEN_244; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_405 = 8'h55 == total_offset_1 ? field_byte_1 : _GEN_245; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_406 = 8'h56 == total_offset_1 ? field_byte_1 : _GEN_246; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_407 = 8'h57 == total_offset_1 ? field_byte_1 : _GEN_247; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_408 = 8'h58 == total_offset_1 ? field_byte_1 : _GEN_248; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_409 = 8'h59 == total_offset_1 ? field_byte_1 : _GEN_249; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_410 = 8'h5a == total_offset_1 ? field_byte_1 : _GEN_250; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_411 = 8'h5b == total_offset_1 ? field_byte_1 : _GEN_251; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_412 = 8'h5c == total_offset_1 ? field_byte_1 : _GEN_252; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_413 = 8'h5d == total_offset_1 ? field_byte_1 : _GEN_253; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_414 = 8'h5e == total_offset_1 ? field_byte_1 : _GEN_254; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_415 = 8'h5f == total_offset_1 ? field_byte_1 : _GEN_255; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_416 = 8'h60 == total_offset_1 ? field_byte_1 : _GEN_256; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_417 = 8'h61 == total_offset_1 ? field_byte_1 : _GEN_257; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_418 = 8'h62 == total_offset_1 ? field_byte_1 : _GEN_258; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_419 = 8'h63 == total_offset_1 ? field_byte_1 : _GEN_259; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_420 = 8'h64 == total_offset_1 ? field_byte_1 : _GEN_260; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_421 = 8'h65 == total_offset_1 ? field_byte_1 : _GEN_261; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_422 = 8'h66 == total_offset_1 ? field_byte_1 : _GEN_262; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_423 = 8'h67 == total_offset_1 ? field_byte_1 : _GEN_263; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_424 = 8'h68 == total_offset_1 ? field_byte_1 : _GEN_264; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_425 = 8'h69 == total_offset_1 ? field_byte_1 : _GEN_265; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_426 = 8'h6a == total_offset_1 ? field_byte_1 : _GEN_266; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_427 = 8'h6b == total_offset_1 ? field_byte_1 : _GEN_267; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_428 = 8'h6c == total_offset_1 ? field_byte_1 : _GEN_268; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_429 = 8'h6d == total_offset_1 ? field_byte_1 : _GEN_269; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_430 = 8'h6e == total_offset_1 ? field_byte_1 : _GEN_270; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_431 = 8'h6f == total_offset_1 ? field_byte_1 : _GEN_271; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_432 = 8'h70 == total_offset_1 ? field_byte_1 : _GEN_272; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_433 = 8'h71 == total_offset_1 ? field_byte_1 : _GEN_273; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_434 = 8'h72 == total_offset_1 ? field_byte_1 : _GEN_274; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_435 = 8'h73 == total_offset_1 ? field_byte_1 : _GEN_275; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_436 = 8'h74 == total_offset_1 ? field_byte_1 : _GEN_276; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_437 = 8'h75 == total_offset_1 ? field_byte_1 : _GEN_277; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_438 = 8'h76 == total_offset_1 ? field_byte_1 : _GEN_278; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_439 = 8'h77 == total_offset_1 ? field_byte_1 : _GEN_279; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_440 = 8'h78 == total_offset_1 ? field_byte_1 : _GEN_280; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_441 = 8'h79 == total_offset_1 ? field_byte_1 : _GEN_281; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_442 = 8'h7a == total_offset_1 ? field_byte_1 : _GEN_282; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_443 = 8'h7b == total_offset_1 ? field_byte_1 : _GEN_283; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_444 = 8'h7c == total_offset_1 ? field_byte_1 : _GEN_284; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_445 = 8'h7d == total_offset_1 ? field_byte_1 : _GEN_285; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_446 = 8'h7e == total_offset_1 ? field_byte_1 : _GEN_286; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_447 = 8'h7f == total_offset_1 ? field_byte_1 : _GEN_287; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_448 = 8'h80 == total_offset_1 ? field_byte_1 : _GEN_288; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_449 = 8'h81 == total_offset_1 ? field_byte_1 : _GEN_289; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_450 = 8'h82 == total_offset_1 ? field_byte_1 : _GEN_290; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_451 = 8'h83 == total_offset_1 ? field_byte_1 : _GEN_291; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_452 = 8'h84 == total_offset_1 ? field_byte_1 : _GEN_292; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_453 = 8'h85 == total_offset_1 ? field_byte_1 : _GEN_293; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_454 = 8'h86 == total_offset_1 ? field_byte_1 : _GEN_294; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_455 = 8'h87 == total_offset_1 ? field_byte_1 : _GEN_295; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_456 = 8'h88 == total_offset_1 ? field_byte_1 : _GEN_296; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_457 = 8'h89 == total_offset_1 ? field_byte_1 : _GEN_297; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_458 = 8'h8a == total_offset_1 ? field_byte_1 : _GEN_298; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_459 = 8'h8b == total_offset_1 ? field_byte_1 : _GEN_299; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_460 = 8'h8c == total_offset_1 ? field_byte_1 : _GEN_300; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_461 = 8'h8d == total_offset_1 ? field_byte_1 : _GEN_301; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_462 = 8'h8e == total_offset_1 ? field_byte_1 : _GEN_302; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_463 = 8'h8f == total_offset_1 ? field_byte_1 : _GEN_303; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_464 = 8'h90 == total_offset_1 ? field_byte_1 : _GEN_304; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_465 = 8'h91 == total_offset_1 ? field_byte_1 : _GEN_305; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_466 = 8'h92 == total_offset_1 ? field_byte_1 : _GEN_306; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_467 = 8'h93 == total_offset_1 ? field_byte_1 : _GEN_307; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_468 = 8'h94 == total_offset_1 ? field_byte_1 : _GEN_308; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_469 = 8'h95 == total_offset_1 ? field_byte_1 : _GEN_309; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_470 = 8'h96 == total_offset_1 ? field_byte_1 : _GEN_310; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_471 = 8'h97 == total_offset_1 ? field_byte_1 : _GEN_311; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_472 = 8'h98 == total_offset_1 ? field_byte_1 : _GEN_312; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_473 = 8'h99 == total_offset_1 ? field_byte_1 : _GEN_313; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_474 = 8'h9a == total_offset_1 ? field_byte_1 : _GEN_314; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_475 = 8'h9b == total_offset_1 ? field_byte_1 : _GEN_315; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_476 = 8'h9c == total_offset_1 ? field_byte_1 : _GEN_316; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_477 = 8'h9d == total_offset_1 ? field_byte_1 : _GEN_317; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_478 = 8'h9e == total_offset_1 ? field_byte_1 : _GEN_318; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_479 = 8'h9f == total_offset_1 ? field_byte_1 : _GEN_319; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_480 = 8'h1 < length_0 ? _GEN_320 : _GEN_160; // @[executor.scala 308:60]
  wire [7:0] _GEN_481 = 8'h1 < length_0 ? _GEN_321 : _GEN_161; // @[executor.scala 308:60]
  wire [7:0] _GEN_482 = 8'h1 < length_0 ? _GEN_322 : _GEN_162; // @[executor.scala 308:60]
  wire [7:0] _GEN_483 = 8'h1 < length_0 ? _GEN_323 : _GEN_163; // @[executor.scala 308:60]
  wire [7:0] _GEN_484 = 8'h1 < length_0 ? _GEN_324 : _GEN_164; // @[executor.scala 308:60]
  wire [7:0] _GEN_485 = 8'h1 < length_0 ? _GEN_325 : _GEN_165; // @[executor.scala 308:60]
  wire [7:0] _GEN_486 = 8'h1 < length_0 ? _GEN_326 : _GEN_166; // @[executor.scala 308:60]
  wire [7:0] _GEN_487 = 8'h1 < length_0 ? _GEN_327 : _GEN_167; // @[executor.scala 308:60]
  wire [7:0] _GEN_488 = 8'h1 < length_0 ? _GEN_328 : _GEN_168; // @[executor.scala 308:60]
  wire [7:0] _GEN_489 = 8'h1 < length_0 ? _GEN_329 : _GEN_169; // @[executor.scala 308:60]
  wire [7:0] _GEN_490 = 8'h1 < length_0 ? _GEN_330 : _GEN_170; // @[executor.scala 308:60]
  wire [7:0] _GEN_491 = 8'h1 < length_0 ? _GEN_331 : _GEN_171; // @[executor.scala 308:60]
  wire [7:0] _GEN_492 = 8'h1 < length_0 ? _GEN_332 : _GEN_172; // @[executor.scala 308:60]
  wire [7:0] _GEN_493 = 8'h1 < length_0 ? _GEN_333 : _GEN_173; // @[executor.scala 308:60]
  wire [7:0] _GEN_494 = 8'h1 < length_0 ? _GEN_334 : _GEN_174; // @[executor.scala 308:60]
  wire [7:0] _GEN_495 = 8'h1 < length_0 ? _GEN_335 : _GEN_175; // @[executor.scala 308:60]
  wire [7:0] _GEN_496 = 8'h1 < length_0 ? _GEN_336 : _GEN_176; // @[executor.scala 308:60]
  wire [7:0] _GEN_497 = 8'h1 < length_0 ? _GEN_337 : _GEN_177; // @[executor.scala 308:60]
  wire [7:0] _GEN_498 = 8'h1 < length_0 ? _GEN_338 : _GEN_178; // @[executor.scala 308:60]
  wire [7:0] _GEN_499 = 8'h1 < length_0 ? _GEN_339 : _GEN_179; // @[executor.scala 308:60]
  wire [7:0] _GEN_500 = 8'h1 < length_0 ? _GEN_340 : _GEN_180; // @[executor.scala 308:60]
  wire [7:0] _GEN_501 = 8'h1 < length_0 ? _GEN_341 : _GEN_181; // @[executor.scala 308:60]
  wire [7:0] _GEN_502 = 8'h1 < length_0 ? _GEN_342 : _GEN_182; // @[executor.scala 308:60]
  wire [7:0] _GEN_503 = 8'h1 < length_0 ? _GEN_343 : _GEN_183; // @[executor.scala 308:60]
  wire [7:0] _GEN_504 = 8'h1 < length_0 ? _GEN_344 : _GEN_184; // @[executor.scala 308:60]
  wire [7:0] _GEN_505 = 8'h1 < length_0 ? _GEN_345 : _GEN_185; // @[executor.scala 308:60]
  wire [7:0] _GEN_506 = 8'h1 < length_0 ? _GEN_346 : _GEN_186; // @[executor.scala 308:60]
  wire [7:0] _GEN_507 = 8'h1 < length_0 ? _GEN_347 : _GEN_187; // @[executor.scala 308:60]
  wire [7:0] _GEN_508 = 8'h1 < length_0 ? _GEN_348 : _GEN_188; // @[executor.scala 308:60]
  wire [7:0] _GEN_509 = 8'h1 < length_0 ? _GEN_349 : _GEN_189; // @[executor.scala 308:60]
  wire [7:0] _GEN_510 = 8'h1 < length_0 ? _GEN_350 : _GEN_190; // @[executor.scala 308:60]
  wire [7:0] _GEN_511 = 8'h1 < length_0 ? _GEN_351 : _GEN_191; // @[executor.scala 308:60]
  wire [7:0] _GEN_512 = 8'h1 < length_0 ? _GEN_352 : _GEN_192; // @[executor.scala 308:60]
  wire [7:0] _GEN_513 = 8'h1 < length_0 ? _GEN_353 : _GEN_193; // @[executor.scala 308:60]
  wire [7:0] _GEN_514 = 8'h1 < length_0 ? _GEN_354 : _GEN_194; // @[executor.scala 308:60]
  wire [7:0] _GEN_515 = 8'h1 < length_0 ? _GEN_355 : _GEN_195; // @[executor.scala 308:60]
  wire [7:0] _GEN_516 = 8'h1 < length_0 ? _GEN_356 : _GEN_196; // @[executor.scala 308:60]
  wire [7:0] _GEN_517 = 8'h1 < length_0 ? _GEN_357 : _GEN_197; // @[executor.scala 308:60]
  wire [7:0] _GEN_518 = 8'h1 < length_0 ? _GEN_358 : _GEN_198; // @[executor.scala 308:60]
  wire [7:0] _GEN_519 = 8'h1 < length_0 ? _GEN_359 : _GEN_199; // @[executor.scala 308:60]
  wire [7:0] _GEN_520 = 8'h1 < length_0 ? _GEN_360 : _GEN_200; // @[executor.scala 308:60]
  wire [7:0] _GEN_521 = 8'h1 < length_0 ? _GEN_361 : _GEN_201; // @[executor.scala 308:60]
  wire [7:0] _GEN_522 = 8'h1 < length_0 ? _GEN_362 : _GEN_202; // @[executor.scala 308:60]
  wire [7:0] _GEN_523 = 8'h1 < length_0 ? _GEN_363 : _GEN_203; // @[executor.scala 308:60]
  wire [7:0] _GEN_524 = 8'h1 < length_0 ? _GEN_364 : _GEN_204; // @[executor.scala 308:60]
  wire [7:0] _GEN_525 = 8'h1 < length_0 ? _GEN_365 : _GEN_205; // @[executor.scala 308:60]
  wire [7:0] _GEN_526 = 8'h1 < length_0 ? _GEN_366 : _GEN_206; // @[executor.scala 308:60]
  wire [7:0] _GEN_527 = 8'h1 < length_0 ? _GEN_367 : _GEN_207; // @[executor.scala 308:60]
  wire [7:0] _GEN_528 = 8'h1 < length_0 ? _GEN_368 : _GEN_208; // @[executor.scala 308:60]
  wire [7:0] _GEN_529 = 8'h1 < length_0 ? _GEN_369 : _GEN_209; // @[executor.scala 308:60]
  wire [7:0] _GEN_530 = 8'h1 < length_0 ? _GEN_370 : _GEN_210; // @[executor.scala 308:60]
  wire [7:0] _GEN_531 = 8'h1 < length_0 ? _GEN_371 : _GEN_211; // @[executor.scala 308:60]
  wire [7:0] _GEN_532 = 8'h1 < length_0 ? _GEN_372 : _GEN_212; // @[executor.scala 308:60]
  wire [7:0] _GEN_533 = 8'h1 < length_0 ? _GEN_373 : _GEN_213; // @[executor.scala 308:60]
  wire [7:0] _GEN_534 = 8'h1 < length_0 ? _GEN_374 : _GEN_214; // @[executor.scala 308:60]
  wire [7:0] _GEN_535 = 8'h1 < length_0 ? _GEN_375 : _GEN_215; // @[executor.scala 308:60]
  wire [7:0] _GEN_536 = 8'h1 < length_0 ? _GEN_376 : _GEN_216; // @[executor.scala 308:60]
  wire [7:0] _GEN_537 = 8'h1 < length_0 ? _GEN_377 : _GEN_217; // @[executor.scala 308:60]
  wire [7:0] _GEN_538 = 8'h1 < length_0 ? _GEN_378 : _GEN_218; // @[executor.scala 308:60]
  wire [7:0] _GEN_539 = 8'h1 < length_0 ? _GEN_379 : _GEN_219; // @[executor.scala 308:60]
  wire [7:0] _GEN_540 = 8'h1 < length_0 ? _GEN_380 : _GEN_220; // @[executor.scala 308:60]
  wire [7:0] _GEN_541 = 8'h1 < length_0 ? _GEN_381 : _GEN_221; // @[executor.scala 308:60]
  wire [7:0] _GEN_542 = 8'h1 < length_0 ? _GEN_382 : _GEN_222; // @[executor.scala 308:60]
  wire [7:0] _GEN_543 = 8'h1 < length_0 ? _GEN_383 : _GEN_223; // @[executor.scala 308:60]
  wire [7:0] _GEN_544 = 8'h1 < length_0 ? _GEN_384 : _GEN_224; // @[executor.scala 308:60]
  wire [7:0] _GEN_545 = 8'h1 < length_0 ? _GEN_385 : _GEN_225; // @[executor.scala 308:60]
  wire [7:0] _GEN_546 = 8'h1 < length_0 ? _GEN_386 : _GEN_226; // @[executor.scala 308:60]
  wire [7:0] _GEN_547 = 8'h1 < length_0 ? _GEN_387 : _GEN_227; // @[executor.scala 308:60]
  wire [7:0] _GEN_548 = 8'h1 < length_0 ? _GEN_388 : _GEN_228; // @[executor.scala 308:60]
  wire [7:0] _GEN_549 = 8'h1 < length_0 ? _GEN_389 : _GEN_229; // @[executor.scala 308:60]
  wire [7:0] _GEN_550 = 8'h1 < length_0 ? _GEN_390 : _GEN_230; // @[executor.scala 308:60]
  wire [7:0] _GEN_551 = 8'h1 < length_0 ? _GEN_391 : _GEN_231; // @[executor.scala 308:60]
  wire [7:0] _GEN_552 = 8'h1 < length_0 ? _GEN_392 : _GEN_232; // @[executor.scala 308:60]
  wire [7:0] _GEN_553 = 8'h1 < length_0 ? _GEN_393 : _GEN_233; // @[executor.scala 308:60]
  wire [7:0] _GEN_554 = 8'h1 < length_0 ? _GEN_394 : _GEN_234; // @[executor.scala 308:60]
  wire [7:0] _GEN_555 = 8'h1 < length_0 ? _GEN_395 : _GEN_235; // @[executor.scala 308:60]
  wire [7:0] _GEN_556 = 8'h1 < length_0 ? _GEN_396 : _GEN_236; // @[executor.scala 308:60]
  wire [7:0] _GEN_557 = 8'h1 < length_0 ? _GEN_397 : _GEN_237; // @[executor.scala 308:60]
  wire [7:0] _GEN_558 = 8'h1 < length_0 ? _GEN_398 : _GEN_238; // @[executor.scala 308:60]
  wire [7:0] _GEN_559 = 8'h1 < length_0 ? _GEN_399 : _GEN_239; // @[executor.scala 308:60]
  wire [7:0] _GEN_560 = 8'h1 < length_0 ? _GEN_400 : _GEN_240; // @[executor.scala 308:60]
  wire [7:0] _GEN_561 = 8'h1 < length_0 ? _GEN_401 : _GEN_241; // @[executor.scala 308:60]
  wire [7:0] _GEN_562 = 8'h1 < length_0 ? _GEN_402 : _GEN_242; // @[executor.scala 308:60]
  wire [7:0] _GEN_563 = 8'h1 < length_0 ? _GEN_403 : _GEN_243; // @[executor.scala 308:60]
  wire [7:0] _GEN_564 = 8'h1 < length_0 ? _GEN_404 : _GEN_244; // @[executor.scala 308:60]
  wire [7:0] _GEN_565 = 8'h1 < length_0 ? _GEN_405 : _GEN_245; // @[executor.scala 308:60]
  wire [7:0] _GEN_566 = 8'h1 < length_0 ? _GEN_406 : _GEN_246; // @[executor.scala 308:60]
  wire [7:0] _GEN_567 = 8'h1 < length_0 ? _GEN_407 : _GEN_247; // @[executor.scala 308:60]
  wire [7:0] _GEN_568 = 8'h1 < length_0 ? _GEN_408 : _GEN_248; // @[executor.scala 308:60]
  wire [7:0] _GEN_569 = 8'h1 < length_0 ? _GEN_409 : _GEN_249; // @[executor.scala 308:60]
  wire [7:0] _GEN_570 = 8'h1 < length_0 ? _GEN_410 : _GEN_250; // @[executor.scala 308:60]
  wire [7:0] _GEN_571 = 8'h1 < length_0 ? _GEN_411 : _GEN_251; // @[executor.scala 308:60]
  wire [7:0] _GEN_572 = 8'h1 < length_0 ? _GEN_412 : _GEN_252; // @[executor.scala 308:60]
  wire [7:0] _GEN_573 = 8'h1 < length_0 ? _GEN_413 : _GEN_253; // @[executor.scala 308:60]
  wire [7:0] _GEN_574 = 8'h1 < length_0 ? _GEN_414 : _GEN_254; // @[executor.scala 308:60]
  wire [7:0] _GEN_575 = 8'h1 < length_0 ? _GEN_415 : _GEN_255; // @[executor.scala 308:60]
  wire [7:0] _GEN_576 = 8'h1 < length_0 ? _GEN_416 : _GEN_256; // @[executor.scala 308:60]
  wire [7:0] _GEN_577 = 8'h1 < length_0 ? _GEN_417 : _GEN_257; // @[executor.scala 308:60]
  wire [7:0] _GEN_578 = 8'h1 < length_0 ? _GEN_418 : _GEN_258; // @[executor.scala 308:60]
  wire [7:0] _GEN_579 = 8'h1 < length_0 ? _GEN_419 : _GEN_259; // @[executor.scala 308:60]
  wire [7:0] _GEN_580 = 8'h1 < length_0 ? _GEN_420 : _GEN_260; // @[executor.scala 308:60]
  wire [7:0] _GEN_581 = 8'h1 < length_0 ? _GEN_421 : _GEN_261; // @[executor.scala 308:60]
  wire [7:0] _GEN_582 = 8'h1 < length_0 ? _GEN_422 : _GEN_262; // @[executor.scala 308:60]
  wire [7:0] _GEN_583 = 8'h1 < length_0 ? _GEN_423 : _GEN_263; // @[executor.scala 308:60]
  wire [7:0] _GEN_584 = 8'h1 < length_0 ? _GEN_424 : _GEN_264; // @[executor.scala 308:60]
  wire [7:0] _GEN_585 = 8'h1 < length_0 ? _GEN_425 : _GEN_265; // @[executor.scala 308:60]
  wire [7:0] _GEN_586 = 8'h1 < length_0 ? _GEN_426 : _GEN_266; // @[executor.scala 308:60]
  wire [7:0] _GEN_587 = 8'h1 < length_0 ? _GEN_427 : _GEN_267; // @[executor.scala 308:60]
  wire [7:0] _GEN_588 = 8'h1 < length_0 ? _GEN_428 : _GEN_268; // @[executor.scala 308:60]
  wire [7:0] _GEN_589 = 8'h1 < length_0 ? _GEN_429 : _GEN_269; // @[executor.scala 308:60]
  wire [7:0] _GEN_590 = 8'h1 < length_0 ? _GEN_430 : _GEN_270; // @[executor.scala 308:60]
  wire [7:0] _GEN_591 = 8'h1 < length_0 ? _GEN_431 : _GEN_271; // @[executor.scala 308:60]
  wire [7:0] _GEN_592 = 8'h1 < length_0 ? _GEN_432 : _GEN_272; // @[executor.scala 308:60]
  wire [7:0] _GEN_593 = 8'h1 < length_0 ? _GEN_433 : _GEN_273; // @[executor.scala 308:60]
  wire [7:0] _GEN_594 = 8'h1 < length_0 ? _GEN_434 : _GEN_274; // @[executor.scala 308:60]
  wire [7:0] _GEN_595 = 8'h1 < length_0 ? _GEN_435 : _GEN_275; // @[executor.scala 308:60]
  wire [7:0] _GEN_596 = 8'h1 < length_0 ? _GEN_436 : _GEN_276; // @[executor.scala 308:60]
  wire [7:0] _GEN_597 = 8'h1 < length_0 ? _GEN_437 : _GEN_277; // @[executor.scala 308:60]
  wire [7:0] _GEN_598 = 8'h1 < length_0 ? _GEN_438 : _GEN_278; // @[executor.scala 308:60]
  wire [7:0] _GEN_599 = 8'h1 < length_0 ? _GEN_439 : _GEN_279; // @[executor.scala 308:60]
  wire [7:0] _GEN_600 = 8'h1 < length_0 ? _GEN_440 : _GEN_280; // @[executor.scala 308:60]
  wire [7:0] _GEN_601 = 8'h1 < length_0 ? _GEN_441 : _GEN_281; // @[executor.scala 308:60]
  wire [7:0] _GEN_602 = 8'h1 < length_0 ? _GEN_442 : _GEN_282; // @[executor.scala 308:60]
  wire [7:0] _GEN_603 = 8'h1 < length_0 ? _GEN_443 : _GEN_283; // @[executor.scala 308:60]
  wire [7:0] _GEN_604 = 8'h1 < length_0 ? _GEN_444 : _GEN_284; // @[executor.scala 308:60]
  wire [7:0] _GEN_605 = 8'h1 < length_0 ? _GEN_445 : _GEN_285; // @[executor.scala 308:60]
  wire [7:0] _GEN_606 = 8'h1 < length_0 ? _GEN_446 : _GEN_286; // @[executor.scala 308:60]
  wire [7:0] _GEN_607 = 8'h1 < length_0 ? _GEN_447 : _GEN_287; // @[executor.scala 308:60]
  wire [7:0] _GEN_608 = 8'h1 < length_0 ? _GEN_448 : _GEN_288; // @[executor.scala 308:60]
  wire [7:0] _GEN_609 = 8'h1 < length_0 ? _GEN_449 : _GEN_289; // @[executor.scala 308:60]
  wire [7:0] _GEN_610 = 8'h1 < length_0 ? _GEN_450 : _GEN_290; // @[executor.scala 308:60]
  wire [7:0] _GEN_611 = 8'h1 < length_0 ? _GEN_451 : _GEN_291; // @[executor.scala 308:60]
  wire [7:0] _GEN_612 = 8'h1 < length_0 ? _GEN_452 : _GEN_292; // @[executor.scala 308:60]
  wire [7:0] _GEN_613 = 8'h1 < length_0 ? _GEN_453 : _GEN_293; // @[executor.scala 308:60]
  wire [7:0] _GEN_614 = 8'h1 < length_0 ? _GEN_454 : _GEN_294; // @[executor.scala 308:60]
  wire [7:0] _GEN_615 = 8'h1 < length_0 ? _GEN_455 : _GEN_295; // @[executor.scala 308:60]
  wire [7:0] _GEN_616 = 8'h1 < length_0 ? _GEN_456 : _GEN_296; // @[executor.scala 308:60]
  wire [7:0] _GEN_617 = 8'h1 < length_0 ? _GEN_457 : _GEN_297; // @[executor.scala 308:60]
  wire [7:0] _GEN_618 = 8'h1 < length_0 ? _GEN_458 : _GEN_298; // @[executor.scala 308:60]
  wire [7:0] _GEN_619 = 8'h1 < length_0 ? _GEN_459 : _GEN_299; // @[executor.scala 308:60]
  wire [7:0] _GEN_620 = 8'h1 < length_0 ? _GEN_460 : _GEN_300; // @[executor.scala 308:60]
  wire [7:0] _GEN_621 = 8'h1 < length_0 ? _GEN_461 : _GEN_301; // @[executor.scala 308:60]
  wire [7:0] _GEN_622 = 8'h1 < length_0 ? _GEN_462 : _GEN_302; // @[executor.scala 308:60]
  wire [7:0] _GEN_623 = 8'h1 < length_0 ? _GEN_463 : _GEN_303; // @[executor.scala 308:60]
  wire [7:0] _GEN_624 = 8'h1 < length_0 ? _GEN_464 : _GEN_304; // @[executor.scala 308:60]
  wire [7:0] _GEN_625 = 8'h1 < length_0 ? _GEN_465 : _GEN_305; // @[executor.scala 308:60]
  wire [7:0] _GEN_626 = 8'h1 < length_0 ? _GEN_466 : _GEN_306; // @[executor.scala 308:60]
  wire [7:0] _GEN_627 = 8'h1 < length_0 ? _GEN_467 : _GEN_307; // @[executor.scala 308:60]
  wire [7:0] _GEN_628 = 8'h1 < length_0 ? _GEN_468 : _GEN_308; // @[executor.scala 308:60]
  wire [7:0] _GEN_629 = 8'h1 < length_0 ? _GEN_469 : _GEN_309; // @[executor.scala 308:60]
  wire [7:0] _GEN_630 = 8'h1 < length_0 ? _GEN_470 : _GEN_310; // @[executor.scala 308:60]
  wire [7:0] _GEN_631 = 8'h1 < length_0 ? _GEN_471 : _GEN_311; // @[executor.scala 308:60]
  wire [7:0] _GEN_632 = 8'h1 < length_0 ? _GEN_472 : _GEN_312; // @[executor.scala 308:60]
  wire [7:0] _GEN_633 = 8'h1 < length_0 ? _GEN_473 : _GEN_313; // @[executor.scala 308:60]
  wire [7:0] _GEN_634 = 8'h1 < length_0 ? _GEN_474 : _GEN_314; // @[executor.scala 308:60]
  wire [7:0] _GEN_635 = 8'h1 < length_0 ? _GEN_475 : _GEN_315; // @[executor.scala 308:60]
  wire [7:0] _GEN_636 = 8'h1 < length_0 ? _GEN_476 : _GEN_316; // @[executor.scala 308:60]
  wire [7:0] _GEN_637 = 8'h1 < length_0 ? _GEN_477 : _GEN_317; // @[executor.scala 308:60]
  wire [7:0] _GEN_638 = 8'h1 < length_0 ? _GEN_478 : _GEN_318; // @[executor.scala 308:60]
  wire [7:0] _GEN_639 = 8'h1 < length_0 ? _GEN_479 : _GEN_319; // @[executor.scala 308:60]
  wire [7:0] field_byte_2 = field_0[47:40]; // @[executor.scala 305:57]
  wire [7:0] total_offset_2 = offset_0 + 8'h2; // @[executor.scala 307:57]
  wire [7:0] _GEN_640 = 8'h0 == total_offset_2 ? field_byte_2 : _GEN_480; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_641 = 8'h1 == total_offset_2 ? field_byte_2 : _GEN_481; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_642 = 8'h2 == total_offset_2 ? field_byte_2 : _GEN_482; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_643 = 8'h3 == total_offset_2 ? field_byte_2 : _GEN_483; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_644 = 8'h4 == total_offset_2 ? field_byte_2 : _GEN_484; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_645 = 8'h5 == total_offset_2 ? field_byte_2 : _GEN_485; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_646 = 8'h6 == total_offset_2 ? field_byte_2 : _GEN_486; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_647 = 8'h7 == total_offset_2 ? field_byte_2 : _GEN_487; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_648 = 8'h8 == total_offset_2 ? field_byte_2 : _GEN_488; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_649 = 8'h9 == total_offset_2 ? field_byte_2 : _GEN_489; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_650 = 8'ha == total_offset_2 ? field_byte_2 : _GEN_490; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_651 = 8'hb == total_offset_2 ? field_byte_2 : _GEN_491; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_652 = 8'hc == total_offset_2 ? field_byte_2 : _GEN_492; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_653 = 8'hd == total_offset_2 ? field_byte_2 : _GEN_493; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_654 = 8'he == total_offset_2 ? field_byte_2 : _GEN_494; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_655 = 8'hf == total_offset_2 ? field_byte_2 : _GEN_495; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_656 = 8'h10 == total_offset_2 ? field_byte_2 : _GEN_496; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_657 = 8'h11 == total_offset_2 ? field_byte_2 : _GEN_497; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_658 = 8'h12 == total_offset_2 ? field_byte_2 : _GEN_498; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_659 = 8'h13 == total_offset_2 ? field_byte_2 : _GEN_499; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_660 = 8'h14 == total_offset_2 ? field_byte_2 : _GEN_500; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_661 = 8'h15 == total_offset_2 ? field_byte_2 : _GEN_501; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_662 = 8'h16 == total_offset_2 ? field_byte_2 : _GEN_502; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_663 = 8'h17 == total_offset_2 ? field_byte_2 : _GEN_503; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_664 = 8'h18 == total_offset_2 ? field_byte_2 : _GEN_504; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_665 = 8'h19 == total_offset_2 ? field_byte_2 : _GEN_505; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_666 = 8'h1a == total_offset_2 ? field_byte_2 : _GEN_506; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_667 = 8'h1b == total_offset_2 ? field_byte_2 : _GEN_507; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_668 = 8'h1c == total_offset_2 ? field_byte_2 : _GEN_508; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_669 = 8'h1d == total_offset_2 ? field_byte_2 : _GEN_509; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_670 = 8'h1e == total_offset_2 ? field_byte_2 : _GEN_510; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_671 = 8'h1f == total_offset_2 ? field_byte_2 : _GEN_511; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_672 = 8'h20 == total_offset_2 ? field_byte_2 : _GEN_512; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_673 = 8'h21 == total_offset_2 ? field_byte_2 : _GEN_513; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_674 = 8'h22 == total_offset_2 ? field_byte_2 : _GEN_514; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_675 = 8'h23 == total_offset_2 ? field_byte_2 : _GEN_515; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_676 = 8'h24 == total_offset_2 ? field_byte_2 : _GEN_516; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_677 = 8'h25 == total_offset_2 ? field_byte_2 : _GEN_517; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_678 = 8'h26 == total_offset_2 ? field_byte_2 : _GEN_518; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_679 = 8'h27 == total_offset_2 ? field_byte_2 : _GEN_519; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_680 = 8'h28 == total_offset_2 ? field_byte_2 : _GEN_520; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_681 = 8'h29 == total_offset_2 ? field_byte_2 : _GEN_521; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_682 = 8'h2a == total_offset_2 ? field_byte_2 : _GEN_522; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_683 = 8'h2b == total_offset_2 ? field_byte_2 : _GEN_523; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_684 = 8'h2c == total_offset_2 ? field_byte_2 : _GEN_524; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_685 = 8'h2d == total_offset_2 ? field_byte_2 : _GEN_525; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_686 = 8'h2e == total_offset_2 ? field_byte_2 : _GEN_526; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_687 = 8'h2f == total_offset_2 ? field_byte_2 : _GEN_527; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_688 = 8'h30 == total_offset_2 ? field_byte_2 : _GEN_528; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_689 = 8'h31 == total_offset_2 ? field_byte_2 : _GEN_529; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_690 = 8'h32 == total_offset_2 ? field_byte_2 : _GEN_530; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_691 = 8'h33 == total_offset_2 ? field_byte_2 : _GEN_531; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_692 = 8'h34 == total_offset_2 ? field_byte_2 : _GEN_532; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_693 = 8'h35 == total_offset_2 ? field_byte_2 : _GEN_533; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_694 = 8'h36 == total_offset_2 ? field_byte_2 : _GEN_534; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_695 = 8'h37 == total_offset_2 ? field_byte_2 : _GEN_535; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_696 = 8'h38 == total_offset_2 ? field_byte_2 : _GEN_536; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_697 = 8'h39 == total_offset_2 ? field_byte_2 : _GEN_537; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_698 = 8'h3a == total_offset_2 ? field_byte_2 : _GEN_538; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_699 = 8'h3b == total_offset_2 ? field_byte_2 : _GEN_539; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_700 = 8'h3c == total_offset_2 ? field_byte_2 : _GEN_540; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_701 = 8'h3d == total_offset_2 ? field_byte_2 : _GEN_541; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_702 = 8'h3e == total_offset_2 ? field_byte_2 : _GEN_542; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_703 = 8'h3f == total_offset_2 ? field_byte_2 : _GEN_543; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_704 = 8'h40 == total_offset_2 ? field_byte_2 : _GEN_544; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_705 = 8'h41 == total_offset_2 ? field_byte_2 : _GEN_545; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_706 = 8'h42 == total_offset_2 ? field_byte_2 : _GEN_546; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_707 = 8'h43 == total_offset_2 ? field_byte_2 : _GEN_547; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_708 = 8'h44 == total_offset_2 ? field_byte_2 : _GEN_548; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_709 = 8'h45 == total_offset_2 ? field_byte_2 : _GEN_549; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_710 = 8'h46 == total_offset_2 ? field_byte_2 : _GEN_550; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_711 = 8'h47 == total_offset_2 ? field_byte_2 : _GEN_551; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_712 = 8'h48 == total_offset_2 ? field_byte_2 : _GEN_552; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_713 = 8'h49 == total_offset_2 ? field_byte_2 : _GEN_553; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_714 = 8'h4a == total_offset_2 ? field_byte_2 : _GEN_554; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_715 = 8'h4b == total_offset_2 ? field_byte_2 : _GEN_555; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_716 = 8'h4c == total_offset_2 ? field_byte_2 : _GEN_556; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_717 = 8'h4d == total_offset_2 ? field_byte_2 : _GEN_557; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_718 = 8'h4e == total_offset_2 ? field_byte_2 : _GEN_558; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_719 = 8'h4f == total_offset_2 ? field_byte_2 : _GEN_559; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_720 = 8'h50 == total_offset_2 ? field_byte_2 : _GEN_560; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_721 = 8'h51 == total_offset_2 ? field_byte_2 : _GEN_561; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_722 = 8'h52 == total_offset_2 ? field_byte_2 : _GEN_562; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_723 = 8'h53 == total_offset_2 ? field_byte_2 : _GEN_563; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_724 = 8'h54 == total_offset_2 ? field_byte_2 : _GEN_564; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_725 = 8'h55 == total_offset_2 ? field_byte_2 : _GEN_565; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_726 = 8'h56 == total_offset_2 ? field_byte_2 : _GEN_566; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_727 = 8'h57 == total_offset_2 ? field_byte_2 : _GEN_567; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_728 = 8'h58 == total_offset_2 ? field_byte_2 : _GEN_568; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_729 = 8'h59 == total_offset_2 ? field_byte_2 : _GEN_569; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_730 = 8'h5a == total_offset_2 ? field_byte_2 : _GEN_570; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_731 = 8'h5b == total_offset_2 ? field_byte_2 : _GEN_571; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_732 = 8'h5c == total_offset_2 ? field_byte_2 : _GEN_572; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_733 = 8'h5d == total_offset_2 ? field_byte_2 : _GEN_573; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_734 = 8'h5e == total_offset_2 ? field_byte_2 : _GEN_574; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_735 = 8'h5f == total_offset_2 ? field_byte_2 : _GEN_575; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_736 = 8'h60 == total_offset_2 ? field_byte_2 : _GEN_576; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_737 = 8'h61 == total_offset_2 ? field_byte_2 : _GEN_577; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_738 = 8'h62 == total_offset_2 ? field_byte_2 : _GEN_578; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_739 = 8'h63 == total_offset_2 ? field_byte_2 : _GEN_579; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_740 = 8'h64 == total_offset_2 ? field_byte_2 : _GEN_580; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_741 = 8'h65 == total_offset_2 ? field_byte_2 : _GEN_581; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_742 = 8'h66 == total_offset_2 ? field_byte_2 : _GEN_582; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_743 = 8'h67 == total_offset_2 ? field_byte_2 : _GEN_583; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_744 = 8'h68 == total_offset_2 ? field_byte_2 : _GEN_584; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_745 = 8'h69 == total_offset_2 ? field_byte_2 : _GEN_585; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_746 = 8'h6a == total_offset_2 ? field_byte_2 : _GEN_586; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_747 = 8'h6b == total_offset_2 ? field_byte_2 : _GEN_587; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_748 = 8'h6c == total_offset_2 ? field_byte_2 : _GEN_588; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_749 = 8'h6d == total_offset_2 ? field_byte_2 : _GEN_589; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_750 = 8'h6e == total_offset_2 ? field_byte_2 : _GEN_590; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_751 = 8'h6f == total_offset_2 ? field_byte_2 : _GEN_591; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_752 = 8'h70 == total_offset_2 ? field_byte_2 : _GEN_592; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_753 = 8'h71 == total_offset_2 ? field_byte_2 : _GEN_593; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_754 = 8'h72 == total_offset_2 ? field_byte_2 : _GEN_594; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_755 = 8'h73 == total_offset_2 ? field_byte_2 : _GEN_595; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_756 = 8'h74 == total_offset_2 ? field_byte_2 : _GEN_596; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_757 = 8'h75 == total_offset_2 ? field_byte_2 : _GEN_597; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_758 = 8'h76 == total_offset_2 ? field_byte_2 : _GEN_598; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_759 = 8'h77 == total_offset_2 ? field_byte_2 : _GEN_599; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_760 = 8'h78 == total_offset_2 ? field_byte_2 : _GEN_600; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_761 = 8'h79 == total_offset_2 ? field_byte_2 : _GEN_601; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_762 = 8'h7a == total_offset_2 ? field_byte_2 : _GEN_602; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_763 = 8'h7b == total_offset_2 ? field_byte_2 : _GEN_603; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_764 = 8'h7c == total_offset_2 ? field_byte_2 : _GEN_604; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_765 = 8'h7d == total_offset_2 ? field_byte_2 : _GEN_605; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_766 = 8'h7e == total_offset_2 ? field_byte_2 : _GEN_606; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_767 = 8'h7f == total_offset_2 ? field_byte_2 : _GEN_607; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_768 = 8'h80 == total_offset_2 ? field_byte_2 : _GEN_608; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_769 = 8'h81 == total_offset_2 ? field_byte_2 : _GEN_609; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_770 = 8'h82 == total_offset_2 ? field_byte_2 : _GEN_610; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_771 = 8'h83 == total_offset_2 ? field_byte_2 : _GEN_611; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_772 = 8'h84 == total_offset_2 ? field_byte_2 : _GEN_612; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_773 = 8'h85 == total_offset_2 ? field_byte_2 : _GEN_613; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_774 = 8'h86 == total_offset_2 ? field_byte_2 : _GEN_614; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_775 = 8'h87 == total_offset_2 ? field_byte_2 : _GEN_615; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_776 = 8'h88 == total_offset_2 ? field_byte_2 : _GEN_616; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_777 = 8'h89 == total_offset_2 ? field_byte_2 : _GEN_617; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_778 = 8'h8a == total_offset_2 ? field_byte_2 : _GEN_618; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_779 = 8'h8b == total_offset_2 ? field_byte_2 : _GEN_619; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_780 = 8'h8c == total_offset_2 ? field_byte_2 : _GEN_620; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_781 = 8'h8d == total_offset_2 ? field_byte_2 : _GEN_621; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_782 = 8'h8e == total_offset_2 ? field_byte_2 : _GEN_622; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_783 = 8'h8f == total_offset_2 ? field_byte_2 : _GEN_623; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_784 = 8'h90 == total_offset_2 ? field_byte_2 : _GEN_624; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_785 = 8'h91 == total_offset_2 ? field_byte_2 : _GEN_625; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_786 = 8'h92 == total_offset_2 ? field_byte_2 : _GEN_626; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_787 = 8'h93 == total_offset_2 ? field_byte_2 : _GEN_627; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_788 = 8'h94 == total_offset_2 ? field_byte_2 : _GEN_628; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_789 = 8'h95 == total_offset_2 ? field_byte_2 : _GEN_629; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_790 = 8'h96 == total_offset_2 ? field_byte_2 : _GEN_630; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_791 = 8'h97 == total_offset_2 ? field_byte_2 : _GEN_631; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_792 = 8'h98 == total_offset_2 ? field_byte_2 : _GEN_632; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_793 = 8'h99 == total_offset_2 ? field_byte_2 : _GEN_633; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_794 = 8'h9a == total_offset_2 ? field_byte_2 : _GEN_634; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_795 = 8'h9b == total_offset_2 ? field_byte_2 : _GEN_635; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_796 = 8'h9c == total_offset_2 ? field_byte_2 : _GEN_636; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_797 = 8'h9d == total_offset_2 ? field_byte_2 : _GEN_637; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_798 = 8'h9e == total_offset_2 ? field_byte_2 : _GEN_638; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_799 = 8'h9f == total_offset_2 ? field_byte_2 : _GEN_639; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_800 = 8'h2 < length_0 ? _GEN_640 : _GEN_480; // @[executor.scala 308:60]
  wire [7:0] _GEN_801 = 8'h2 < length_0 ? _GEN_641 : _GEN_481; // @[executor.scala 308:60]
  wire [7:0] _GEN_802 = 8'h2 < length_0 ? _GEN_642 : _GEN_482; // @[executor.scala 308:60]
  wire [7:0] _GEN_803 = 8'h2 < length_0 ? _GEN_643 : _GEN_483; // @[executor.scala 308:60]
  wire [7:0] _GEN_804 = 8'h2 < length_0 ? _GEN_644 : _GEN_484; // @[executor.scala 308:60]
  wire [7:0] _GEN_805 = 8'h2 < length_0 ? _GEN_645 : _GEN_485; // @[executor.scala 308:60]
  wire [7:0] _GEN_806 = 8'h2 < length_0 ? _GEN_646 : _GEN_486; // @[executor.scala 308:60]
  wire [7:0] _GEN_807 = 8'h2 < length_0 ? _GEN_647 : _GEN_487; // @[executor.scala 308:60]
  wire [7:0] _GEN_808 = 8'h2 < length_0 ? _GEN_648 : _GEN_488; // @[executor.scala 308:60]
  wire [7:0] _GEN_809 = 8'h2 < length_0 ? _GEN_649 : _GEN_489; // @[executor.scala 308:60]
  wire [7:0] _GEN_810 = 8'h2 < length_0 ? _GEN_650 : _GEN_490; // @[executor.scala 308:60]
  wire [7:0] _GEN_811 = 8'h2 < length_0 ? _GEN_651 : _GEN_491; // @[executor.scala 308:60]
  wire [7:0] _GEN_812 = 8'h2 < length_0 ? _GEN_652 : _GEN_492; // @[executor.scala 308:60]
  wire [7:0] _GEN_813 = 8'h2 < length_0 ? _GEN_653 : _GEN_493; // @[executor.scala 308:60]
  wire [7:0] _GEN_814 = 8'h2 < length_0 ? _GEN_654 : _GEN_494; // @[executor.scala 308:60]
  wire [7:0] _GEN_815 = 8'h2 < length_0 ? _GEN_655 : _GEN_495; // @[executor.scala 308:60]
  wire [7:0] _GEN_816 = 8'h2 < length_0 ? _GEN_656 : _GEN_496; // @[executor.scala 308:60]
  wire [7:0] _GEN_817 = 8'h2 < length_0 ? _GEN_657 : _GEN_497; // @[executor.scala 308:60]
  wire [7:0] _GEN_818 = 8'h2 < length_0 ? _GEN_658 : _GEN_498; // @[executor.scala 308:60]
  wire [7:0] _GEN_819 = 8'h2 < length_0 ? _GEN_659 : _GEN_499; // @[executor.scala 308:60]
  wire [7:0] _GEN_820 = 8'h2 < length_0 ? _GEN_660 : _GEN_500; // @[executor.scala 308:60]
  wire [7:0] _GEN_821 = 8'h2 < length_0 ? _GEN_661 : _GEN_501; // @[executor.scala 308:60]
  wire [7:0] _GEN_822 = 8'h2 < length_0 ? _GEN_662 : _GEN_502; // @[executor.scala 308:60]
  wire [7:0] _GEN_823 = 8'h2 < length_0 ? _GEN_663 : _GEN_503; // @[executor.scala 308:60]
  wire [7:0] _GEN_824 = 8'h2 < length_0 ? _GEN_664 : _GEN_504; // @[executor.scala 308:60]
  wire [7:0] _GEN_825 = 8'h2 < length_0 ? _GEN_665 : _GEN_505; // @[executor.scala 308:60]
  wire [7:0] _GEN_826 = 8'h2 < length_0 ? _GEN_666 : _GEN_506; // @[executor.scala 308:60]
  wire [7:0] _GEN_827 = 8'h2 < length_0 ? _GEN_667 : _GEN_507; // @[executor.scala 308:60]
  wire [7:0] _GEN_828 = 8'h2 < length_0 ? _GEN_668 : _GEN_508; // @[executor.scala 308:60]
  wire [7:0] _GEN_829 = 8'h2 < length_0 ? _GEN_669 : _GEN_509; // @[executor.scala 308:60]
  wire [7:0] _GEN_830 = 8'h2 < length_0 ? _GEN_670 : _GEN_510; // @[executor.scala 308:60]
  wire [7:0] _GEN_831 = 8'h2 < length_0 ? _GEN_671 : _GEN_511; // @[executor.scala 308:60]
  wire [7:0] _GEN_832 = 8'h2 < length_0 ? _GEN_672 : _GEN_512; // @[executor.scala 308:60]
  wire [7:0] _GEN_833 = 8'h2 < length_0 ? _GEN_673 : _GEN_513; // @[executor.scala 308:60]
  wire [7:0] _GEN_834 = 8'h2 < length_0 ? _GEN_674 : _GEN_514; // @[executor.scala 308:60]
  wire [7:0] _GEN_835 = 8'h2 < length_0 ? _GEN_675 : _GEN_515; // @[executor.scala 308:60]
  wire [7:0] _GEN_836 = 8'h2 < length_0 ? _GEN_676 : _GEN_516; // @[executor.scala 308:60]
  wire [7:0] _GEN_837 = 8'h2 < length_0 ? _GEN_677 : _GEN_517; // @[executor.scala 308:60]
  wire [7:0] _GEN_838 = 8'h2 < length_0 ? _GEN_678 : _GEN_518; // @[executor.scala 308:60]
  wire [7:0] _GEN_839 = 8'h2 < length_0 ? _GEN_679 : _GEN_519; // @[executor.scala 308:60]
  wire [7:0] _GEN_840 = 8'h2 < length_0 ? _GEN_680 : _GEN_520; // @[executor.scala 308:60]
  wire [7:0] _GEN_841 = 8'h2 < length_0 ? _GEN_681 : _GEN_521; // @[executor.scala 308:60]
  wire [7:0] _GEN_842 = 8'h2 < length_0 ? _GEN_682 : _GEN_522; // @[executor.scala 308:60]
  wire [7:0] _GEN_843 = 8'h2 < length_0 ? _GEN_683 : _GEN_523; // @[executor.scala 308:60]
  wire [7:0] _GEN_844 = 8'h2 < length_0 ? _GEN_684 : _GEN_524; // @[executor.scala 308:60]
  wire [7:0] _GEN_845 = 8'h2 < length_0 ? _GEN_685 : _GEN_525; // @[executor.scala 308:60]
  wire [7:0] _GEN_846 = 8'h2 < length_0 ? _GEN_686 : _GEN_526; // @[executor.scala 308:60]
  wire [7:0] _GEN_847 = 8'h2 < length_0 ? _GEN_687 : _GEN_527; // @[executor.scala 308:60]
  wire [7:0] _GEN_848 = 8'h2 < length_0 ? _GEN_688 : _GEN_528; // @[executor.scala 308:60]
  wire [7:0] _GEN_849 = 8'h2 < length_0 ? _GEN_689 : _GEN_529; // @[executor.scala 308:60]
  wire [7:0] _GEN_850 = 8'h2 < length_0 ? _GEN_690 : _GEN_530; // @[executor.scala 308:60]
  wire [7:0] _GEN_851 = 8'h2 < length_0 ? _GEN_691 : _GEN_531; // @[executor.scala 308:60]
  wire [7:0] _GEN_852 = 8'h2 < length_0 ? _GEN_692 : _GEN_532; // @[executor.scala 308:60]
  wire [7:0] _GEN_853 = 8'h2 < length_0 ? _GEN_693 : _GEN_533; // @[executor.scala 308:60]
  wire [7:0] _GEN_854 = 8'h2 < length_0 ? _GEN_694 : _GEN_534; // @[executor.scala 308:60]
  wire [7:0] _GEN_855 = 8'h2 < length_0 ? _GEN_695 : _GEN_535; // @[executor.scala 308:60]
  wire [7:0] _GEN_856 = 8'h2 < length_0 ? _GEN_696 : _GEN_536; // @[executor.scala 308:60]
  wire [7:0] _GEN_857 = 8'h2 < length_0 ? _GEN_697 : _GEN_537; // @[executor.scala 308:60]
  wire [7:0] _GEN_858 = 8'h2 < length_0 ? _GEN_698 : _GEN_538; // @[executor.scala 308:60]
  wire [7:0] _GEN_859 = 8'h2 < length_0 ? _GEN_699 : _GEN_539; // @[executor.scala 308:60]
  wire [7:0] _GEN_860 = 8'h2 < length_0 ? _GEN_700 : _GEN_540; // @[executor.scala 308:60]
  wire [7:0] _GEN_861 = 8'h2 < length_0 ? _GEN_701 : _GEN_541; // @[executor.scala 308:60]
  wire [7:0] _GEN_862 = 8'h2 < length_0 ? _GEN_702 : _GEN_542; // @[executor.scala 308:60]
  wire [7:0] _GEN_863 = 8'h2 < length_0 ? _GEN_703 : _GEN_543; // @[executor.scala 308:60]
  wire [7:0] _GEN_864 = 8'h2 < length_0 ? _GEN_704 : _GEN_544; // @[executor.scala 308:60]
  wire [7:0] _GEN_865 = 8'h2 < length_0 ? _GEN_705 : _GEN_545; // @[executor.scala 308:60]
  wire [7:0] _GEN_866 = 8'h2 < length_0 ? _GEN_706 : _GEN_546; // @[executor.scala 308:60]
  wire [7:0] _GEN_867 = 8'h2 < length_0 ? _GEN_707 : _GEN_547; // @[executor.scala 308:60]
  wire [7:0] _GEN_868 = 8'h2 < length_0 ? _GEN_708 : _GEN_548; // @[executor.scala 308:60]
  wire [7:0] _GEN_869 = 8'h2 < length_0 ? _GEN_709 : _GEN_549; // @[executor.scala 308:60]
  wire [7:0] _GEN_870 = 8'h2 < length_0 ? _GEN_710 : _GEN_550; // @[executor.scala 308:60]
  wire [7:0] _GEN_871 = 8'h2 < length_0 ? _GEN_711 : _GEN_551; // @[executor.scala 308:60]
  wire [7:0] _GEN_872 = 8'h2 < length_0 ? _GEN_712 : _GEN_552; // @[executor.scala 308:60]
  wire [7:0] _GEN_873 = 8'h2 < length_0 ? _GEN_713 : _GEN_553; // @[executor.scala 308:60]
  wire [7:0] _GEN_874 = 8'h2 < length_0 ? _GEN_714 : _GEN_554; // @[executor.scala 308:60]
  wire [7:0] _GEN_875 = 8'h2 < length_0 ? _GEN_715 : _GEN_555; // @[executor.scala 308:60]
  wire [7:0] _GEN_876 = 8'h2 < length_0 ? _GEN_716 : _GEN_556; // @[executor.scala 308:60]
  wire [7:0] _GEN_877 = 8'h2 < length_0 ? _GEN_717 : _GEN_557; // @[executor.scala 308:60]
  wire [7:0] _GEN_878 = 8'h2 < length_0 ? _GEN_718 : _GEN_558; // @[executor.scala 308:60]
  wire [7:0] _GEN_879 = 8'h2 < length_0 ? _GEN_719 : _GEN_559; // @[executor.scala 308:60]
  wire [7:0] _GEN_880 = 8'h2 < length_0 ? _GEN_720 : _GEN_560; // @[executor.scala 308:60]
  wire [7:0] _GEN_881 = 8'h2 < length_0 ? _GEN_721 : _GEN_561; // @[executor.scala 308:60]
  wire [7:0] _GEN_882 = 8'h2 < length_0 ? _GEN_722 : _GEN_562; // @[executor.scala 308:60]
  wire [7:0] _GEN_883 = 8'h2 < length_0 ? _GEN_723 : _GEN_563; // @[executor.scala 308:60]
  wire [7:0] _GEN_884 = 8'h2 < length_0 ? _GEN_724 : _GEN_564; // @[executor.scala 308:60]
  wire [7:0] _GEN_885 = 8'h2 < length_0 ? _GEN_725 : _GEN_565; // @[executor.scala 308:60]
  wire [7:0] _GEN_886 = 8'h2 < length_0 ? _GEN_726 : _GEN_566; // @[executor.scala 308:60]
  wire [7:0] _GEN_887 = 8'h2 < length_0 ? _GEN_727 : _GEN_567; // @[executor.scala 308:60]
  wire [7:0] _GEN_888 = 8'h2 < length_0 ? _GEN_728 : _GEN_568; // @[executor.scala 308:60]
  wire [7:0] _GEN_889 = 8'h2 < length_0 ? _GEN_729 : _GEN_569; // @[executor.scala 308:60]
  wire [7:0] _GEN_890 = 8'h2 < length_0 ? _GEN_730 : _GEN_570; // @[executor.scala 308:60]
  wire [7:0] _GEN_891 = 8'h2 < length_0 ? _GEN_731 : _GEN_571; // @[executor.scala 308:60]
  wire [7:0] _GEN_892 = 8'h2 < length_0 ? _GEN_732 : _GEN_572; // @[executor.scala 308:60]
  wire [7:0] _GEN_893 = 8'h2 < length_0 ? _GEN_733 : _GEN_573; // @[executor.scala 308:60]
  wire [7:0] _GEN_894 = 8'h2 < length_0 ? _GEN_734 : _GEN_574; // @[executor.scala 308:60]
  wire [7:0] _GEN_895 = 8'h2 < length_0 ? _GEN_735 : _GEN_575; // @[executor.scala 308:60]
  wire [7:0] _GEN_896 = 8'h2 < length_0 ? _GEN_736 : _GEN_576; // @[executor.scala 308:60]
  wire [7:0] _GEN_897 = 8'h2 < length_0 ? _GEN_737 : _GEN_577; // @[executor.scala 308:60]
  wire [7:0] _GEN_898 = 8'h2 < length_0 ? _GEN_738 : _GEN_578; // @[executor.scala 308:60]
  wire [7:0] _GEN_899 = 8'h2 < length_0 ? _GEN_739 : _GEN_579; // @[executor.scala 308:60]
  wire [7:0] _GEN_900 = 8'h2 < length_0 ? _GEN_740 : _GEN_580; // @[executor.scala 308:60]
  wire [7:0] _GEN_901 = 8'h2 < length_0 ? _GEN_741 : _GEN_581; // @[executor.scala 308:60]
  wire [7:0] _GEN_902 = 8'h2 < length_0 ? _GEN_742 : _GEN_582; // @[executor.scala 308:60]
  wire [7:0] _GEN_903 = 8'h2 < length_0 ? _GEN_743 : _GEN_583; // @[executor.scala 308:60]
  wire [7:0] _GEN_904 = 8'h2 < length_0 ? _GEN_744 : _GEN_584; // @[executor.scala 308:60]
  wire [7:0] _GEN_905 = 8'h2 < length_0 ? _GEN_745 : _GEN_585; // @[executor.scala 308:60]
  wire [7:0] _GEN_906 = 8'h2 < length_0 ? _GEN_746 : _GEN_586; // @[executor.scala 308:60]
  wire [7:0] _GEN_907 = 8'h2 < length_0 ? _GEN_747 : _GEN_587; // @[executor.scala 308:60]
  wire [7:0] _GEN_908 = 8'h2 < length_0 ? _GEN_748 : _GEN_588; // @[executor.scala 308:60]
  wire [7:0] _GEN_909 = 8'h2 < length_0 ? _GEN_749 : _GEN_589; // @[executor.scala 308:60]
  wire [7:0] _GEN_910 = 8'h2 < length_0 ? _GEN_750 : _GEN_590; // @[executor.scala 308:60]
  wire [7:0] _GEN_911 = 8'h2 < length_0 ? _GEN_751 : _GEN_591; // @[executor.scala 308:60]
  wire [7:0] _GEN_912 = 8'h2 < length_0 ? _GEN_752 : _GEN_592; // @[executor.scala 308:60]
  wire [7:0] _GEN_913 = 8'h2 < length_0 ? _GEN_753 : _GEN_593; // @[executor.scala 308:60]
  wire [7:0] _GEN_914 = 8'h2 < length_0 ? _GEN_754 : _GEN_594; // @[executor.scala 308:60]
  wire [7:0] _GEN_915 = 8'h2 < length_0 ? _GEN_755 : _GEN_595; // @[executor.scala 308:60]
  wire [7:0] _GEN_916 = 8'h2 < length_0 ? _GEN_756 : _GEN_596; // @[executor.scala 308:60]
  wire [7:0] _GEN_917 = 8'h2 < length_0 ? _GEN_757 : _GEN_597; // @[executor.scala 308:60]
  wire [7:0] _GEN_918 = 8'h2 < length_0 ? _GEN_758 : _GEN_598; // @[executor.scala 308:60]
  wire [7:0] _GEN_919 = 8'h2 < length_0 ? _GEN_759 : _GEN_599; // @[executor.scala 308:60]
  wire [7:0] _GEN_920 = 8'h2 < length_0 ? _GEN_760 : _GEN_600; // @[executor.scala 308:60]
  wire [7:0] _GEN_921 = 8'h2 < length_0 ? _GEN_761 : _GEN_601; // @[executor.scala 308:60]
  wire [7:0] _GEN_922 = 8'h2 < length_0 ? _GEN_762 : _GEN_602; // @[executor.scala 308:60]
  wire [7:0] _GEN_923 = 8'h2 < length_0 ? _GEN_763 : _GEN_603; // @[executor.scala 308:60]
  wire [7:0] _GEN_924 = 8'h2 < length_0 ? _GEN_764 : _GEN_604; // @[executor.scala 308:60]
  wire [7:0] _GEN_925 = 8'h2 < length_0 ? _GEN_765 : _GEN_605; // @[executor.scala 308:60]
  wire [7:0] _GEN_926 = 8'h2 < length_0 ? _GEN_766 : _GEN_606; // @[executor.scala 308:60]
  wire [7:0] _GEN_927 = 8'h2 < length_0 ? _GEN_767 : _GEN_607; // @[executor.scala 308:60]
  wire [7:0] _GEN_928 = 8'h2 < length_0 ? _GEN_768 : _GEN_608; // @[executor.scala 308:60]
  wire [7:0] _GEN_929 = 8'h2 < length_0 ? _GEN_769 : _GEN_609; // @[executor.scala 308:60]
  wire [7:0] _GEN_930 = 8'h2 < length_0 ? _GEN_770 : _GEN_610; // @[executor.scala 308:60]
  wire [7:0] _GEN_931 = 8'h2 < length_0 ? _GEN_771 : _GEN_611; // @[executor.scala 308:60]
  wire [7:0] _GEN_932 = 8'h2 < length_0 ? _GEN_772 : _GEN_612; // @[executor.scala 308:60]
  wire [7:0] _GEN_933 = 8'h2 < length_0 ? _GEN_773 : _GEN_613; // @[executor.scala 308:60]
  wire [7:0] _GEN_934 = 8'h2 < length_0 ? _GEN_774 : _GEN_614; // @[executor.scala 308:60]
  wire [7:0] _GEN_935 = 8'h2 < length_0 ? _GEN_775 : _GEN_615; // @[executor.scala 308:60]
  wire [7:0] _GEN_936 = 8'h2 < length_0 ? _GEN_776 : _GEN_616; // @[executor.scala 308:60]
  wire [7:0] _GEN_937 = 8'h2 < length_0 ? _GEN_777 : _GEN_617; // @[executor.scala 308:60]
  wire [7:0] _GEN_938 = 8'h2 < length_0 ? _GEN_778 : _GEN_618; // @[executor.scala 308:60]
  wire [7:0] _GEN_939 = 8'h2 < length_0 ? _GEN_779 : _GEN_619; // @[executor.scala 308:60]
  wire [7:0] _GEN_940 = 8'h2 < length_0 ? _GEN_780 : _GEN_620; // @[executor.scala 308:60]
  wire [7:0] _GEN_941 = 8'h2 < length_0 ? _GEN_781 : _GEN_621; // @[executor.scala 308:60]
  wire [7:0] _GEN_942 = 8'h2 < length_0 ? _GEN_782 : _GEN_622; // @[executor.scala 308:60]
  wire [7:0] _GEN_943 = 8'h2 < length_0 ? _GEN_783 : _GEN_623; // @[executor.scala 308:60]
  wire [7:0] _GEN_944 = 8'h2 < length_0 ? _GEN_784 : _GEN_624; // @[executor.scala 308:60]
  wire [7:0] _GEN_945 = 8'h2 < length_0 ? _GEN_785 : _GEN_625; // @[executor.scala 308:60]
  wire [7:0] _GEN_946 = 8'h2 < length_0 ? _GEN_786 : _GEN_626; // @[executor.scala 308:60]
  wire [7:0] _GEN_947 = 8'h2 < length_0 ? _GEN_787 : _GEN_627; // @[executor.scala 308:60]
  wire [7:0] _GEN_948 = 8'h2 < length_0 ? _GEN_788 : _GEN_628; // @[executor.scala 308:60]
  wire [7:0] _GEN_949 = 8'h2 < length_0 ? _GEN_789 : _GEN_629; // @[executor.scala 308:60]
  wire [7:0] _GEN_950 = 8'h2 < length_0 ? _GEN_790 : _GEN_630; // @[executor.scala 308:60]
  wire [7:0] _GEN_951 = 8'h2 < length_0 ? _GEN_791 : _GEN_631; // @[executor.scala 308:60]
  wire [7:0] _GEN_952 = 8'h2 < length_0 ? _GEN_792 : _GEN_632; // @[executor.scala 308:60]
  wire [7:0] _GEN_953 = 8'h2 < length_0 ? _GEN_793 : _GEN_633; // @[executor.scala 308:60]
  wire [7:0] _GEN_954 = 8'h2 < length_0 ? _GEN_794 : _GEN_634; // @[executor.scala 308:60]
  wire [7:0] _GEN_955 = 8'h2 < length_0 ? _GEN_795 : _GEN_635; // @[executor.scala 308:60]
  wire [7:0] _GEN_956 = 8'h2 < length_0 ? _GEN_796 : _GEN_636; // @[executor.scala 308:60]
  wire [7:0] _GEN_957 = 8'h2 < length_0 ? _GEN_797 : _GEN_637; // @[executor.scala 308:60]
  wire [7:0] _GEN_958 = 8'h2 < length_0 ? _GEN_798 : _GEN_638; // @[executor.scala 308:60]
  wire [7:0] _GEN_959 = 8'h2 < length_0 ? _GEN_799 : _GEN_639; // @[executor.scala 308:60]
  wire [7:0] field_byte_3 = field_0[39:32]; // @[executor.scala 305:57]
  wire [7:0] total_offset_3 = offset_0 + 8'h3; // @[executor.scala 307:57]
  wire [7:0] _GEN_960 = 8'h0 == total_offset_3 ? field_byte_3 : _GEN_800; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_961 = 8'h1 == total_offset_3 ? field_byte_3 : _GEN_801; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_962 = 8'h2 == total_offset_3 ? field_byte_3 : _GEN_802; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_963 = 8'h3 == total_offset_3 ? field_byte_3 : _GEN_803; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_964 = 8'h4 == total_offset_3 ? field_byte_3 : _GEN_804; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_965 = 8'h5 == total_offset_3 ? field_byte_3 : _GEN_805; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_966 = 8'h6 == total_offset_3 ? field_byte_3 : _GEN_806; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_967 = 8'h7 == total_offset_3 ? field_byte_3 : _GEN_807; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_968 = 8'h8 == total_offset_3 ? field_byte_3 : _GEN_808; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_969 = 8'h9 == total_offset_3 ? field_byte_3 : _GEN_809; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_970 = 8'ha == total_offset_3 ? field_byte_3 : _GEN_810; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_971 = 8'hb == total_offset_3 ? field_byte_3 : _GEN_811; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_972 = 8'hc == total_offset_3 ? field_byte_3 : _GEN_812; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_973 = 8'hd == total_offset_3 ? field_byte_3 : _GEN_813; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_974 = 8'he == total_offset_3 ? field_byte_3 : _GEN_814; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_975 = 8'hf == total_offset_3 ? field_byte_3 : _GEN_815; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_976 = 8'h10 == total_offset_3 ? field_byte_3 : _GEN_816; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_977 = 8'h11 == total_offset_3 ? field_byte_3 : _GEN_817; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_978 = 8'h12 == total_offset_3 ? field_byte_3 : _GEN_818; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_979 = 8'h13 == total_offset_3 ? field_byte_3 : _GEN_819; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_980 = 8'h14 == total_offset_3 ? field_byte_3 : _GEN_820; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_981 = 8'h15 == total_offset_3 ? field_byte_3 : _GEN_821; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_982 = 8'h16 == total_offset_3 ? field_byte_3 : _GEN_822; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_983 = 8'h17 == total_offset_3 ? field_byte_3 : _GEN_823; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_984 = 8'h18 == total_offset_3 ? field_byte_3 : _GEN_824; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_985 = 8'h19 == total_offset_3 ? field_byte_3 : _GEN_825; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_986 = 8'h1a == total_offset_3 ? field_byte_3 : _GEN_826; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_987 = 8'h1b == total_offset_3 ? field_byte_3 : _GEN_827; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_988 = 8'h1c == total_offset_3 ? field_byte_3 : _GEN_828; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_989 = 8'h1d == total_offset_3 ? field_byte_3 : _GEN_829; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_990 = 8'h1e == total_offset_3 ? field_byte_3 : _GEN_830; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_991 = 8'h1f == total_offset_3 ? field_byte_3 : _GEN_831; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_992 = 8'h20 == total_offset_3 ? field_byte_3 : _GEN_832; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_993 = 8'h21 == total_offset_3 ? field_byte_3 : _GEN_833; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_994 = 8'h22 == total_offset_3 ? field_byte_3 : _GEN_834; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_995 = 8'h23 == total_offset_3 ? field_byte_3 : _GEN_835; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_996 = 8'h24 == total_offset_3 ? field_byte_3 : _GEN_836; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_997 = 8'h25 == total_offset_3 ? field_byte_3 : _GEN_837; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_998 = 8'h26 == total_offset_3 ? field_byte_3 : _GEN_838; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_999 = 8'h27 == total_offset_3 ? field_byte_3 : _GEN_839; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1000 = 8'h28 == total_offset_3 ? field_byte_3 : _GEN_840; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1001 = 8'h29 == total_offset_3 ? field_byte_3 : _GEN_841; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1002 = 8'h2a == total_offset_3 ? field_byte_3 : _GEN_842; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1003 = 8'h2b == total_offset_3 ? field_byte_3 : _GEN_843; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1004 = 8'h2c == total_offset_3 ? field_byte_3 : _GEN_844; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1005 = 8'h2d == total_offset_3 ? field_byte_3 : _GEN_845; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1006 = 8'h2e == total_offset_3 ? field_byte_3 : _GEN_846; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1007 = 8'h2f == total_offset_3 ? field_byte_3 : _GEN_847; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1008 = 8'h30 == total_offset_3 ? field_byte_3 : _GEN_848; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1009 = 8'h31 == total_offset_3 ? field_byte_3 : _GEN_849; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1010 = 8'h32 == total_offset_3 ? field_byte_3 : _GEN_850; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1011 = 8'h33 == total_offset_3 ? field_byte_3 : _GEN_851; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1012 = 8'h34 == total_offset_3 ? field_byte_3 : _GEN_852; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1013 = 8'h35 == total_offset_3 ? field_byte_3 : _GEN_853; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1014 = 8'h36 == total_offset_3 ? field_byte_3 : _GEN_854; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1015 = 8'h37 == total_offset_3 ? field_byte_3 : _GEN_855; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1016 = 8'h38 == total_offset_3 ? field_byte_3 : _GEN_856; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1017 = 8'h39 == total_offset_3 ? field_byte_3 : _GEN_857; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1018 = 8'h3a == total_offset_3 ? field_byte_3 : _GEN_858; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1019 = 8'h3b == total_offset_3 ? field_byte_3 : _GEN_859; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1020 = 8'h3c == total_offset_3 ? field_byte_3 : _GEN_860; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1021 = 8'h3d == total_offset_3 ? field_byte_3 : _GEN_861; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1022 = 8'h3e == total_offset_3 ? field_byte_3 : _GEN_862; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1023 = 8'h3f == total_offset_3 ? field_byte_3 : _GEN_863; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1024 = 8'h40 == total_offset_3 ? field_byte_3 : _GEN_864; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1025 = 8'h41 == total_offset_3 ? field_byte_3 : _GEN_865; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1026 = 8'h42 == total_offset_3 ? field_byte_3 : _GEN_866; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1027 = 8'h43 == total_offset_3 ? field_byte_3 : _GEN_867; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1028 = 8'h44 == total_offset_3 ? field_byte_3 : _GEN_868; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1029 = 8'h45 == total_offset_3 ? field_byte_3 : _GEN_869; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1030 = 8'h46 == total_offset_3 ? field_byte_3 : _GEN_870; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1031 = 8'h47 == total_offset_3 ? field_byte_3 : _GEN_871; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1032 = 8'h48 == total_offset_3 ? field_byte_3 : _GEN_872; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1033 = 8'h49 == total_offset_3 ? field_byte_3 : _GEN_873; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1034 = 8'h4a == total_offset_3 ? field_byte_3 : _GEN_874; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1035 = 8'h4b == total_offset_3 ? field_byte_3 : _GEN_875; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1036 = 8'h4c == total_offset_3 ? field_byte_3 : _GEN_876; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1037 = 8'h4d == total_offset_3 ? field_byte_3 : _GEN_877; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1038 = 8'h4e == total_offset_3 ? field_byte_3 : _GEN_878; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1039 = 8'h4f == total_offset_3 ? field_byte_3 : _GEN_879; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1040 = 8'h50 == total_offset_3 ? field_byte_3 : _GEN_880; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1041 = 8'h51 == total_offset_3 ? field_byte_3 : _GEN_881; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1042 = 8'h52 == total_offset_3 ? field_byte_3 : _GEN_882; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1043 = 8'h53 == total_offset_3 ? field_byte_3 : _GEN_883; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1044 = 8'h54 == total_offset_3 ? field_byte_3 : _GEN_884; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1045 = 8'h55 == total_offset_3 ? field_byte_3 : _GEN_885; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1046 = 8'h56 == total_offset_3 ? field_byte_3 : _GEN_886; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1047 = 8'h57 == total_offset_3 ? field_byte_3 : _GEN_887; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1048 = 8'h58 == total_offset_3 ? field_byte_3 : _GEN_888; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1049 = 8'h59 == total_offset_3 ? field_byte_3 : _GEN_889; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1050 = 8'h5a == total_offset_3 ? field_byte_3 : _GEN_890; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1051 = 8'h5b == total_offset_3 ? field_byte_3 : _GEN_891; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1052 = 8'h5c == total_offset_3 ? field_byte_3 : _GEN_892; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1053 = 8'h5d == total_offset_3 ? field_byte_3 : _GEN_893; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1054 = 8'h5e == total_offset_3 ? field_byte_3 : _GEN_894; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1055 = 8'h5f == total_offset_3 ? field_byte_3 : _GEN_895; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1056 = 8'h60 == total_offset_3 ? field_byte_3 : _GEN_896; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1057 = 8'h61 == total_offset_3 ? field_byte_3 : _GEN_897; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1058 = 8'h62 == total_offset_3 ? field_byte_3 : _GEN_898; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1059 = 8'h63 == total_offset_3 ? field_byte_3 : _GEN_899; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1060 = 8'h64 == total_offset_3 ? field_byte_3 : _GEN_900; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1061 = 8'h65 == total_offset_3 ? field_byte_3 : _GEN_901; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1062 = 8'h66 == total_offset_3 ? field_byte_3 : _GEN_902; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1063 = 8'h67 == total_offset_3 ? field_byte_3 : _GEN_903; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1064 = 8'h68 == total_offset_3 ? field_byte_3 : _GEN_904; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1065 = 8'h69 == total_offset_3 ? field_byte_3 : _GEN_905; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1066 = 8'h6a == total_offset_3 ? field_byte_3 : _GEN_906; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1067 = 8'h6b == total_offset_3 ? field_byte_3 : _GEN_907; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1068 = 8'h6c == total_offset_3 ? field_byte_3 : _GEN_908; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1069 = 8'h6d == total_offset_3 ? field_byte_3 : _GEN_909; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1070 = 8'h6e == total_offset_3 ? field_byte_3 : _GEN_910; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1071 = 8'h6f == total_offset_3 ? field_byte_3 : _GEN_911; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1072 = 8'h70 == total_offset_3 ? field_byte_3 : _GEN_912; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1073 = 8'h71 == total_offset_3 ? field_byte_3 : _GEN_913; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1074 = 8'h72 == total_offset_3 ? field_byte_3 : _GEN_914; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1075 = 8'h73 == total_offset_3 ? field_byte_3 : _GEN_915; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1076 = 8'h74 == total_offset_3 ? field_byte_3 : _GEN_916; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1077 = 8'h75 == total_offset_3 ? field_byte_3 : _GEN_917; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1078 = 8'h76 == total_offset_3 ? field_byte_3 : _GEN_918; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1079 = 8'h77 == total_offset_3 ? field_byte_3 : _GEN_919; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1080 = 8'h78 == total_offset_3 ? field_byte_3 : _GEN_920; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1081 = 8'h79 == total_offset_3 ? field_byte_3 : _GEN_921; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1082 = 8'h7a == total_offset_3 ? field_byte_3 : _GEN_922; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1083 = 8'h7b == total_offset_3 ? field_byte_3 : _GEN_923; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1084 = 8'h7c == total_offset_3 ? field_byte_3 : _GEN_924; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1085 = 8'h7d == total_offset_3 ? field_byte_3 : _GEN_925; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1086 = 8'h7e == total_offset_3 ? field_byte_3 : _GEN_926; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1087 = 8'h7f == total_offset_3 ? field_byte_3 : _GEN_927; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1088 = 8'h80 == total_offset_3 ? field_byte_3 : _GEN_928; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1089 = 8'h81 == total_offset_3 ? field_byte_3 : _GEN_929; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1090 = 8'h82 == total_offset_3 ? field_byte_3 : _GEN_930; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1091 = 8'h83 == total_offset_3 ? field_byte_3 : _GEN_931; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1092 = 8'h84 == total_offset_3 ? field_byte_3 : _GEN_932; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1093 = 8'h85 == total_offset_3 ? field_byte_3 : _GEN_933; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1094 = 8'h86 == total_offset_3 ? field_byte_3 : _GEN_934; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1095 = 8'h87 == total_offset_3 ? field_byte_3 : _GEN_935; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1096 = 8'h88 == total_offset_3 ? field_byte_3 : _GEN_936; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1097 = 8'h89 == total_offset_3 ? field_byte_3 : _GEN_937; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1098 = 8'h8a == total_offset_3 ? field_byte_3 : _GEN_938; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1099 = 8'h8b == total_offset_3 ? field_byte_3 : _GEN_939; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1100 = 8'h8c == total_offset_3 ? field_byte_3 : _GEN_940; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1101 = 8'h8d == total_offset_3 ? field_byte_3 : _GEN_941; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1102 = 8'h8e == total_offset_3 ? field_byte_3 : _GEN_942; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1103 = 8'h8f == total_offset_3 ? field_byte_3 : _GEN_943; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1104 = 8'h90 == total_offset_3 ? field_byte_3 : _GEN_944; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1105 = 8'h91 == total_offset_3 ? field_byte_3 : _GEN_945; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1106 = 8'h92 == total_offset_3 ? field_byte_3 : _GEN_946; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1107 = 8'h93 == total_offset_3 ? field_byte_3 : _GEN_947; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1108 = 8'h94 == total_offset_3 ? field_byte_3 : _GEN_948; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1109 = 8'h95 == total_offset_3 ? field_byte_3 : _GEN_949; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1110 = 8'h96 == total_offset_3 ? field_byte_3 : _GEN_950; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1111 = 8'h97 == total_offset_3 ? field_byte_3 : _GEN_951; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1112 = 8'h98 == total_offset_3 ? field_byte_3 : _GEN_952; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1113 = 8'h99 == total_offset_3 ? field_byte_3 : _GEN_953; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1114 = 8'h9a == total_offset_3 ? field_byte_3 : _GEN_954; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1115 = 8'h9b == total_offset_3 ? field_byte_3 : _GEN_955; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1116 = 8'h9c == total_offset_3 ? field_byte_3 : _GEN_956; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1117 = 8'h9d == total_offset_3 ? field_byte_3 : _GEN_957; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1118 = 8'h9e == total_offset_3 ? field_byte_3 : _GEN_958; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1119 = 8'h9f == total_offset_3 ? field_byte_3 : _GEN_959; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1120 = 8'h3 < length_0 ? _GEN_960 : _GEN_800; // @[executor.scala 308:60]
  wire [7:0] _GEN_1121 = 8'h3 < length_0 ? _GEN_961 : _GEN_801; // @[executor.scala 308:60]
  wire [7:0] _GEN_1122 = 8'h3 < length_0 ? _GEN_962 : _GEN_802; // @[executor.scala 308:60]
  wire [7:0] _GEN_1123 = 8'h3 < length_0 ? _GEN_963 : _GEN_803; // @[executor.scala 308:60]
  wire [7:0] _GEN_1124 = 8'h3 < length_0 ? _GEN_964 : _GEN_804; // @[executor.scala 308:60]
  wire [7:0] _GEN_1125 = 8'h3 < length_0 ? _GEN_965 : _GEN_805; // @[executor.scala 308:60]
  wire [7:0] _GEN_1126 = 8'h3 < length_0 ? _GEN_966 : _GEN_806; // @[executor.scala 308:60]
  wire [7:0] _GEN_1127 = 8'h3 < length_0 ? _GEN_967 : _GEN_807; // @[executor.scala 308:60]
  wire [7:0] _GEN_1128 = 8'h3 < length_0 ? _GEN_968 : _GEN_808; // @[executor.scala 308:60]
  wire [7:0] _GEN_1129 = 8'h3 < length_0 ? _GEN_969 : _GEN_809; // @[executor.scala 308:60]
  wire [7:0] _GEN_1130 = 8'h3 < length_0 ? _GEN_970 : _GEN_810; // @[executor.scala 308:60]
  wire [7:0] _GEN_1131 = 8'h3 < length_0 ? _GEN_971 : _GEN_811; // @[executor.scala 308:60]
  wire [7:0] _GEN_1132 = 8'h3 < length_0 ? _GEN_972 : _GEN_812; // @[executor.scala 308:60]
  wire [7:0] _GEN_1133 = 8'h3 < length_0 ? _GEN_973 : _GEN_813; // @[executor.scala 308:60]
  wire [7:0] _GEN_1134 = 8'h3 < length_0 ? _GEN_974 : _GEN_814; // @[executor.scala 308:60]
  wire [7:0] _GEN_1135 = 8'h3 < length_0 ? _GEN_975 : _GEN_815; // @[executor.scala 308:60]
  wire [7:0] _GEN_1136 = 8'h3 < length_0 ? _GEN_976 : _GEN_816; // @[executor.scala 308:60]
  wire [7:0] _GEN_1137 = 8'h3 < length_0 ? _GEN_977 : _GEN_817; // @[executor.scala 308:60]
  wire [7:0] _GEN_1138 = 8'h3 < length_0 ? _GEN_978 : _GEN_818; // @[executor.scala 308:60]
  wire [7:0] _GEN_1139 = 8'h3 < length_0 ? _GEN_979 : _GEN_819; // @[executor.scala 308:60]
  wire [7:0] _GEN_1140 = 8'h3 < length_0 ? _GEN_980 : _GEN_820; // @[executor.scala 308:60]
  wire [7:0] _GEN_1141 = 8'h3 < length_0 ? _GEN_981 : _GEN_821; // @[executor.scala 308:60]
  wire [7:0] _GEN_1142 = 8'h3 < length_0 ? _GEN_982 : _GEN_822; // @[executor.scala 308:60]
  wire [7:0] _GEN_1143 = 8'h3 < length_0 ? _GEN_983 : _GEN_823; // @[executor.scala 308:60]
  wire [7:0] _GEN_1144 = 8'h3 < length_0 ? _GEN_984 : _GEN_824; // @[executor.scala 308:60]
  wire [7:0] _GEN_1145 = 8'h3 < length_0 ? _GEN_985 : _GEN_825; // @[executor.scala 308:60]
  wire [7:0] _GEN_1146 = 8'h3 < length_0 ? _GEN_986 : _GEN_826; // @[executor.scala 308:60]
  wire [7:0] _GEN_1147 = 8'h3 < length_0 ? _GEN_987 : _GEN_827; // @[executor.scala 308:60]
  wire [7:0] _GEN_1148 = 8'h3 < length_0 ? _GEN_988 : _GEN_828; // @[executor.scala 308:60]
  wire [7:0] _GEN_1149 = 8'h3 < length_0 ? _GEN_989 : _GEN_829; // @[executor.scala 308:60]
  wire [7:0] _GEN_1150 = 8'h3 < length_0 ? _GEN_990 : _GEN_830; // @[executor.scala 308:60]
  wire [7:0] _GEN_1151 = 8'h3 < length_0 ? _GEN_991 : _GEN_831; // @[executor.scala 308:60]
  wire [7:0] _GEN_1152 = 8'h3 < length_0 ? _GEN_992 : _GEN_832; // @[executor.scala 308:60]
  wire [7:0] _GEN_1153 = 8'h3 < length_0 ? _GEN_993 : _GEN_833; // @[executor.scala 308:60]
  wire [7:0] _GEN_1154 = 8'h3 < length_0 ? _GEN_994 : _GEN_834; // @[executor.scala 308:60]
  wire [7:0] _GEN_1155 = 8'h3 < length_0 ? _GEN_995 : _GEN_835; // @[executor.scala 308:60]
  wire [7:0] _GEN_1156 = 8'h3 < length_0 ? _GEN_996 : _GEN_836; // @[executor.scala 308:60]
  wire [7:0] _GEN_1157 = 8'h3 < length_0 ? _GEN_997 : _GEN_837; // @[executor.scala 308:60]
  wire [7:0] _GEN_1158 = 8'h3 < length_0 ? _GEN_998 : _GEN_838; // @[executor.scala 308:60]
  wire [7:0] _GEN_1159 = 8'h3 < length_0 ? _GEN_999 : _GEN_839; // @[executor.scala 308:60]
  wire [7:0] _GEN_1160 = 8'h3 < length_0 ? _GEN_1000 : _GEN_840; // @[executor.scala 308:60]
  wire [7:0] _GEN_1161 = 8'h3 < length_0 ? _GEN_1001 : _GEN_841; // @[executor.scala 308:60]
  wire [7:0] _GEN_1162 = 8'h3 < length_0 ? _GEN_1002 : _GEN_842; // @[executor.scala 308:60]
  wire [7:0] _GEN_1163 = 8'h3 < length_0 ? _GEN_1003 : _GEN_843; // @[executor.scala 308:60]
  wire [7:0] _GEN_1164 = 8'h3 < length_0 ? _GEN_1004 : _GEN_844; // @[executor.scala 308:60]
  wire [7:0] _GEN_1165 = 8'h3 < length_0 ? _GEN_1005 : _GEN_845; // @[executor.scala 308:60]
  wire [7:0] _GEN_1166 = 8'h3 < length_0 ? _GEN_1006 : _GEN_846; // @[executor.scala 308:60]
  wire [7:0] _GEN_1167 = 8'h3 < length_0 ? _GEN_1007 : _GEN_847; // @[executor.scala 308:60]
  wire [7:0] _GEN_1168 = 8'h3 < length_0 ? _GEN_1008 : _GEN_848; // @[executor.scala 308:60]
  wire [7:0] _GEN_1169 = 8'h3 < length_0 ? _GEN_1009 : _GEN_849; // @[executor.scala 308:60]
  wire [7:0] _GEN_1170 = 8'h3 < length_0 ? _GEN_1010 : _GEN_850; // @[executor.scala 308:60]
  wire [7:0] _GEN_1171 = 8'h3 < length_0 ? _GEN_1011 : _GEN_851; // @[executor.scala 308:60]
  wire [7:0] _GEN_1172 = 8'h3 < length_0 ? _GEN_1012 : _GEN_852; // @[executor.scala 308:60]
  wire [7:0] _GEN_1173 = 8'h3 < length_0 ? _GEN_1013 : _GEN_853; // @[executor.scala 308:60]
  wire [7:0] _GEN_1174 = 8'h3 < length_0 ? _GEN_1014 : _GEN_854; // @[executor.scala 308:60]
  wire [7:0] _GEN_1175 = 8'h3 < length_0 ? _GEN_1015 : _GEN_855; // @[executor.scala 308:60]
  wire [7:0] _GEN_1176 = 8'h3 < length_0 ? _GEN_1016 : _GEN_856; // @[executor.scala 308:60]
  wire [7:0] _GEN_1177 = 8'h3 < length_0 ? _GEN_1017 : _GEN_857; // @[executor.scala 308:60]
  wire [7:0] _GEN_1178 = 8'h3 < length_0 ? _GEN_1018 : _GEN_858; // @[executor.scala 308:60]
  wire [7:0] _GEN_1179 = 8'h3 < length_0 ? _GEN_1019 : _GEN_859; // @[executor.scala 308:60]
  wire [7:0] _GEN_1180 = 8'h3 < length_0 ? _GEN_1020 : _GEN_860; // @[executor.scala 308:60]
  wire [7:0] _GEN_1181 = 8'h3 < length_0 ? _GEN_1021 : _GEN_861; // @[executor.scala 308:60]
  wire [7:0] _GEN_1182 = 8'h3 < length_0 ? _GEN_1022 : _GEN_862; // @[executor.scala 308:60]
  wire [7:0] _GEN_1183 = 8'h3 < length_0 ? _GEN_1023 : _GEN_863; // @[executor.scala 308:60]
  wire [7:0] _GEN_1184 = 8'h3 < length_0 ? _GEN_1024 : _GEN_864; // @[executor.scala 308:60]
  wire [7:0] _GEN_1185 = 8'h3 < length_0 ? _GEN_1025 : _GEN_865; // @[executor.scala 308:60]
  wire [7:0] _GEN_1186 = 8'h3 < length_0 ? _GEN_1026 : _GEN_866; // @[executor.scala 308:60]
  wire [7:0] _GEN_1187 = 8'h3 < length_0 ? _GEN_1027 : _GEN_867; // @[executor.scala 308:60]
  wire [7:0] _GEN_1188 = 8'h3 < length_0 ? _GEN_1028 : _GEN_868; // @[executor.scala 308:60]
  wire [7:0] _GEN_1189 = 8'h3 < length_0 ? _GEN_1029 : _GEN_869; // @[executor.scala 308:60]
  wire [7:0] _GEN_1190 = 8'h3 < length_0 ? _GEN_1030 : _GEN_870; // @[executor.scala 308:60]
  wire [7:0] _GEN_1191 = 8'h3 < length_0 ? _GEN_1031 : _GEN_871; // @[executor.scala 308:60]
  wire [7:0] _GEN_1192 = 8'h3 < length_0 ? _GEN_1032 : _GEN_872; // @[executor.scala 308:60]
  wire [7:0] _GEN_1193 = 8'h3 < length_0 ? _GEN_1033 : _GEN_873; // @[executor.scala 308:60]
  wire [7:0] _GEN_1194 = 8'h3 < length_0 ? _GEN_1034 : _GEN_874; // @[executor.scala 308:60]
  wire [7:0] _GEN_1195 = 8'h3 < length_0 ? _GEN_1035 : _GEN_875; // @[executor.scala 308:60]
  wire [7:0] _GEN_1196 = 8'h3 < length_0 ? _GEN_1036 : _GEN_876; // @[executor.scala 308:60]
  wire [7:0] _GEN_1197 = 8'h3 < length_0 ? _GEN_1037 : _GEN_877; // @[executor.scala 308:60]
  wire [7:0] _GEN_1198 = 8'h3 < length_0 ? _GEN_1038 : _GEN_878; // @[executor.scala 308:60]
  wire [7:0] _GEN_1199 = 8'h3 < length_0 ? _GEN_1039 : _GEN_879; // @[executor.scala 308:60]
  wire [7:0] _GEN_1200 = 8'h3 < length_0 ? _GEN_1040 : _GEN_880; // @[executor.scala 308:60]
  wire [7:0] _GEN_1201 = 8'h3 < length_0 ? _GEN_1041 : _GEN_881; // @[executor.scala 308:60]
  wire [7:0] _GEN_1202 = 8'h3 < length_0 ? _GEN_1042 : _GEN_882; // @[executor.scala 308:60]
  wire [7:0] _GEN_1203 = 8'h3 < length_0 ? _GEN_1043 : _GEN_883; // @[executor.scala 308:60]
  wire [7:0] _GEN_1204 = 8'h3 < length_0 ? _GEN_1044 : _GEN_884; // @[executor.scala 308:60]
  wire [7:0] _GEN_1205 = 8'h3 < length_0 ? _GEN_1045 : _GEN_885; // @[executor.scala 308:60]
  wire [7:0] _GEN_1206 = 8'h3 < length_0 ? _GEN_1046 : _GEN_886; // @[executor.scala 308:60]
  wire [7:0] _GEN_1207 = 8'h3 < length_0 ? _GEN_1047 : _GEN_887; // @[executor.scala 308:60]
  wire [7:0] _GEN_1208 = 8'h3 < length_0 ? _GEN_1048 : _GEN_888; // @[executor.scala 308:60]
  wire [7:0] _GEN_1209 = 8'h3 < length_0 ? _GEN_1049 : _GEN_889; // @[executor.scala 308:60]
  wire [7:0] _GEN_1210 = 8'h3 < length_0 ? _GEN_1050 : _GEN_890; // @[executor.scala 308:60]
  wire [7:0] _GEN_1211 = 8'h3 < length_0 ? _GEN_1051 : _GEN_891; // @[executor.scala 308:60]
  wire [7:0] _GEN_1212 = 8'h3 < length_0 ? _GEN_1052 : _GEN_892; // @[executor.scala 308:60]
  wire [7:0] _GEN_1213 = 8'h3 < length_0 ? _GEN_1053 : _GEN_893; // @[executor.scala 308:60]
  wire [7:0] _GEN_1214 = 8'h3 < length_0 ? _GEN_1054 : _GEN_894; // @[executor.scala 308:60]
  wire [7:0] _GEN_1215 = 8'h3 < length_0 ? _GEN_1055 : _GEN_895; // @[executor.scala 308:60]
  wire [7:0] _GEN_1216 = 8'h3 < length_0 ? _GEN_1056 : _GEN_896; // @[executor.scala 308:60]
  wire [7:0] _GEN_1217 = 8'h3 < length_0 ? _GEN_1057 : _GEN_897; // @[executor.scala 308:60]
  wire [7:0] _GEN_1218 = 8'h3 < length_0 ? _GEN_1058 : _GEN_898; // @[executor.scala 308:60]
  wire [7:0] _GEN_1219 = 8'h3 < length_0 ? _GEN_1059 : _GEN_899; // @[executor.scala 308:60]
  wire [7:0] _GEN_1220 = 8'h3 < length_0 ? _GEN_1060 : _GEN_900; // @[executor.scala 308:60]
  wire [7:0] _GEN_1221 = 8'h3 < length_0 ? _GEN_1061 : _GEN_901; // @[executor.scala 308:60]
  wire [7:0] _GEN_1222 = 8'h3 < length_0 ? _GEN_1062 : _GEN_902; // @[executor.scala 308:60]
  wire [7:0] _GEN_1223 = 8'h3 < length_0 ? _GEN_1063 : _GEN_903; // @[executor.scala 308:60]
  wire [7:0] _GEN_1224 = 8'h3 < length_0 ? _GEN_1064 : _GEN_904; // @[executor.scala 308:60]
  wire [7:0] _GEN_1225 = 8'h3 < length_0 ? _GEN_1065 : _GEN_905; // @[executor.scala 308:60]
  wire [7:0] _GEN_1226 = 8'h3 < length_0 ? _GEN_1066 : _GEN_906; // @[executor.scala 308:60]
  wire [7:0] _GEN_1227 = 8'h3 < length_0 ? _GEN_1067 : _GEN_907; // @[executor.scala 308:60]
  wire [7:0] _GEN_1228 = 8'h3 < length_0 ? _GEN_1068 : _GEN_908; // @[executor.scala 308:60]
  wire [7:0] _GEN_1229 = 8'h3 < length_0 ? _GEN_1069 : _GEN_909; // @[executor.scala 308:60]
  wire [7:0] _GEN_1230 = 8'h3 < length_0 ? _GEN_1070 : _GEN_910; // @[executor.scala 308:60]
  wire [7:0] _GEN_1231 = 8'h3 < length_0 ? _GEN_1071 : _GEN_911; // @[executor.scala 308:60]
  wire [7:0] _GEN_1232 = 8'h3 < length_0 ? _GEN_1072 : _GEN_912; // @[executor.scala 308:60]
  wire [7:0] _GEN_1233 = 8'h3 < length_0 ? _GEN_1073 : _GEN_913; // @[executor.scala 308:60]
  wire [7:0] _GEN_1234 = 8'h3 < length_0 ? _GEN_1074 : _GEN_914; // @[executor.scala 308:60]
  wire [7:0] _GEN_1235 = 8'h3 < length_0 ? _GEN_1075 : _GEN_915; // @[executor.scala 308:60]
  wire [7:0] _GEN_1236 = 8'h3 < length_0 ? _GEN_1076 : _GEN_916; // @[executor.scala 308:60]
  wire [7:0] _GEN_1237 = 8'h3 < length_0 ? _GEN_1077 : _GEN_917; // @[executor.scala 308:60]
  wire [7:0] _GEN_1238 = 8'h3 < length_0 ? _GEN_1078 : _GEN_918; // @[executor.scala 308:60]
  wire [7:0] _GEN_1239 = 8'h3 < length_0 ? _GEN_1079 : _GEN_919; // @[executor.scala 308:60]
  wire [7:0] _GEN_1240 = 8'h3 < length_0 ? _GEN_1080 : _GEN_920; // @[executor.scala 308:60]
  wire [7:0] _GEN_1241 = 8'h3 < length_0 ? _GEN_1081 : _GEN_921; // @[executor.scala 308:60]
  wire [7:0] _GEN_1242 = 8'h3 < length_0 ? _GEN_1082 : _GEN_922; // @[executor.scala 308:60]
  wire [7:0] _GEN_1243 = 8'h3 < length_0 ? _GEN_1083 : _GEN_923; // @[executor.scala 308:60]
  wire [7:0] _GEN_1244 = 8'h3 < length_0 ? _GEN_1084 : _GEN_924; // @[executor.scala 308:60]
  wire [7:0] _GEN_1245 = 8'h3 < length_0 ? _GEN_1085 : _GEN_925; // @[executor.scala 308:60]
  wire [7:0] _GEN_1246 = 8'h3 < length_0 ? _GEN_1086 : _GEN_926; // @[executor.scala 308:60]
  wire [7:0] _GEN_1247 = 8'h3 < length_0 ? _GEN_1087 : _GEN_927; // @[executor.scala 308:60]
  wire [7:0] _GEN_1248 = 8'h3 < length_0 ? _GEN_1088 : _GEN_928; // @[executor.scala 308:60]
  wire [7:0] _GEN_1249 = 8'h3 < length_0 ? _GEN_1089 : _GEN_929; // @[executor.scala 308:60]
  wire [7:0] _GEN_1250 = 8'h3 < length_0 ? _GEN_1090 : _GEN_930; // @[executor.scala 308:60]
  wire [7:0] _GEN_1251 = 8'h3 < length_0 ? _GEN_1091 : _GEN_931; // @[executor.scala 308:60]
  wire [7:0] _GEN_1252 = 8'h3 < length_0 ? _GEN_1092 : _GEN_932; // @[executor.scala 308:60]
  wire [7:0] _GEN_1253 = 8'h3 < length_0 ? _GEN_1093 : _GEN_933; // @[executor.scala 308:60]
  wire [7:0] _GEN_1254 = 8'h3 < length_0 ? _GEN_1094 : _GEN_934; // @[executor.scala 308:60]
  wire [7:0] _GEN_1255 = 8'h3 < length_0 ? _GEN_1095 : _GEN_935; // @[executor.scala 308:60]
  wire [7:0] _GEN_1256 = 8'h3 < length_0 ? _GEN_1096 : _GEN_936; // @[executor.scala 308:60]
  wire [7:0] _GEN_1257 = 8'h3 < length_0 ? _GEN_1097 : _GEN_937; // @[executor.scala 308:60]
  wire [7:0] _GEN_1258 = 8'h3 < length_0 ? _GEN_1098 : _GEN_938; // @[executor.scala 308:60]
  wire [7:0] _GEN_1259 = 8'h3 < length_0 ? _GEN_1099 : _GEN_939; // @[executor.scala 308:60]
  wire [7:0] _GEN_1260 = 8'h3 < length_0 ? _GEN_1100 : _GEN_940; // @[executor.scala 308:60]
  wire [7:0] _GEN_1261 = 8'h3 < length_0 ? _GEN_1101 : _GEN_941; // @[executor.scala 308:60]
  wire [7:0] _GEN_1262 = 8'h3 < length_0 ? _GEN_1102 : _GEN_942; // @[executor.scala 308:60]
  wire [7:0] _GEN_1263 = 8'h3 < length_0 ? _GEN_1103 : _GEN_943; // @[executor.scala 308:60]
  wire [7:0] _GEN_1264 = 8'h3 < length_0 ? _GEN_1104 : _GEN_944; // @[executor.scala 308:60]
  wire [7:0] _GEN_1265 = 8'h3 < length_0 ? _GEN_1105 : _GEN_945; // @[executor.scala 308:60]
  wire [7:0] _GEN_1266 = 8'h3 < length_0 ? _GEN_1106 : _GEN_946; // @[executor.scala 308:60]
  wire [7:0] _GEN_1267 = 8'h3 < length_0 ? _GEN_1107 : _GEN_947; // @[executor.scala 308:60]
  wire [7:0] _GEN_1268 = 8'h3 < length_0 ? _GEN_1108 : _GEN_948; // @[executor.scala 308:60]
  wire [7:0] _GEN_1269 = 8'h3 < length_0 ? _GEN_1109 : _GEN_949; // @[executor.scala 308:60]
  wire [7:0] _GEN_1270 = 8'h3 < length_0 ? _GEN_1110 : _GEN_950; // @[executor.scala 308:60]
  wire [7:0] _GEN_1271 = 8'h3 < length_0 ? _GEN_1111 : _GEN_951; // @[executor.scala 308:60]
  wire [7:0] _GEN_1272 = 8'h3 < length_0 ? _GEN_1112 : _GEN_952; // @[executor.scala 308:60]
  wire [7:0] _GEN_1273 = 8'h3 < length_0 ? _GEN_1113 : _GEN_953; // @[executor.scala 308:60]
  wire [7:0] _GEN_1274 = 8'h3 < length_0 ? _GEN_1114 : _GEN_954; // @[executor.scala 308:60]
  wire [7:0] _GEN_1275 = 8'h3 < length_0 ? _GEN_1115 : _GEN_955; // @[executor.scala 308:60]
  wire [7:0] _GEN_1276 = 8'h3 < length_0 ? _GEN_1116 : _GEN_956; // @[executor.scala 308:60]
  wire [7:0] _GEN_1277 = 8'h3 < length_0 ? _GEN_1117 : _GEN_957; // @[executor.scala 308:60]
  wire [7:0] _GEN_1278 = 8'h3 < length_0 ? _GEN_1118 : _GEN_958; // @[executor.scala 308:60]
  wire [7:0] _GEN_1279 = 8'h3 < length_0 ? _GEN_1119 : _GEN_959; // @[executor.scala 308:60]
  wire [7:0] field_byte_4 = field_0[31:24]; // @[executor.scala 305:57]
  wire [7:0] total_offset_4 = offset_0 + 8'h4; // @[executor.scala 307:57]
  wire [7:0] _GEN_1280 = 8'h0 == total_offset_4 ? field_byte_4 : _GEN_1120; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1281 = 8'h1 == total_offset_4 ? field_byte_4 : _GEN_1121; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1282 = 8'h2 == total_offset_4 ? field_byte_4 : _GEN_1122; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1283 = 8'h3 == total_offset_4 ? field_byte_4 : _GEN_1123; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1284 = 8'h4 == total_offset_4 ? field_byte_4 : _GEN_1124; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1285 = 8'h5 == total_offset_4 ? field_byte_4 : _GEN_1125; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1286 = 8'h6 == total_offset_4 ? field_byte_4 : _GEN_1126; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1287 = 8'h7 == total_offset_4 ? field_byte_4 : _GEN_1127; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1288 = 8'h8 == total_offset_4 ? field_byte_4 : _GEN_1128; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1289 = 8'h9 == total_offset_4 ? field_byte_4 : _GEN_1129; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1290 = 8'ha == total_offset_4 ? field_byte_4 : _GEN_1130; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1291 = 8'hb == total_offset_4 ? field_byte_4 : _GEN_1131; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1292 = 8'hc == total_offset_4 ? field_byte_4 : _GEN_1132; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1293 = 8'hd == total_offset_4 ? field_byte_4 : _GEN_1133; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1294 = 8'he == total_offset_4 ? field_byte_4 : _GEN_1134; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1295 = 8'hf == total_offset_4 ? field_byte_4 : _GEN_1135; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1296 = 8'h10 == total_offset_4 ? field_byte_4 : _GEN_1136; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1297 = 8'h11 == total_offset_4 ? field_byte_4 : _GEN_1137; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1298 = 8'h12 == total_offset_4 ? field_byte_4 : _GEN_1138; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1299 = 8'h13 == total_offset_4 ? field_byte_4 : _GEN_1139; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1300 = 8'h14 == total_offset_4 ? field_byte_4 : _GEN_1140; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1301 = 8'h15 == total_offset_4 ? field_byte_4 : _GEN_1141; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1302 = 8'h16 == total_offset_4 ? field_byte_4 : _GEN_1142; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1303 = 8'h17 == total_offset_4 ? field_byte_4 : _GEN_1143; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1304 = 8'h18 == total_offset_4 ? field_byte_4 : _GEN_1144; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1305 = 8'h19 == total_offset_4 ? field_byte_4 : _GEN_1145; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1306 = 8'h1a == total_offset_4 ? field_byte_4 : _GEN_1146; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1307 = 8'h1b == total_offset_4 ? field_byte_4 : _GEN_1147; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1308 = 8'h1c == total_offset_4 ? field_byte_4 : _GEN_1148; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1309 = 8'h1d == total_offset_4 ? field_byte_4 : _GEN_1149; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1310 = 8'h1e == total_offset_4 ? field_byte_4 : _GEN_1150; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1311 = 8'h1f == total_offset_4 ? field_byte_4 : _GEN_1151; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1312 = 8'h20 == total_offset_4 ? field_byte_4 : _GEN_1152; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1313 = 8'h21 == total_offset_4 ? field_byte_4 : _GEN_1153; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1314 = 8'h22 == total_offset_4 ? field_byte_4 : _GEN_1154; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1315 = 8'h23 == total_offset_4 ? field_byte_4 : _GEN_1155; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1316 = 8'h24 == total_offset_4 ? field_byte_4 : _GEN_1156; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1317 = 8'h25 == total_offset_4 ? field_byte_4 : _GEN_1157; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1318 = 8'h26 == total_offset_4 ? field_byte_4 : _GEN_1158; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1319 = 8'h27 == total_offset_4 ? field_byte_4 : _GEN_1159; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1320 = 8'h28 == total_offset_4 ? field_byte_4 : _GEN_1160; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1321 = 8'h29 == total_offset_4 ? field_byte_4 : _GEN_1161; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1322 = 8'h2a == total_offset_4 ? field_byte_4 : _GEN_1162; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1323 = 8'h2b == total_offset_4 ? field_byte_4 : _GEN_1163; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1324 = 8'h2c == total_offset_4 ? field_byte_4 : _GEN_1164; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1325 = 8'h2d == total_offset_4 ? field_byte_4 : _GEN_1165; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1326 = 8'h2e == total_offset_4 ? field_byte_4 : _GEN_1166; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1327 = 8'h2f == total_offset_4 ? field_byte_4 : _GEN_1167; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1328 = 8'h30 == total_offset_4 ? field_byte_4 : _GEN_1168; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1329 = 8'h31 == total_offset_4 ? field_byte_4 : _GEN_1169; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1330 = 8'h32 == total_offset_4 ? field_byte_4 : _GEN_1170; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1331 = 8'h33 == total_offset_4 ? field_byte_4 : _GEN_1171; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1332 = 8'h34 == total_offset_4 ? field_byte_4 : _GEN_1172; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1333 = 8'h35 == total_offset_4 ? field_byte_4 : _GEN_1173; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1334 = 8'h36 == total_offset_4 ? field_byte_4 : _GEN_1174; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1335 = 8'h37 == total_offset_4 ? field_byte_4 : _GEN_1175; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1336 = 8'h38 == total_offset_4 ? field_byte_4 : _GEN_1176; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1337 = 8'h39 == total_offset_4 ? field_byte_4 : _GEN_1177; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1338 = 8'h3a == total_offset_4 ? field_byte_4 : _GEN_1178; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1339 = 8'h3b == total_offset_4 ? field_byte_4 : _GEN_1179; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1340 = 8'h3c == total_offset_4 ? field_byte_4 : _GEN_1180; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1341 = 8'h3d == total_offset_4 ? field_byte_4 : _GEN_1181; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1342 = 8'h3e == total_offset_4 ? field_byte_4 : _GEN_1182; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1343 = 8'h3f == total_offset_4 ? field_byte_4 : _GEN_1183; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1344 = 8'h40 == total_offset_4 ? field_byte_4 : _GEN_1184; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1345 = 8'h41 == total_offset_4 ? field_byte_4 : _GEN_1185; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1346 = 8'h42 == total_offset_4 ? field_byte_4 : _GEN_1186; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1347 = 8'h43 == total_offset_4 ? field_byte_4 : _GEN_1187; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1348 = 8'h44 == total_offset_4 ? field_byte_4 : _GEN_1188; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1349 = 8'h45 == total_offset_4 ? field_byte_4 : _GEN_1189; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1350 = 8'h46 == total_offset_4 ? field_byte_4 : _GEN_1190; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1351 = 8'h47 == total_offset_4 ? field_byte_4 : _GEN_1191; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1352 = 8'h48 == total_offset_4 ? field_byte_4 : _GEN_1192; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1353 = 8'h49 == total_offset_4 ? field_byte_4 : _GEN_1193; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1354 = 8'h4a == total_offset_4 ? field_byte_4 : _GEN_1194; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1355 = 8'h4b == total_offset_4 ? field_byte_4 : _GEN_1195; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1356 = 8'h4c == total_offset_4 ? field_byte_4 : _GEN_1196; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1357 = 8'h4d == total_offset_4 ? field_byte_4 : _GEN_1197; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1358 = 8'h4e == total_offset_4 ? field_byte_4 : _GEN_1198; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1359 = 8'h4f == total_offset_4 ? field_byte_4 : _GEN_1199; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1360 = 8'h50 == total_offset_4 ? field_byte_4 : _GEN_1200; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1361 = 8'h51 == total_offset_4 ? field_byte_4 : _GEN_1201; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1362 = 8'h52 == total_offset_4 ? field_byte_4 : _GEN_1202; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1363 = 8'h53 == total_offset_4 ? field_byte_4 : _GEN_1203; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1364 = 8'h54 == total_offset_4 ? field_byte_4 : _GEN_1204; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1365 = 8'h55 == total_offset_4 ? field_byte_4 : _GEN_1205; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1366 = 8'h56 == total_offset_4 ? field_byte_4 : _GEN_1206; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1367 = 8'h57 == total_offset_4 ? field_byte_4 : _GEN_1207; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1368 = 8'h58 == total_offset_4 ? field_byte_4 : _GEN_1208; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1369 = 8'h59 == total_offset_4 ? field_byte_4 : _GEN_1209; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1370 = 8'h5a == total_offset_4 ? field_byte_4 : _GEN_1210; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1371 = 8'h5b == total_offset_4 ? field_byte_4 : _GEN_1211; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1372 = 8'h5c == total_offset_4 ? field_byte_4 : _GEN_1212; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1373 = 8'h5d == total_offset_4 ? field_byte_4 : _GEN_1213; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1374 = 8'h5e == total_offset_4 ? field_byte_4 : _GEN_1214; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1375 = 8'h5f == total_offset_4 ? field_byte_4 : _GEN_1215; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1376 = 8'h60 == total_offset_4 ? field_byte_4 : _GEN_1216; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1377 = 8'h61 == total_offset_4 ? field_byte_4 : _GEN_1217; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1378 = 8'h62 == total_offset_4 ? field_byte_4 : _GEN_1218; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1379 = 8'h63 == total_offset_4 ? field_byte_4 : _GEN_1219; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1380 = 8'h64 == total_offset_4 ? field_byte_4 : _GEN_1220; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1381 = 8'h65 == total_offset_4 ? field_byte_4 : _GEN_1221; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1382 = 8'h66 == total_offset_4 ? field_byte_4 : _GEN_1222; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1383 = 8'h67 == total_offset_4 ? field_byte_4 : _GEN_1223; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1384 = 8'h68 == total_offset_4 ? field_byte_4 : _GEN_1224; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1385 = 8'h69 == total_offset_4 ? field_byte_4 : _GEN_1225; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1386 = 8'h6a == total_offset_4 ? field_byte_4 : _GEN_1226; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1387 = 8'h6b == total_offset_4 ? field_byte_4 : _GEN_1227; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1388 = 8'h6c == total_offset_4 ? field_byte_4 : _GEN_1228; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1389 = 8'h6d == total_offset_4 ? field_byte_4 : _GEN_1229; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1390 = 8'h6e == total_offset_4 ? field_byte_4 : _GEN_1230; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1391 = 8'h6f == total_offset_4 ? field_byte_4 : _GEN_1231; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1392 = 8'h70 == total_offset_4 ? field_byte_4 : _GEN_1232; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1393 = 8'h71 == total_offset_4 ? field_byte_4 : _GEN_1233; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1394 = 8'h72 == total_offset_4 ? field_byte_4 : _GEN_1234; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1395 = 8'h73 == total_offset_4 ? field_byte_4 : _GEN_1235; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1396 = 8'h74 == total_offset_4 ? field_byte_4 : _GEN_1236; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1397 = 8'h75 == total_offset_4 ? field_byte_4 : _GEN_1237; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1398 = 8'h76 == total_offset_4 ? field_byte_4 : _GEN_1238; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1399 = 8'h77 == total_offset_4 ? field_byte_4 : _GEN_1239; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1400 = 8'h78 == total_offset_4 ? field_byte_4 : _GEN_1240; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1401 = 8'h79 == total_offset_4 ? field_byte_4 : _GEN_1241; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1402 = 8'h7a == total_offset_4 ? field_byte_4 : _GEN_1242; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1403 = 8'h7b == total_offset_4 ? field_byte_4 : _GEN_1243; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1404 = 8'h7c == total_offset_4 ? field_byte_4 : _GEN_1244; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1405 = 8'h7d == total_offset_4 ? field_byte_4 : _GEN_1245; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1406 = 8'h7e == total_offset_4 ? field_byte_4 : _GEN_1246; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1407 = 8'h7f == total_offset_4 ? field_byte_4 : _GEN_1247; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1408 = 8'h80 == total_offset_4 ? field_byte_4 : _GEN_1248; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1409 = 8'h81 == total_offset_4 ? field_byte_4 : _GEN_1249; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1410 = 8'h82 == total_offset_4 ? field_byte_4 : _GEN_1250; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1411 = 8'h83 == total_offset_4 ? field_byte_4 : _GEN_1251; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1412 = 8'h84 == total_offset_4 ? field_byte_4 : _GEN_1252; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1413 = 8'h85 == total_offset_4 ? field_byte_4 : _GEN_1253; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1414 = 8'h86 == total_offset_4 ? field_byte_4 : _GEN_1254; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1415 = 8'h87 == total_offset_4 ? field_byte_4 : _GEN_1255; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1416 = 8'h88 == total_offset_4 ? field_byte_4 : _GEN_1256; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1417 = 8'h89 == total_offset_4 ? field_byte_4 : _GEN_1257; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1418 = 8'h8a == total_offset_4 ? field_byte_4 : _GEN_1258; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1419 = 8'h8b == total_offset_4 ? field_byte_4 : _GEN_1259; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1420 = 8'h8c == total_offset_4 ? field_byte_4 : _GEN_1260; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1421 = 8'h8d == total_offset_4 ? field_byte_4 : _GEN_1261; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1422 = 8'h8e == total_offset_4 ? field_byte_4 : _GEN_1262; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1423 = 8'h8f == total_offset_4 ? field_byte_4 : _GEN_1263; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1424 = 8'h90 == total_offset_4 ? field_byte_4 : _GEN_1264; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1425 = 8'h91 == total_offset_4 ? field_byte_4 : _GEN_1265; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1426 = 8'h92 == total_offset_4 ? field_byte_4 : _GEN_1266; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1427 = 8'h93 == total_offset_4 ? field_byte_4 : _GEN_1267; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1428 = 8'h94 == total_offset_4 ? field_byte_4 : _GEN_1268; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1429 = 8'h95 == total_offset_4 ? field_byte_4 : _GEN_1269; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1430 = 8'h96 == total_offset_4 ? field_byte_4 : _GEN_1270; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1431 = 8'h97 == total_offset_4 ? field_byte_4 : _GEN_1271; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1432 = 8'h98 == total_offset_4 ? field_byte_4 : _GEN_1272; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1433 = 8'h99 == total_offset_4 ? field_byte_4 : _GEN_1273; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1434 = 8'h9a == total_offset_4 ? field_byte_4 : _GEN_1274; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1435 = 8'h9b == total_offset_4 ? field_byte_4 : _GEN_1275; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1436 = 8'h9c == total_offset_4 ? field_byte_4 : _GEN_1276; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1437 = 8'h9d == total_offset_4 ? field_byte_4 : _GEN_1277; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1438 = 8'h9e == total_offset_4 ? field_byte_4 : _GEN_1278; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1439 = 8'h9f == total_offset_4 ? field_byte_4 : _GEN_1279; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1440 = 8'h4 < length_0 ? _GEN_1280 : _GEN_1120; // @[executor.scala 308:60]
  wire [7:0] _GEN_1441 = 8'h4 < length_0 ? _GEN_1281 : _GEN_1121; // @[executor.scala 308:60]
  wire [7:0] _GEN_1442 = 8'h4 < length_0 ? _GEN_1282 : _GEN_1122; // @[executor.scala 308:60]
  wire [7:0] _GEN_1443 = 8'h4 < length_0 ? _GEN_1283 : _GEN_1123; // @[executor.scala 308:60]
  wire [7:0] _GEN_1444 = 8'h4 < length_0 ? _GEN_1284 : _GEN_1124; // @[executor.scala 308:60]
  wire [7:0] _GEN_1445 = 8'h4 < length_0 ? _GEN_1285 : _GEN_1125; // @[executor.scala 308:60]
  wire [7:0] _GEN_1446 = 8'h4 < length_0 ? _GEN_1286 : _GEN_1126; // @[executor.scala 308:60]
  wire [7:0] _GEN_1447 = 8'h4 < length_0 ? _GEN_1287 : _GEN_1127; // @[executor.scala 308:60]
  wire [7:0] _GEN_1448 = 8'h4 < length_0 ? _GEN_1288 : _GEN_1128; // @[executor.scala 308:60]
  wire [7:0] _GEN_1449 = 8'h4 < length_0 ? _GEN_1289 : _GEN_1129; // @[executor.scala 308:60]
  wire [7:0] _GEN_1450 = 8'h4 < length_0 ? _GEN_1290 : _GEN_1130; // @[executor.scala 308:60]
  wire [7:0] _GEN_1451 = 8'h4 < length_0 ? _GEN_1291 : _GEN_1131; // @[executor.scala 308:60]
  wire [7:0] _GEN_1452 = 8'h4 < length_0 ? _GEN_1292 : _GEN_1132; // @[executor.scala 308:60]
  wire [7:0] _GEN_1453 = 8'h4 < length_0 ? _GEN_1293 : _GEN_1133; // @[executor.scala 308:60]
  wire [7:0] _GEN_1454 = 8'h4 < length_0 ? _GEN_1294 : _GEN_1134; // @[executor.scala 308:60]
  wire [7:0] _GEN_1455 = 8'h4 < length_0 ? _GEN_1295 : _GEN_1135; // @[executor.scala 308:60]
  wire [7:0] _GEN_1456 = 8'h4 < length_0 ? _GEN_1296 : _GEN_1136; // @[executor.scala 308:60]
  wire [7:0] _GEN_1457 = 8'h4 < length_0 ? _GEN_1297 : _GEN_1137; // @[executor.scala 308:60]
  wire [7:0] _GEN_1458 = 8'h4 < length_0 ? _GEN_1298 : _GEN_1138; // @[executor.scala 308:60]
  wire [7:0] _GEN_1459 = 8'h4 < length_0 ? _GEN_1299 : _GEN_1139; // @[executor.scala 308:60]
  wire [7:0] _GEN_1460 = 8'h4 < length_0 ? _GEN_1300 : _GEN_1140; // @[executor.scala 308:60]
  wire [7:0] _GEN_1461 = 8'h4 < length_0 ? _GEN_1301 : _GEN_1141; // @[executor.scala 308:60]
  wire [7:0] _GEN_1462 = 8'h4 < length_0 ? _GEN_1302 : _GEN_1142; // @[executor.scala 308:60]
  wire [7:0] _GEN_1463 = 8'h4 < length_0 ? _GEN_1303 : _GEN_1143; // @[executor.scala 308:60]
  wire [7:0] _GEN_1464 = 8'h4 < length_0 ? _GEN_1304 : _GEN_1144; // @[executor.scala 308:60]
  wire [7:0] _GEN_1465 = 8'h4 < length_0 ? _GEN_1305 : _GEN_1145; // @[executor.scala 308:60]
  wire [7:0] _GEN_1466 = 8'h4 < length_0 ? _GEN_1306 : _GEN_1146; // @[executor.scala 308:60]
  wire [7:0] _GEN_1467 = 8'h4 < length_0 ? _GEN_1307 : _GEN_1147; // @[executor.scala 308:60]
  wire [7:0] _GEN_1468 = 8'h4 < length_0 ? _GEN_1308 : _GEN_1148; // @[executor.scala 308:60]
  wire [7:0] _GEN_1469 = 8'h4 < length_0 ? _GEN_1309 : _GEN_1149; // @[executor.scala 308:60]
  wire [7:0] _GEN_1470 = 8'h4 < length_0 ? _GEN_1310 : _GEN_1150; // @[executor.scala 308:60]
  wire [7:0] _GEN_1471 = 8'h4 < length_0 ? _GEN_1311 : _GEN_1151; // @[executor.scala 308:60]
  wire [7:0] _GEN_1472 = 8'h4 < length_0 ? _GEN_1312 : _GEN_1152; // @[executor.scala 308:60]
  wire [7:0] _GEN_1473 = 8'h4 < length_0 ? _GEN_1313 : _GEN_1153; // @[executor.scala 308:60]
  wire [7:0] _GEN_1474 = 8'h4 < length_0 ? _GEN_1314 : _GEN_1154; // @[executor.scala 308:60]
  wire [7:0] _GEN_1475 = 8'h4 < length_0 ? _GEN_1315 : _GEN_1155; // @[executor.scala 308:60]
  wire [7:0] _GEN_1476 = 8'h4 < length_0 ? _GEN_1316 : _GEN_1156; // @[executor.scala 308:60]
  wire [7:0] _GEN_1477 = 8'h4 < length_0 ? _GEN_1317 : _GEN_1157; // @[executor.scala 308:60]
  wire [7:0] _GEN_1478 = 8'h4 < length_0 ? _GEN_1318 : _GEN_1158; // @[executor.scala 308:60]
  wire [7:0] _GEN_1479 = 8'h4 < length_0 ? _GEN_1319 : _GEN_1159; // @[executor.scala 308:60]
  wire [7:0] _GEN_1480 = 8'h4 < length_0 ? _GEN_1320 : _GEN_1160; // @[executor.scala 308:60]
  wire [7:0] _GEN_1481 = 8'h4 < length_0 ? _GEN_1321 : _GEN_1161; // @[executor.scala 308:60]
  wire [7:0] _GEN_1482 = 8'h4 < length_0 ? _GEN_1322 : _GEN_1162; // @[executor.scala 308:60]
  wire [7:0] _GEN_1483 = 8'h4 < length_0 ? _GEN_1323 : _GEN_1163; // @[executor.scala 308:60]
  wire [7:0] _GEN_1484 = 8'h4 < length_0 ? _GEN_1324 : _GEN_1164; // @[executor.scala 308:60]
  wire [7:0] _GEN_1485 = 8'h4 < length_0 ? _GEN_1325 : _GEN_1165; // @[executor.scala 308:60]
  wire [7:0] _GEN_1486 = 8'h4 < length_0 ? _GEN_1326 : _GEN_1166; // @[executor.scala 308:60]
  wire [7:0] _GEN_1487 = 8'h4 < length_0 ? _GEN_1327 : _GEN_1167; // @[executor.scala 308:60]
  wire [7:0] _GEN_1488 = 8'h4 < length_0 ? _GEN_1328 : _GEN_1168; // @[executor.scala 308:60]
  wire [7:0] _GEN_1489 = 8'h4 < length_0 ? _GEN_1329 : _GEN_1169; // @[executor.scala 308:60]
  wire [7:0] _GEN_1490 = 8'h4 < length_0 ? _GEN_1330 : _GEN_1170; // @[executor.scala 308:60]
  wire [7:0] _GEN_1491 = 8'h4 < length_0 ? _GEN_1331 : _GEN_1171; // @[executor.scala 308:60]
  wire [7:0] _GEN_1492 = 8'h4 < length_0 ? _GEN_1332 : _GEN_1172; // @[executor.scala 308:60]
  wire [7:0] _GEN_1493 = 8'h4 < length_0 ? _GEN_1333 : _GEN_1173; // @[executor.scala 308:60]
  wire [7:0] _GEN_1494 = 8'h4 < length_0 ? _GEN_1334 : _GEN_1174; // @[executor.scala 308:60]
  wire [7:0] _GEN_1495 = 8'h4 < length_0 ? _GEN_1335 : _GEN_1175; // @[executor.scala 308:60]
  wire [7:0] _GEN_1496 = 8'h4 < length_0 ? _GEN_1336 : _GEN_1176; // @[executor.scala 308:60]
  wire [7:0] _GEN_1497 = 8'h4 < length_0 ? _GEN_1337 : _GEN_1177; // @[executor.scala 308:60]
  wire [7:0] _GEN_1498 = 8'h4 < length_0 ? _GEN_1338 : _GEN_1178; // @[executor.scala 308:60]
  wire [7:0] _GEN_1499 = 8'h4 < length_0 ? _GEN_1339 : _GEN_1179; // @[executor.scala 308:60]
  wire [7:0] _GEN_1500 = 8'h4 < length_0 ? _GEN_1340 : _GEN_1180; // @[executor.scala 308:60]
  wire [7:0] _GEN_1501 = 8'h4 < length_0 ? _GEN_1341 : _GEN_1181; // @[executor.scala 308:60]
  wire [7:0] _GEN_1502 = 8'h4 < length_0 ? _GEN_1342 : _GEN_1182; // @[executor.scala 308:60]
  wire [7:0] _GEN_1503 = 8'h4 < length_0 ? _GEN_1343 : _GEN_1183; // @[executor.scala 308:60]
  wire [7:0] _GEN_1504 = 8'h4 < length_0 ? _GEN_1344 : _GEN_1184; // @[executor.scala 308:60]
  wire [7:0] _GEN_1505 = 8'h4 < length_0 ? _GEN_1345 : _GEN_1185; // @[executor.scala 308:60]
  wire [7:0] _GEN_1506 = 8'h4 < length_0 ? _GEN_1346 : _GEN_1186; // @[executor.scala 308:60]
  wire [7:0] _GEN_1507 = 8'h4 < length_0 ? _GEN_1347 : _GEN_1187; // @[executor.scala 308:60]
  wire [7:0] _GEN_1508 = 8'h4 < length_0 ? _GEN_1348 : _GEN_1188; // @[executor.scala 308:60]
  wire [7:0] _GEN_1509 = 8'h4 < length_0 ? _GEN_1349 : _GEN_1189; // @[executor.scala 308:60]
  wire [7:0] _GEN_1510 = 8'h4 < length_0 ? _GEN_1350 : _GEN_1190; // @[executor.scala 308:60]
  wire [7:0] _GEN_1511 = 8'h4 < length_0 ? _GEN_1351 : _GEN_1191; // @[executor.scala 308:60]
  wire [7:0] _GEN_1512 = 8'h4 < length_0 ? _GEN_1352 : _GEN_1192; // @[executor.scala 308:60]
  wire [7:0] _GEN_1513 = 8'h4 < length_0 ? _GEN_1353 : _GEN_1193; // @[executor.scala 308:60]
  wire [7:0] _GEN_1514 = 8'h4 < length_0 ? _GEN_1354 : _GEN_1194; // @[executor.scala 308:60]
  wire [7:0] _GEN_1515 = 8'h4 < length_0 ? _GEN_1355 : _GEN_1195; // @[executor.scala 308:60]
  wire [7:0] _GEN_1516 = 8'h4 < length_0 ? _GEN_1356 : _GEN_1196; // @[executor.scala 308:60]
  wire [7:0] _GEN_1517 = 8'h4 < length_0 ? _GEN_1357 : _GEN_1197; // @[executor.scala 308:60]
  wire [7:0] _GEN_1518 = 8'h4 < length_0 ? _GEN_1358 : _GEN_1198; // @[executor.scala 308:60]
  wire [7:0] _GEN_1519 = 8'h4 < length_0 ? _GEN_1359 : _GEN_1199; // @[executor.scala 308:60]
  wire [7:0] _GEN_1520 = 8'h4 < length_0 ? _GEN_1360 : _GEN_1200; // @[executor.scala 308:60]
  wire [7:0] _GEN_1521 = 8'h4 < length_0 ? _GEN_1361 : _GEN_1201; // @[executor.scala 308:60]
  wire [7:0] _GEN_1522 = 8'h4 < length_0 ? _GEN_1362 : _GEN_1202; // @[executor.scala 308:60]
  wire [7:0] _GEN_1523 = 8'h4 < length_0 ? _GEN_1363 : _GEN_1203; // @[executor.scala 308:60]
  wire [7:0] _GEN_1524 = 8'h4 < length_0 ? _GEN_1364 : _GEN_1204; // @[executor.scala 308:60]
  wire [7:0] _GEN_1525 = 8'h4 < length_0 ? _GEN_1365 : _GEN_1205; // @[executor.scala 308:60]
  wire [7:0] _GEN_1526 = 8'h4 < length_0 ? _GEN_1366 : _GEN_1206; // @[executor.scala 308:60]
  wire [7:0] _GEN_1527 = 8'h4 < length_0 ? _GEN_1367 : _GEN_1207; // @[executor.scala 308:60]
  wire [7:0] _GEN_1528 = 8'h4 < length_0 ? _GEN_1368 : _GEN_1208; // @[executor.scala 308:60]
  wire [7:0] _GEN_1529 = 8'h4 < length_0 ? _GEN_1369 : _GEN_1209; // @[executor.scala 308:60]
  wire [7:0] _GEN_1530 = 8'h4 < length_0 ? _GEN_1370 : _GEN_1210; // @[executor.scala 308:60]
  wire [7:0] _GEN_1531 = 8'h4 < length_0 ? _GEN_1371 : _GEN_1211; // @[executor.scala 308:60]
  wire [7:0] _GEN_1532 = 8'h4 < length_0 ? _GEN_1372 : _GEN_1212; // @[executor.scala 308:60]
  wire [7:0] _GEN_1533 = 8'h4 < length_0 ? _GEN_1373 : _GEN_1213; // @[executor.scala 308:60]
  wire [7:0] _GEN_1534 = 8'h4 < length_0 ? _GEN_1374 : _GEN_1214; // @[executor.scala 308:60]
  wire [7:0] _GEN_1535 = 8'h4 < length_0 ? _GEN_1375 : _GEN_1215; // @[executor.scala 308:60]
  wire [7:0] _GEN_1536 = 8'h4 < length_0 ? _GEN_1376 : _GEN_1216; // @[executor.scala 308:60]
  wire [7:0] _GEN_1537 = 8'h4 < length_0 ? _GEN_1377 : _GEN_1217; // @[executor.scala 308:60]
  wire [7:0] _GEN_1538 = 8'h4 < length_0 ? _GEN_1378 : _GEN_1218; // @[executor.scala 308:60]
  wire [7:0] _GEN_1539 = 8'h4 < length_0 ? _GEN_1379 : _GEN_1219; // @[executor.scala 308:60]
  wire [7:0] _GEN_1540 = 8'h4 < length_0 ? _GEN_1380 : _GEN_1220; // @[executor.scala 308:60]
  wire [7:0] _GEN_1541 = 8'h4 < length_0 ? _GEN_1381 : _GEN_1221; // @[executor.scala 308:60]
  wire [7:0] _GEN_1542 = 8'h4 < length_0 ? _GEN_1382 : _GEN_1222; // @[executor.scala 308:60]
  wire [7:0] _GEN_1543 = 8'h4 < length_0 ? _GEN_1383 : _GEN_1223; // @[executor.scala 308:60]
  wire [7:0] _GEN_1544 = 8'h4 < length_0 ? _GEN_1384 : _GEN_1224; // @[executor.scala 308:60]
  wire [7:0] _GEN_1545 = 8'h4 < length_0 ? _GEN_1385 : _GEN_1225; // @[executor.scala 308:60]
  wire [7:0] _GEN_1546 = 8'h4 < length_0 ? _GEN_1386 : _GEN_1226; // @[executor.scala 308:60]
  wire [7:0] _GEN_1547 = 8'h4 < length_0 ? _GEN_1387 : _GEN_1227; // @[executor.scala 308:60]
  wire [7:0] _GEN_1548 = 8'h4 < length_0 ? _GEN_1388 : _GEN_1228; // @[executor.scala 308:60]
  wire [7:0] _GEN_1549 = 8'h4 < length_0 ? _GEN_1389 : _GEN_1229; // @[executor.scala 308:60]
  wire [7:0] _GEN_1550 = 8'h4 < length_0 ? _GEN_1390 : _GEN_1230; // @[executor.scala 308:60]
  wire [7:0] _GEN_1551 = 8'h4 < length_0 ? _GEN_1391 : _GEN_1231; // @[executor.scala 308:60]
  wire [7:0] _GEN_1552 = 8'h4 < length_0 ? _GEN_1392 : _GEN_1232; // @[executor.scala 308:60]
  wire [7:0] _GEN_1553 = 8'h4 < length_0 ? _GEN_1393 : _GEN_1233; // @[executor.scala 308:60]
  wire [7:0] _GEN_1554 = 8'h4 < length_0 ? _GEN_1394 : _GEN_1234; // @[executor.scala 308:60]
  wire [7:0] _GEN_1555 = 8'h4 < length_0 ? _GEN_1395 : _GEN_1235; // @[executor.scala 308:60]
  wire [7:0] _GEN_1556 = 8'h4 < length_0 ? _GEN_1396 : _GEN_1236; // @[executor.scala 308:60]
  wire [7:0] _GEN_1557 = 8'h4 < length_0 ? _GEN_1397 : _GEN_1237; // @[executor.scala 308:60]
  wire [7:0] _GEN_1558 = 8'h4 < length_0 ? _GEN_1398 : _GEN_1238; // @[executor.scala 308:60]
  wire [7:0] _GEN_1559 = 8'h4 < length_0 ? _GEN_1399 : _GEN_1239; // @[executor.scala 308:60]
  wire [7:0] _GEN_1560 = 8'h4 < length_0 ? _GEN_1400 : _GEN_1240; // @[executor.scala 308:60]
  wire [7:0] _GEN_1561 = 8'h4 < length_0 ? _GEN_1401 : _GEN_1241; // @[executor.scala 308:60]
  wire [7:0] _GEN_1562 = 8'h4 < length_0 ? _GEN_1402 : _GEN_1242; // @[executor.scala 308:60]
  wire [7:0] _GEN_1563 = 8'h4 < length_0 ? _GEN_1403 : _GEN_1243; // @[executor.scala 308:60]
  wire [7:0] _GEN_1564 = 8'h4 < length_0 ? _GEN_1404 : _GEN_1244; // @[executor.scala 308:60]
  wire [7:0] _GEN_1565 = 8'h4 < length_0 ? _GEN_1405 : _GEN_1245; // @[executor.scala 308:60]
  wire [7:0] _GEN_1566 = 8'h4 < length_0 ? _GEN_1406 : _GEN_1246; // @[executor.scala 308:60]
  wire [7:0] _GEN_1567 = 8'h4 < length_0 ? _GEN_1407 : _GEN_1247; // @[executor.scala 308:60]
  wire [7:0] _GEN_1568 = 8'h4 < length_0 ? _GEN_1408 : _GEN_1248; // @[executor.scala 308:60]
  wire [7:0] _GEN_1569 = 8'h4 < length_0 ? _GEN_1409 : _GEN_1249; // @[executor.scala 308:60]
  wire [7:0] _GEN_1570 = 8'h4 < length_0 ? _GEN_1410 : _GEN_1250; // @[executor.scala 308:60]
  wire [7:0] _GEN_1571 = 8'h4 < length_0 ? _GEN_1411 : _GEN_1251; // @[executor.scala 308:60]
  wire [7:0] _GEN_1572 = 8'h4 < length_0 ? _GEN_1412 : _GEN_1252; // @[executor.scala 308:60]
  wire [7:0] _GEN_1573 = 8'h4 < length_0 ? _GEN_1413 : _GEN_1253; // @[executor.scala 308:60]
  wire [7:0] _GEN_1574 = 8'h4 < length_0 ? _GEN_1414 : _GEN_1254; // @[executor.scala 308:60]
  wire [7:0] _GEN_1575 = 8'h4 < length_0 ? _GEN_1415 : _GEN_1255; // @[executor.scala 308:60]
  wire [7:0] _GEN_1576 = 8'h4 < length_0 ? _GEN_1416 : _GEN_1256; // @[executor.scala 308:60]
  wire [7:0] _GEN_1577 = 8'h4 < length_0 ? _GEN_1417 : _GEN_1257; // @[executor.scala 308:60]
  wire [7:0] _GEN_1578 = 8'h4 < length_0 ? _GEN_1418 : _GEN_1258; // @[executor.scala 308:60]
  wire [7:0] _GEN_1579 = 8'h4 < length_0 ? _GEN_1419 : _GEN_1259; // @[executor.scala 308:60]
  wire [7:0] _GEN_1580 = 8'h4 < length_0 ? _GEN_1420 : _GEN_1260; // @[executor.scala 308:60]
  wire [7:0] _GEN_1581 = 8'h4 < length_0 ? _GEN_1421 : _GEN_1261; // @[executor.scala 308:60]
  wire [7:0] _GEN_1582 = 8'h4 < length_0 ? _GEN_1422 : _GEN_1262; // @[executor.scala 308:60]
  wire [7:0] _GEN_1583 = 8'h4 < length_0 ? _GEN_1423 : _GEN_1263; // @[executor.scala 308:60]
  wire [7:0] _GEN_1584 = 8'h4 < length_0 ? _GEN_1424 : _GEN_1264; // @[executor.scala 308:60]
  wire [7:0] _GEN_1585 = 8'h4 < length_0 ? _GEN_1425 : _GEN_1265; // @[executor.scala 308:60]
  wire [7:0] _GEN_1586 = 8'h4 < length_0 ? _GEN_1426 : _GEN_1266; // @[executor.scala 308:60]
  wire [7:0] _GEN_1587 = 8'h4 < length_0 ? _GEN_1427 : _GEN_1267; // @[executor.scala 308:60]
  wire [7:0] _GEN_1588 = 8'h4 < length_0 ? _GEN_1428 : _GEN_1268; // @[executor.scala 308:60]
  wire [7:0] _GEN_1589 = 8'h4 < length_0 ? _GEN_1429 : _GEN_1269; // @[executor.scala 308:60]
  wire [7:0] _GEN_1590 = 8'h4 < length_0 ? _GEN_1430 : _GEN_1270; // @[executor.scala 308:60]
  wire [7:0] _GEN_1591 = 8'h4 < length_0 ? _GEN_1431 : _GEN_1271; // @[executor.scala 308:60]
  wire [7:0] _GEN_1592 = 8'h4 < length_0 ? _GEN_1432 : _GEN_1272; // @[executor.scala 308:60]
  wire [7:0] _GEN_1593 = 8'h4 < length_0 ? _GEN_1433 : _GEN_1273; // @[executor.scala 308:60]
  wire [7:0] _GEN_1594 = 8'h4 < length_0 ? _GEN_1434 : _GEN_1274; // @[executor.scala 308:60]
  wire [7:0] _GEN_1595 = 8'h4 < length_0 ? _GEN_1435 : _GEN_1275; // @[executor.scala 308:60]
  wire [7:0] _GEN_1596 = 8'h4 < length_0 ? _GEN_1436 : _GEN_1276; // @[executor.scala 308:60]
  wire [7:0] _GEN_1597 = 8'h4 < length_0 ? _GEN_1437 : _GEN_1277; // @[executor.scala 308:60]
  wire [7:0] _GEN_1598 = 8'h4 < length_0 ? _GEN_1438 : _GEN_1278; // @[executor.scala 308:60]
  wire [7:0] _GEN_1599 = 8'h4 < length_0 ? _GEN_1439 : _GEN_1279; // @[executor.scala 308:60]
  wire [7:0] field_byte_5 = field_0[23:16]; // @[executor.scala 305:57]
  wire [7:0] total_offset_5 = offset_0 + 8'h5; // @[executor.scala 307:57]
  wire [7:0] _GEN_1600 = 8'h0 == total_offset_5 ? field_byte_5 : _GEN_1440; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1601 = 8'h1 == total_offset_5 ? field_byte_5 : _GEN_1441; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1602 = 8'h2 == total_offset_5 ? field_byte_5 : _GEN_1442; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1603 = 8'h3 == total_offset_5 ? field_byte_5 : _GEN_1443; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1604 = 8'h4 == total_offset_5 ? field_byte_5 : _GEN_1444; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1605 = 8'h5 == total_offset_5 ? field_byte_5 : _GEN_1445; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1606 = 8'h6 == total_offset_5 ? field_byte_5 : _GEN_1446; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1607 = 8'h7 == total_offset_5 ? field_byte_5 : _GEN_1447; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1608 = 8'h8 == total_offset_5 ? field_byte_5 : _GEN_1448; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1609 = 8'h9 == total_offset_5 ? field_byte_5 : _GEN_1449; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1610 = 8'ha == total_offset_5 ? field_byte_5 : _GEN_1450; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1611 = 8'hb == total_offset_5 ? field_byte_5 : _GEN_1451; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1612 = 8'hc == total_offset_5 ? field_byte_5 : _GEN_1452; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1613 = 8'hd == total_offset_5 ? field_byte_5 : _GEN_1453; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1614 = 8'he == total_offset_5 ? field_byte_5 : _GEN_1454; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1615 = 8'hf == total_offset_5 ? field_byte_5 : _GEN_1455; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1616 = 8'h10 == total_offset_5 ? field_byte_5 : _GEN_1456; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1617 = 8'h11 == total_offset_5 ? field_byte_5 : _GEN_1457; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1618 = 8'h12 == total_offset_5 ? field_byte_5 : _GEN_1458; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1619 = 8'h13 == total_offset_5 ? field_byte_5 : _GEN_1459; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1620 = 8'h14 == total_offset_5 ? field_byte_5 : _GEN_1460; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1621 = 8'h15 == total_offset_5 ? field_byte_5 : _GEN_1461; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1622 = 8'h16 == total_offset_5 ? field_byte_5 : _GEN_1462; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1623 = 8'h17 == total_offset_5 ? field_byte_5 : _GEN_1463; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1624 = 8'h18 == total_offset_5 ? field_byte_5 : _GEN_1464; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1625 = 8'h19 == total_offset_5 ? field_byte_5 : _GEN_1465; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1626 = 8'h1a == total_offset_5 ? field_byte_5 : _GEN_1466; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1627 = 8'h1b == total_offset_5 ? field_byte_5 : _GEN_1467; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1628 = 8'h1c == total_offset_5 ? field_byte_5 : _GEN_1468; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1629 = 8'h1d == total_offset_5 ? field_byte_5 : _GEN_1469; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1630 = 8'h1e == total_offset_5 ? field_byte_5 : _GEN_1470; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1631 = 8'h1f == total_offset_5 ? field_byte_5 : _GEN_1471; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1632 = 8'h20 == total_offset_5 ? field_byte_5 : _GEN_1472; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1633 = 8'h21 == total_offset_5 ? field_byte_5 : _GEN_1473; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1634 = 8'h22 == total_offset_5 ? field_byte_5 : _GEN_1474; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1635 = 8'h23 == total_offset_5 ? field_byte_5 : _GEN_1475; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1636 = 8'h24 == total_offset_5 ? field_byte_5 : _GEN_1476; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1637 = 8'h25 == total_offset_5 ? field_byte_5 : _GEN_1477; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1638 = 8'h26 == total_offset_5 ? field_byte_5 : _GEN_1478; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1639 = 8'h27 == total_offset_5 ? field_byte_5 : _GEN_1479; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1640 = 8'h28 == total_offset_5 ? field_byte_5 : _GEN_1480; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1641 = 8'h29 == total_offset_5 ? field_byte_5 : _GEN_1481; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1642 = 8'h2a == total_offset_5 ? field_byte_5 : _GEN_1482; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1643 = 8'h2b == total_offset_5 ? field_byte_5 : _GEN_1483; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1644 = 8'h2c == total_offset_5 ? field_byte_5 : _GEN_1484; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1645 = 8'h2d == total_offset_5 ? field_byte_5 : _GEN_1485; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1646 = 8'h2e == total_offset_5 ? field_byte_5 : _GEN_1486; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1647 = 8'h2f == total_offset_5 ? field_byte_5 : _GEN_1487; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1648 = 8'h30 == total_offset_5 ? field_byte_5 : _GEN_1488; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1649 = 8'h31 == total_offset_5 ? field_byte_5 : _GEN_1489; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1650 = 8'h32 == total_offset_5 ? field_byte_5 : _GEN_1490; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1651 = 8'h33 == total_offset_5 ? field_byte_5 : _GEN_1491; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1652 = 8'h34 == total_offset_5 ? field_byte_5 : _GEN_1492; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1653 = 8'h35 == total_offset_5 ? field_byte_5 : _GEN_1493; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1654 = 8'h36 == total_offset_5 ? field_byte_5 : _GEN_1494; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1655 = 8'h37 == total_offset_5 ? field_byte_5 : _GEN_1495; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1656 = 8'h38 == total_offset_5 ? field_byte_5 : _GEN_1496; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1657 = 8'h39 == total_offset_5 ? field_byte_5 : _GEN_1497; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1658 = 8'h3a == total_offset_5 ? field_byte_5 : _GEN_1498; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1659 = 8'h3b == total_offset_5 ? field_byte_5 : _GEN_1499; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1660 = 8'h3c == total_offset_5 ? field_byte_5 : _GEN_1500; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1661 = 8'h3d == total_offset_5 ? field_byte_5 : _GEN_1501; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1662 = 8'h3e == total_offset_5 ? field_byte_5 : _GEN_1502; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1663 = 8'h3f == total_offset_5 ? field_byte_5 : _GEN_1503; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1664 = 8'h40 == total_offset_5 ? field_byte_5 : _GEN_1504; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1665 = 8'h41 == total_offset_5 ? field_byte_5 : _GEN_1505; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1666 = 8'h42 == total_offset_5 ? field_byte_5 : _GEN_1506; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1667 = 8'h43 == total_offset_5 ? field_byte_5 : _GEN_1507; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1668 = 8'h44 == total_offset_5 ? field_byte_5 : _GEN_1508; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1669 = 8'h45 == total_offset_5 ? field_byte_5 : _GEN_1509; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1670 = 8'h46 == total_offset_5 ? field_byte_5 : _GEN_1510; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1671 = 8'h47 == total_offset_5 ? field_byte_5 : _GEN_1511; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1672 = 8'h48 == total_offset_5 ? field_byte_5 : _GEN_1512; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1673 = 8'h49 == total_offset_5 ? field_byte_5 : _GEN_1513; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1674 = 8'h4a == total_offset_5 ? field_byte_5 : _GEN_1514; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1675 = 8'h4b == total_offset_5 ? field_byte_5 : _GEN_1515; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1676 = 8'h4c == total_offset_5 ? field_byte_5 : _GEN_1516; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1677 = 8'h4d == total_offset_5 ? field_byte_5 : _GEN_1517; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1678 = 8'h4e == total_offset_5 ? field_byte_5 : _GEN_1518; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1679 = 8'h4f == total_offset_5 ? field_byte_5 : _GEN_1519; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1680 = 8'h50 == total_offset_5 ? field_byte_5 : _GEN_1520; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1681 = 8'h51 == total_offset_5 ? field_byte_5 : _GEN_1521; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1682 = 8'h52 == total_offset_5 ? field_byte_5 : _GEN_1522; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1683 = 8'h53 == total_offset_5 ? field_byte_5 : _GEN_1523; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1684 = 8'h54 == total_offset_5 ? field_byte_5 : _GEN_1524; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1685 = 8'h55 == total_offset_5 ? field_byte_5 : _GEN_1525; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1686 = 8'h56 == total_offset_5 ? field_byte_5 : _GEN_1526; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1687 = 8'h57 == total_offset_5 ? field_byte_5 : _GEN_1527; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1688 = 8'h58 == total_offset_5 ? field_byte_5 : _GEN_1528; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1689 = 8'h59 == total_offset_5 ? field_byte_5 : _GEN_1529; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1690 = 8'h5a == total_offset_5 ? field_byte_5 : _GEN_1530; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1691 = 8'h5b == total_offset_5 ? field_byte_5 : _GEN_1531; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1692 = 8'h5c == total_offset_5 ? field_byte_5 : _GEN_1532; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1693 = 8'h5d == total_offset_5 ? field_byte_5 : _GEN_1533; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1694 = 8'h5e == total_offset_5 ? field_byte_5 : _GEN_1534; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1695 = 8'h5f == total_offset_5 ? field_byte_5 : _GEN_1535; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1696 = 8'h60 == total_offset_5 ? field_byte_5 : _GEN_1536; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1697 = 8'h61 == total_offset_5 ? field_byte_5 : _GEN_1537; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1698 = 8'h62 == total_offset_5 ? field_byte_5 : _GEN_1538; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1699 = 8'h63 == total_offset_5 ? field_byte_5 : _GEN_1539; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1700 = 8'h64 == total_offset_5 ? field_byte_5 : _GEN_1540; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1701 = 8'h65 == total_offset_5 ? field_byte_5 : _GEN_1541; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1702 = 8'h66 == total_offset_5 ? field_byte_5 : _GEN_1542; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1703 = 8'h67 == total_offset_5 ? field_byte_5 : _GEN_1543; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1704 = 8'h68 == total_offset_5 ? field_byte_5 : _GEN_1544; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1705 = 8'h69 == total_offset_5 ? field_byte_5 : _GEN_1545; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1706 = 8'h6a == total_offset_5 ? field_byte_5 : _GEN_1546; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1707 = 8'h6b == total_offset_5 ? field_byte_5 : _GEN_1547; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1708 = 8'h6c == total_offset_5 ? field_byte_5 : _GEN_1548; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1709 = 8'h6d == total_offset_5 ? field_byte_5 : _GEN_1549; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1710 = 8'h6e == total_offset_5 ? field_byte_5 : _GEN_1550; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1711 = 8'h6f == total_offset_5 ? field_byte_5 : _GEN_1551; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1712 = 8'h70 == total_offset_5 ? field_byte_5 : _GEN_1552; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1713 = 8'h71 == total_offset_5 ? field_byte_5 : _GEN_1553; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1714 = 8'h72 == total_offset_5 ? field_byte_5 : _GEN_1554; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1715 = 8'h73 == total_offset_5 ? field_byte_5 : _GEN_1555; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1716 = 8'h74 == total_offset_5 ? field_byte_5 : _GEN_1556; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1717 = 8'h75 == total_offset_5 ? field_byte_5 : _GEN_1557; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1718 = 8'h76 == total_offset_5 ? field_byte_5 : _GEN_1558; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1719 = 8'h77 == total_offset_5 ? field_byte_5 : _GEN_1559; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1720 = 8'h78 == total_offset_5 ? field_byte_5 : _GEN_1560; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1721 = 8'h79 == total_offset_5 ? field_byte_5 : _GEN_1561; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1722 = 8'h7a == total_offset_5 ? field_byte_5 : _GEN_1562; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1723 = 8'h7b == total_offset_5 ? field_byte_5 : _GEN_1563; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1724 = 8'h7c == total_offset_5 ? field_byte_5 : _GEN_1564; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1725 = 8'h7d == total_offset_5 ? field_byte_5 : _GEN_1565; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1726 = 8'h7e == total_offset_5 ? field_byte_5 : _GEN_1566; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1727 = 8'h7f == total_offset_5 ? field_byte_5 : _GEN_1567; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1728 = 8'h80 == total_offset_5 ? field_byte_5 : _GEN_1568; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1729 = 8'h81 == total_offset_5 ? field_byte_5 : _GEN_1569; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1730 = 8'h82 == total_offset_5 ? field_byte_5 : _GEN_1570; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1731 = 8'h83 == total_offset_5 ? field_byte_5 : _GEN_1571; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1732 = 8'h84 == total_offset_5 ? field_byte_5 : _GEN_1572; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1733 = 8'h85 == total_offset_5 ? field_byte_5 : _GEN_1573; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1734 = 8'h86 == total_offset_5 ? field_byte_5 : _GEN_1574; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1735 = 8'h87 == total_offset_5 ? field_byte_5 : _GEN_1575; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1736 = 8'h88 == total_offset_5 ? field_byte_5 : _GEN_1576; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1737 = 8'h89 == total_offset_5 ? field_byte_5 : _GEN_1577; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1738 = 8'h8a == total_offset_5 ? field_byte_5 : _GEN_1578; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1739 = 8'h8b == total_offset_5 ? field_byte_5 : _GEN_1579; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1740 = 8'h8c == total_offset_5 ? field_byte_5 : _GEN_1580; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1741 = 8'h8d == total_offset_5 ? field_byte_5 : _GEN_1581; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1742 = 8'h8e == total_offset_5 ? field_byte_5 : _GEN_1582; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1743 = 8'h8f == total_offset_5 ? field_byte_5 : _GEN_1583; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1744 = 8'h90 == total_offset_5 ? field_byte_5 : _GEN_1584; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1745 = 8'h91 == total_offset_5 ? field_byte_5 : _GEN_1585; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1746 = 8'h92 == total_offset_5 ? field_byte_5 : _GEN_1586; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1747 = 8'h93 == total_offset_5 ? field_byte_5 : _GEN_1587; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1748 = 8'h94 == total_offset_5 ? field_byte_5 : _GEN_1588; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1749 = 8'h95 == total_offset_5 ? field_byte_5 : _GEN_1589; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1750 = 8'h96 == total_offset_5 ? field_byte_5 : _GEN_1590; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1751 = 8'h97 == total_offset_5 ? field_byte_5 : _GEN_1591; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1752 = 8'h98 == total_offset_5 ? field_byte_5 : _GEN_1592; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1753 = 8'h99 == total_offset_5 ? field_byte_5 : _GEN_1593; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1754 = 8'h9a == total_offset_5 ? field_byte_5 : _GEN_1594; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1755 = 8'h9b == total_offset_5 ? field_byte_5 : _GEN_1595; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1756 = 8'h9c == total_offset_5 ? field_byte_5 : _GEN_1596; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1757 = 8'h9d == total_offset_5 ? field_byte_5 : _GEN_1597; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1758 = 8'h9e == total_offset_5 ? field_byte_5 : _GEN_1598; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1759 = 8'h9f == total_offset_5 ? field_byte_5 : _GEN_1599; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1760 = 8'h5 < length_0 ? _GEN_1600 : _GEN_1440; // @[executor.scala 308:60]
  wire [7:0] _GEN_1761 = 8'h5 < length_0 ? _GEN_1601 : _GEN_1441; // @[executor.scala 308:60]
  wire [7:0] _GEN_1762 = 8'h5 < length_0 ? _GEN_1602 : _GEN_1442; // @[executor.scala 308:60]
  wire [7:0] _GEN_1763 = 8'h5 < length_0 ? _GEN_1603 : _GEN_1443; // @[executor.scala 308:60]
  wire [7:0] _GEN_1764 = 8'h5 < length_0 ? _GEN_1604 : _GEN_1444; // @[executor.scala 308:60]
  wire [7:0] _GEN_1765 = 8'h5 < length_0 ? _GEN_1605 : _GEN_1445; // @[executor.scala 308:60]
  wire [7:0] _GEN_1766 = 8'h5 < length_0 ? _GEN_1606 : _GEN_1446; // @[executor.scala 308:60]
  wire [7:0] _GEN_1767 = 8'h5 < length_0 ? _GEN_1607 : _GEN_1447; // @[executor.scala 308:60]
  wire [7:0] _GEN_1768 = 8'h5 < length_0 ? _GEN_1608 : _GEN_1448; // @[executor.scala 308:60]
  wire [7:0] _GEN_1769 = 8'h5 < length_0 ? _GEN_1609 : _GEN_1449; // @[executor.scala 308:60]
  wire [7:0] _GEN_1770 = 8'h5 < length_0 ? _GEN_1610 : _GEN_1450; // @[executor.scala 308:60]
  wire [7:0] _GEN_1771 = 8'h5 < length_0 ? _GEN_1611 : _GEN_1451; // @[executor.scala 308:60]
  wire [7:0] _GEN_1772 = 8'h5 < length_0 ? _GEN_1612 : _GEN_1452; // @[executor.scala 308:60]
  wire [7:0] _GEN_1773 = 8'h5 < length_0 ? _GEN_1613 : _GEN_1453; // @[executor.scala 308:60]
  wire [7:0] _GEN_1774 = 8'h5 < length_0 ? _GEN_1614 : _GEN_1454; // @[executor.scala 308:60]
  wire [7:0] _GEN_1775 = 8'h5 < length_0 ? _GEN_1615 : _GEN_1455; // @[executor.scala 308:60]
  wire [7:0] _GEN_1776 = 8'h5 < length_0 ? _GEN_1616 : _GEN_1456; // @[executor.scala 308:60]
  wire [7:0] _GEN_1777 = 8'h5 < length_0 ? _GEN_1617 : _GEN_1457; // @[executor.scala 308:60]
  wire [7:0] _GEN_1778 = 8'h5 < length_0 ? _GEN_1618 : _GEN_1458; // @[executor.scala 308:60]
  wire [7:0] _GEN_1779 = 8'h5 < length_0 ? _GEN_1619 : _GEN_1459; // @[executor.scala 308:60]
  wire [7:0] _GEN_1780 = 8'h5 < length_0 ? _GEN_1620 : _GEN_1460; // @[executor.scala 308:60]
  wire [7:0] _GEN_1781 = 8'h5 < length_0 ? _GEN_1621 : _GEN_1461; // @[executor.scala 308:60]
  wire [7:0] _GEN_1782 = 8'h5 < length_0 ? _GEN_1622 : _GEN_1462; // @[executor.scala 308:60]
  wire [7:0] _GEN_1783 = 8'h5 < length_0 ? _GEN_1623 : _GEN_1463; // @[executor.scala 308:60]
  wire [7:0] _GEN_1784 = 8'h5 < length_0 ? _GEN_1624 : _GEN_1464; // @[executor.scala 308:60]
  wire [7:0] _GEN_1785 = 8'h5 < length_0 ? _GEN_1625 : _GEN_1465; // @[executor.scala 308:60]
  wire [7:0] _GEN_1786 = 8'h5 < length_0 ? _GEN_1626 : _GEN_1466; // @[executor.scala 308:60]
  wire [7:0] _GEN_1787 = 8'h5 < length_0 ? _GEN_1627 : _GEN_1467; // @[executor.scala 308:60]
  wire [7:0] _GEN_1788 = 8'h5 < length_0 ? _GEN_1628 : _GEN_1468; // @[executor.scala 308:60]
  wire [7:0] _GEN_1789 = 8'h5 < length_0 ? _GEN_1629 : _GEN_1469; // @[executor.scala 308:60]
  wire [7:0] _GEN_1790 = 8'h5 < length_0 ? _GEN_1630 : _GEN_1470; // @[executor.scala 308:60]
  wire [7:0] _GEN_1791 = 8'h5 < length_0 ? _GEN_1631 : _GEN_1471; // @[executor.scala 308:60]
  wire [7:0] _GEN_1792 = 8'h5 < length_0 ? _GEN_1632 : _GEN_1472; // @[executor.scala 308:60]
  wire [7:0] _GEN_1793 = 8'h5 < length_0 ? _GEN_1633 : _GEN_1473; // @[executor.scala 308:60]
  wire [7:0] _GEN_1794 = 8'h5 < length_0 ? _GEN_1634 : _GEN_1474; // @[executor.scala 308:60]
  wire [7:0] _GEN_1795 = 8'h5 < length_0 ? _GEN_1635 : _GEN_1475; // @[executor.scala 308:60]
  wire [7:0] _GEN_1796 = 8'h5 < length_0 ? _GEN_1636 : _GEN_1476; // @[executor.scala 308:60]
  wire [7:0] _GEN_1797 = 8'h5 < length_0 ? _GEN_1637 : _GEN_1477; // @[executor.scala 308:60]
  wire [7:0] _GEN_1798 = 8'h5 < length_0 ? _GEN_1638 : _GEN_1478; // @[executor.scala 308:60]
  wire [7:0] _GEN_1799 = 8'h5 < length_0 ? _GEN_1639 : _GEN_1479; // @[executor.scala 308:60]
  wire [7:0] _GEN_1800 = 8'h5 < length_0 ? _GEN_1640 : _GEN_1480; // @[executor.scala 308:60]
  wire [7:0] _GEN_1801 = 8'h5 < length_0 ? _GEN_1641 : _GEN_1481; // @[executor.scala 308:60]
  wire [7:0] _GEN_1802 = 8'h5 < length_0 ? _GEN_1642 : _GEN_1482; // @[executor.scala 308:60]
  wire [7:0] _GEN_1803 = 8'h5 < length_0 ? _GEN_1643 : _GEN_1483; // @[executor.scala 308:60]
  wire [7:0] _GEN_1804 = 8'h5 < length_0 ? _GEN_1644 : _GEN_1484; // @[executor.scala 308:60]
  wire [7:0] _GEN_1805 = 8'h5 < length_0 ? _GEN_1645 : _GEN_1485; // @[executor.scala 308:60]
  wire [7:0] _GEN_1806 = 8'h5 < length_0 ? _GEN_1646 : _GEN_1486; // @[executor.scala 308:60]
  wire [7:0] _GEN_1807 = 8'h5 < length_0 ? _GEN_1647 : _GEN_1487; // @[executor.scala 308:60]
  wire [7:0] _GEN_1808 = 8'h5 < length_0 ? _GEN_1648 : _GEN_1488; // @[executor.scala 308:60]
  wire [7:0] _GEN_1809 = 8'h5 < length_0 ? _GEN_1649 : _GEN_1489; // @[executor.scala 308:60]
  wire [7:0] _GEN_1810 = 8'h5 < length_0 ? _GEN_1650 : _GEN_1490; // @[executor.scala 308:60]
  wire [7:0] _GEN_1811 = 8'h5 < length_0 ? _GEN_1651 : _GEN_1491; // @[executor.scala 308:60]
  wire [7:0] _GEN_1812 = 8'h5 < length_0 ? _GEN_1652 : _GEN_1492; // @[executor.scala 308:60]
  wire [7:0] _GEN_1813 = 8'h5 < length_0 ? _GEN_1653 : _GEN_1493; // @[executor.scala 308:60]
  wire [7:0] _GEN_1814 = 8'h5 < length_0 ? _GEN_1654 : _GEN_1494; // @[executor.scala 308:60]
  wire [7:0] _GEN_1815 = 8'h5 < length_0 ? _GEN_1655 : _GEN_1495; // @[executor.scala 308:60]
  wire [7:0] _GEN_1816 = 8'h5 < length_0 ? _GEN_1656 : _GEN_1496; // @[executor.scala 308:60]
  wire [7:0] _GEN_1817 = 8'h5 < length_0 ? _GEN_1657 : _GEN_1497; // @[executor.scala 308:60]
  wire [7:0] _GEN_1818 = 8'h5 < length_0 ? _GEN_1658 : _GEN_1498; // @[executor.scala 308:60]
  wire [7:0] _GEN_1819 = 8'h5 < length_0 ? _GEN_1659 : _GEN_1499; // @[executor.scala 308:60]
  wire [7:0] _GEN_1820 = 8'h5 < length_0 ? _GEN_1660 : _GEN_1500; // @[executor.scala 308:60]
  wire [7:0] _GEN_1821 = 8'h5 < length_0 ? _GEN_1661 : _GEN_1501; // @[executor.scala 308:60]
  wire [7:0] _GEN_1822 = 8'h5 < length_0 ? _GEN_1662 : _GEN_1502; // @[executor.scala 308:60]
  wire [7:0] _GEN_1823 = 8'h5 < length_0 ? _GEN_1663 : _GEN_1503; // @[executor.scala 308:60]
  wire [7:0] _GEN_1824 = 8'h5 < length_0 ? _GEN_1664 : _GEN_1504; // @[executor.scala 308:60]
  wire [7:0] _GEN_1825 = 8'h5 < length_0 ? _GEN_1665 : _GEN_1505; // @[executor.scala 308:60]
  wire [7:0] _GEN_1826 = 8'h5 < length_0 ? _GEN_1666 : _GEN_1506; // @[executor.scala 308:60]
  wire [7:0] _GEN_1827 = 8'h5 < length_0 ? _GEN_1667 : _GEN_1507; // @[executor.scala 308:60]
  wire [7:0] _GEN_1828 = 8'h5 < length_0 ? _GEN_1668 : _GEN_1508; // @[executor.scala 308:60]
  wire [7:0] _GEN_1829 = 8'h5 < length_0 ? _GEN_1669 : _GEN_1509; // @[executor.scala 308:60]
  wire [7:0] _GEN_1830 = 8'h5 < length_0 ? _GEN_1670 : _GEN_1510; // @[executor.scala 308:60]
  wire [7:0] _GEN_1831 = 8'h5 < length_0 ? _GEN_1671 : _GEN_1511; // @[executor.scala 308:60]
  wire [7:0] _GEN_1832 = 8'h5 < length_0 ? _GEN_1672 : _GEN_1512; // @[executor.scala 308:60]
  wire [7:0] _GEN_1833 = 8'h5 < length_0 ? _GEN_1673 : _GEN_1513; // @[executor.scala 308:60]
  wire [7:0] _GEN_1834 = 8'h5 < length_0 ? _GEN_1674 : _GEN_1514; // @[executor.scala 308:60]
  wire [7:0] _GEN_1835 = 8'h5 < length_0 ? _GEN_1675 : _GEN_1515; // @[executor.scala 308:60]
  wire [7:0] _GEN_1836 = 8'h5 < length_0 ? _GEN_1676 : _GEN_1516; // @[executor.scala 308:60]
  wire [7:0] _GEN_1837 = 8'h5 < length_0 ? _GEN_1677 : _GEN_1517; // @[executor.scala 308:60]
  wire [7:0] _GEN_1838 = 8'h5 < length_0 ? _GEN_1678 : _GEN_1518; // @[executor.scala 308:60]
  wire [7:0] _GEN_1839 = 8'h5 < length_0 ? _GEN_1679 : _GEN_1519; // @[executor.scala 308:60]
  wire [7:0] _GEN_1840 = 8'h5 < length_0 ? _GEN_1680 : _GEN_1520; // @[executor.scala 308:60]
  wire [7:0] _GEN_1841 = 8'h5 < length_0 ? _GEN_1681 : _GEN_1521; // @[executor.scala 308:60]
  wire [7:0] _GEN_1842 = 8'h5 < length_0 ? _GEN_1682 : _GEN_1522; // @[executor.scala 308:60]
  wire [7:0] _GEN_1843 = 8'h5 < length_0 ? _GEN_1683 : _GEN_1523; // @[executor.scala 308:60]
  wire [7:0] _GEN_1844 = 8'h5 < length_0 ? _GEN_1684 : _GEN_1524; // @[executor.scala 308:60]
  wire [7:0] _GEN_1845 = 8'h5 < length_0 ? _GEN_1685 : _GEN_1525; // @[executor.scala 308:60]
  wire [7:0] _GEN_1846 = 8'h5 < length_0 ? _GEN_1686 : _GEN_1526; // @[executor.scala 308:60]
  wire [7:0] _GEN_1847 = 8'h5 < length_0 ? _GEN_1687 : _GEN_1527; // @[executor.scala 308:60]
  wire [7:0] _GEN_1848 = 8'h5 < length_0 ? _GEN_1688 : _GEN_1528; // @[executor.scala 308:60]
  wire [7:0] _GEN_1849 = 8'h5 < length_0 ? _GEN_1689 : _GEN_1529; // @[executor.scala 308:60]
  wire [7:0] _GEN_1850 = 8'h5 < length_0 ? _GEN_1690 : _GEN_1530; // @[executor.scala 308:60]
  wire [7:0] _GEN_1851 = 8'h5 < length_0 ? _GEN_1691 : _GEN_1531; // @[executor.scala 308:60]
  wire [7:0] _GEN_1852 = 8'h5 < length_0 ? _GEN_1692 : _GEN_1532; // @[executor.scala 308:60]
  wire [7:0] _GEN_1853 = 8'h5 < length_0 ? _GEN_1693 : _GEN_1533; // @[executor.scala 308:60]
  wire [7:0] _GEN_1854 = 8'h5 < length_0 ? _GEN_1694 : _GEN_1534; // @[executor.scala 308:60]
  wire [7:0] _GEN_1855 = 8'h5 < length_0 ? _GEN_1695 : _GEN_1535; // @[executor.scala 308:60]
  wire [7:0] _GEN_1856 = 8'h5 < length_0 ? _GEN_1696 : _GEN_1536; // @[executor.scala 308:60]
  wire [7:0] _GEN_1857 = 8'h5 < length_0 ? _GEN_1697 : _GEN_1537; // @[executor.scala 308:60]
  wire [7:0] _GEN_1858 = 8'h5 < length_0 ? _GEN_1698 : _GEN_1538; // @[executor.scala 308:60]
  wire [7:0] _GEN_1859 = 8'h5 < length_0 ? _GEN_1699 : _GEN_1539; // @[executor.scala 308:60]
  wire [7:0] _GEN_1860 = 8'h5 < length_0 ? _GEN_1700 : _GEN_1540; // @[executor.scala 308:60]
  wire [7:0] _GEN_1861 = 8'h5 < length_0 ? _GEN_1701 : _GEN_1541; // @[executor.scala 308:60]
  wire [7:0] _GEN_1862 = 8'h5 < length_0 ? _GEN_1702 : _GEN_1542; // @[executor.scala 308:60]
  wire [7:0] _GEN_1863 = 8'h5 < length_0 ? _GEN_1703 : _GEN_1543; // @[executor.scala 308:60]
  wire [7:0] _GEN_1864 = 8'h5 < length_0 ? _GEN_1704 : _GEN_1544; // @[executor.scala 308:60]
  wire [7:0] _GEN_1865 = 8'h5 < length_0 ? _GEN_1705 : _GEN_1545; // @[executor.scala 308:60]
  wire [7:0] _GEN_1866 = 8'h5 < length_0 ? _GEN_1706 : _GEN_1546; // @[executor.scala 308:60]
  wire [7:0] _GEN_1867 = 8'h5 < length_0 ? _GEN_1707 : _GEN_1547; // @[executor.scala 308:60]
  wire [7:0] _GEN_1868 = 8'h5 < length_0 ? _GEN_1708 : _GEN_1548; // @[executor.scala 308:60]
  wire [7:0] _GEN_1869 = 8'h5 < length_0 ? _GEN_1709 : _GEN_1549; // @[executor.scala 308:60]
  wire [7:0] _GEN_1870 = 8'h5 < length_0 ? _GEN_1710 : _GEN_1550; // @[executor.scala 308:60]
  wire [7:0] _GEN_1871 = 8'h5 < length_0 ? _GEN_1711 : _GEN_1551; // @[executor.scala 308:60]
  wire [7:0] _GEN_1872 = 8'h5 < length_0 ? _GEN_1712 : _GEN_1552; // @[executor.scala 308:60]
  wire [7:0] _GEN_1873 = 8'h5 < length_0 ? _GEN_1713 : _GEN_1553; // @[executor.scala 308:60]
  wire [7:0] _GEN_1874 = 8'h5 < length_0 ? _GEN_1714 : _GEN_1554; // @[executor.scala 308:60]
  wire [7:0] _GEN_1875 = 8'h5 < length_0 ? _GEN_1715 : _GEN_1555; // @[executor.scala 308:60]
  wire [7:0] _GEN_1876 = 8'h5 < length_0 ? _GEN_1716 : _GEN_1556; // @[executor.scala 308:60]
  wire [7:0] _GEN_1877 = 8'h5 < length_0 ? _GEN_1717 : _GEN_1557; // @[executor.scala 308:60]
  wire [7:0] _GEN_1878 = 8'h5 < length_0 ? _GEN_1718 : _GEN_1558; // @[executor.scala 308:60]
  wire [7:0] _GEN_1879 = 8'h5 < length_0 ? _GEN_1719 : _GEN_1559; // @[executor.scala 308:60]
  wire [7:0] _GEN_1880 = 8'h5 < length_0 ? _GEN_1720 : _GEN_1560; // @[executor.scala 308:60]
  wire [7:0] _GEN_1881 = 8'h5 < length_0 ? _GEN_1721 : _GEN_1561; // @[executor.scala 308:60]
  wire [7:0] _GEN_1882 = 8'h5 < length_0 ? _GEN_1722 : _GEN_1562; // @[executor.scala 308:60]
  wire [7:0] _GEN_1883 = 8'h5 < length_0 ? _GEN_1723 : _GEN_1563; // @[executor.scala 308:60]
  wire [7:0] _GEN_1884 = 8'h5 < length_0 ? _GEN_1724 : _GEN_1564; // @[executor.scala 308:60]
  wire [7:0] _GEN_1885 = 8'h5 < length_0 ? _GEN_1725 : _GEN_1565; // @[executor.scala 308:60]
  wire [7:0] _GEN_1886 = 8'h5 < length_0 ? _GEN_1726 : _GEN_1566; // @[executor.scala 308:60]
  wire [7:0] _GEN_1887 = 8'h5 < length_0 ? _GEN_1727 : _GEN_1567; // @[executor.scala 308:60]
  wire [7:0] _GEN_1888 = 8'h5 < length_0 ? _GEN_1728 : _GEN_1568; // @[executor.scala 308:60]
  wire [7:0] _GEN_1889 = 8'h5 < length_0 ? _GEN_1729 : _GEN_1569; // @[executor.scala 308:60]
  wire [7:0] _GEN_1890 = 8'h5 < length_0 ? _GEN_1730 : _GEN_1570; // @[executor.scala 308:60]
  wire [7:0] _GEN_1891 = 8'h5 < length_0 ? _GEN_1731 : _GEN_1571; // @[executor.scala 308:60]
  wire [7:0] _GEN_1892 = 8'h5 < length_0 ? _GEN_1732 : _GEN_1572; // @[executor.scala 308:60]
  wire [7:0] _GEN_1893 = 8'h5 < length_0 ? _GEN_1733 : _GEN_1573; // @[executor.scala 308:60]
  wire [7:0] _GEN_1894 = 8'h5 < length_0 ? _GEN_1734 : _GEN_1574; // @[executor.scala 308:60]
  wire [7:0] _GEN_1895 = 8'h5 < length_0 ? _GEN_1735 : _GEN_1575; // @[executor.scala 308:60]
  wire [7:0] _GEN_1896 = 8'h5 < length_0 ? _GEN_1736 : _GEN_1576; // @[executor.scala 308:60]
  wire [7:0] _GEN_1897 = 8'h5 < length_0 ? _GEN_1737 : _GEN_1577; // @[executor.scala 308:60]
  wire [7:0] _GEN_1898 = 8'h5 < length_0 ? _GEN_1738 : _GEN_1578; // @[executor.scala 308:60]
  wire [7:0] _GEN_1899 = 8'h5 < length_0 ? _GEN_1739 : _GEN_1579; // @[executor.scala 308:60]
  wire [7:0] _GEN_1900 = 8'h5 < length_0 ? _GEN_1740 : _GEN_1580; // @[executor.scala 308:60]
  wire [7:0] _GEN_1901 = 8'h5 < length_0 ? _GEN_1741 : _GEN_1581; // @[executor.scala 308:60]
  wire [7:0] _GEN_1902 = 8'h5 < length_0 ? _GEN_1742 : _GEN_1582; // @[executor.scala 308:60]
  wire [7:0] _GEN_1903 = 8'h5 < length_0 ? _GEN_1743 : _GEN_1583; // @[executor.scala 308:60]
  wire [7:0] _GEN_1904 = 8'h5 < length_0 ? _GEN_1744 : _GEN_1584; // @[executor.scala 308:60]
  wire [7:0] _GEN_1905 = 8'h5 < length_0 ? _GEN_1745 : _GEN_1585; // @[executor.scala 308:60]
  wire [7:0] _GEN_1906 = 8'h5 < length_0 ? _GEN_1746 : _GEN_1586; // @[executor.scala 308:60]
  wire [7:0] _GEN_1907 = 8'h5 < length_0 ? _GEN_1747 : _GEN_1587; // @[executor.scala 308:60]
  wire [7:0] _GEN_1908 = 8'h5 < length_0 ? _GEN_1748 : _GEN_1588; // @[executor.scala 308:60]
  wire [7:0] _GEN_1909 = 8'h5 < length_0 ? _GEN_1749 : _GEN_1589; // @[executor.scala 308:60]
  wire [7:0] _GEN_1910 = 8'h5 < length_0 ? _GEN_1750 : _GEN_1590; // @[executor.scala 308:60]
  wire [7:0] _GEN_1911 = 8'h5 < length_0 ? _GEN_1751 : _GEN_1591; // @[executor.scala 308:60]
  wire [7:0] _GEN_1912 = 8'h5 < length_0 ? _GEN_1752 : _GEN_1592; // @[executor.scala 308:60]
  wire [7:0] _GEN_1913 = 8'h5 < length_0 ? _GEN_1753 : _GEN_1593; // @[executor.scala 308:60]
  wire [7:0] _GEN_1914 = 8'h5 < length_0 ? _GEN_1754 : _GEN_1594; // @[executor.scala 308:60]
  wire [7:0] _GEN_1915 = 8'h5 < length_0 ? _GEN_1755 : _GEN_1595; // @[executor.scala 308:60]
  wire [7:0] _GEN_1916 = 8'h5 < length_0 ? _GEN_1756 : _GEN_1596; // @[executor.scala 308:60]
  wire [7:0] _GEN_1917 = 8'h5 < length_0 ? _GEN_1757 : _GEN_1597; // @[executor.scala 308:60]
  wire [7:0] _GEN_1918 = 8'h5 < length_0 ? _GEN_1758 : _GEN_1598; // @[executor.scala 308:60]
  wire [7:0] _GEN_1919 = 8'h5 < length_0 ? _GEN_1759 : _GEN_1599; // @[executor.scala 308:60]
  wire [7:0] field_byte_6 = field_0[15:8]; // @[executor.scala 305:57]
  wire [7:0] total_offset_6 = offset_0 + 8'h6; // @[executor.scala 307:57]
  wire [7:0] _GEN_1920 = 8'h0 == total_offset_6 ? field_byte_6 : _GEN_1760; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1921 = 8'h1 == total_offset_6 ? field_byte_6 : _GEN_1761; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1922 = 8'h2 == total_offset_6 ? field_byte_6 : _GEN_1762; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1923 = 8'h3 == total_offset_6 ? field_byte_6 : _GEN_1763; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1924 = 8'h4 == total_offset_6 ? field_byte_6 : _GEN_1764; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1925 = 8'h5 == total_offset_6 ? field_byte_6 : _GEN_1765; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1926 = 8'h6 == total_offset_6 ? field_byte_6 : _GEN_1766; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1927 = 8'h7 == total_offset_6 ? field_byte_6 : _GEN_1767; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1928 = 8'h8 == total_offset_6 ? field_byte_6 : _GEN_1768; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1929 = 8'h9 == total_offset_6 ? field_byte_6 : _GEN_1769; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1930 = 8'ha == total_offset_6 ? field_byte_6 : _GEN_1770; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1931 = 8'hb == total_offset_6 ? field_byte_6 : _GEN_1771; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1932 = 8'hc == total_offset_6 ? field_byte_6 : _GEN_1772; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1933 = 8'hd == total_offset_6 ? field_byte_6 : _GEN_1773; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1934 = 8'he == total_offset_6 ? field_byte_6 : _GEN_1774; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1935 = 8'hf == total_offset_6 ? field_byte_6 : _GEN_1775; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1936 = 8'h10 == total_offset_6 ? field_byte_6 : _GEN_1776; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1937 = 8'h11 == total_offset_6 ? field_byte_6 : _GEN_1777; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1938 = 8'h12 == total_offset_6 ? field_byte_6 : _GEN_1778; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1939 = 8'h13 == total_offset_6 ? field_byte_6 : _GEN_1779; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1940 = 8'h14 == total_offset_6 ? field_byte_6 : _GEN_1780; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1941 = 8'h15 == total_offset_6 ? field_byte_6 : _GEN_1781; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1942 = 8'h16 == total_offset_6 ? field_byte_6 : _GEN_1782; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1943 = 8'h17 == total_offset_6 ? field_byte_6 : _GEN_1783; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1944 = 8'h18 == total_offset_6 ? field_byte_6 : _GEN_1784; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1945 = 8'h19 == total_offset_6 ? field_byte_6 : _GEN_1785; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1946 = 8'h1a == total_offset_6 ? field_byte_6 : _GEN_1786; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1947 = 8'h1b == total_offset_6 ? field_byte_6 : _GEN_1787; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1948 = 8'h1c == total_offset_6 ? field_byte_6 : _GEN_1788; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1949 = 8'h1d == total_offset_6 ? field_byte_6 : _GEN_1789; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1950 = 8'h1e == total_offset_6 ? field_byte_6 : _GEN_1790; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1951 = 8'h1f == total_offset_6 ? field_byte_6 : _GEN_1791; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1952 = 8'h20 == total_offset_6 ? field_byte_6 : _GEN_1792; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1953 = 8'h21 == total_offset_6 ? field_byte_6 : _GEN_1793; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1954 = 8'h22 == total_offset_6 ? field_byte_6 : _GEN_1794; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1955 = 8'h23 == total_offset_6 ? field_byte_6 : _GEN_1795; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1956 = 8'h24 == total_offset_6 ? field_byte_6 : _GEN_1796; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1957 = 8'h25 == total_offset_6 ? field_byte_6 : _GEN_1797; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1958 = 8'h26 == total_offset_6 ? field_byte_6 : _GEN_1798; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1959 = 8'h27 == total_offset_6 ? field_byte_6 : _GEN_1799; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1960 = 8'h28 == total_offset_6 ? field_byte_6 : _GEN_1800; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1961 = 8'h29 == total_offset_6 ? field_byte_6 : _GEN_1801; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1962 = 8'h2a == total_offset_6 ? field_byte_6 : _GEN_1802; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1963 = 8'h2b == total_offset_6 ? field_byte_6 : _GEN_1803; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1964 = 8'h2c == total_offset_6 ? field_byte_6 : _GEN_1804; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1965 = 8'h2d == total_offset_6 ? field_byte_6 : _GEN_1805; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1966 = 8'h2e == total_offset_6 ? field_byte_6 : _GEN_1806; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1967 = 8'h2f == total_offset_6 ? field_byte_6 : _GEN_1807; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1968 = 8'h30 == total_offset_6 ? field_byte_6 : _GEN_1808; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1969 = 8'h31 == total_offset_6 ? field_byte_6 : _GEN_1809; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1970 = 8'h32 == total_offset_6 ? field_byte_6 : _GEN_1810; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1971 = 8'h33 == total_offset_6 ? field_byte_6 : _GEN_1811; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1972 = 8'h34 == total_offset_6 ? field_byte_6 : _GEN_1812; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1973 = 8'h35 == total_offset_6 ? field_byte_6 : _GEN_1813; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1974 = 8'h36 == total_offset_6 ? field_byte_6 : _GEN_1814; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1975 = 8'h37 == total_offset_6 ? field_byte_6 : _GEN_1815; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1976 = 8'h38 == total_offset_6 ? field_byte_6 : _GEN_1816; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1977 = 8'h39 == total_offset_6 ? field_byte_6 : _GEN_1817; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1978 = 8'h3a == total_offset_6 ? field_byte_6 : _GEN_1818; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1979 = 8'h3b == total_offset_6 ? field_byte_6 : _GEN_1819; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1980 = 8'h3c == total_offset_6 ? field_byte_6 : _GEN_1820; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1981 = 8'h3d == total_offset_6 ? field_byte_6 : _GEN_1821; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1982 = 8'h3e == total_offset_6 ? field_byte_6 : _GEN_1822; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1983 = 8'h3f == total_offset_6 ? field_byte_6 : _GEN_1823; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1984 = 8'h40 == total_offset_6 ? field_byte_6 : _GEN_1824; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1985 = 8'h41 == total_offset_6 ? field_byte_6 : _GEN_1825; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1986 = 8'h42 == total_offset_6 ? field_byte_6 : _GEN_1826; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1987 = 8'h43 == total_offset_6 ? field_byte_6 : _GEN_1827; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1988 = 8'h44 == total_offset_6 ? field_byte_6 : _GEN_1828; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1989 = 8'h45 == total_offset_6 ? field_byte_6 : _GEN_1829; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1990 = 8'h46 == total_offset_6 ? field_byte_6 : _GEN_1830; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1991 = 8'h47 == total_offset_6 ? field_byte_6 : _GEN_1831; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1992 = 8'h48 == total_offset_6 ? field_byte_6 : _GEN_1832; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1993 = 8'h49 == total_offset_6 ? field_byte_6 : _GEN_1833; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1994 = 8'h4a == total_offset_6 ? field_byte_6 : _GEN_1834; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1995 = 8'h4b == total_offset_6 ? field_byte_6 : _GEN_1835; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1996 = 8'h4c == total_offset_6 ? field_byte_6 : _GEN_1836; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1997 = 8'h4d == total_offset_6 ? field_byte_6 : _GEN_1837; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1998 = 8'h4e == total_offset_6 ? field_byte_6 : _GEN_1838; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_1999 = 8'h4f == total_offset_6 ? field_byte_6 : _GEN_1839; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2000 = 8'h50 == total_offset_6 ? field_byte_6 : _GEN_1840; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2001 = 8'h51 == total_offset_6 ? field_byte_6 : _GEN_1841; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2002 = 8'h52 == total_offset_6 ? field_byte_6 : _GEN_1842; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2003 = 8'h53 == total_offset_6 ? field_byte_6 : _GEN_1843; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2004 = 8'h54 == total_offset_6 ? field_byte_6 : _GEN_1844; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2005 = 8'h55 == total_offset_6 ? field_byte_6 : _GEN_1845; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2006 = 8'h56 == total_offset_6 ? field_byte_6 : _GEN_1846; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2007 = 8'h57 == total_offset_6 ? field_byte_6 : _GEN_1847; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2008 = 8'h58 == total_offset_6 ? field_byte_6 : _GEN_1848; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2009 = 8'h59 == total_offset_6 ? field_byte_6 : _GEN_1849; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2010 = 8'h5a == total_offset_6 ? field_byte_6 : _GEN_1850; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2011 = 8'h5b == total_offset_6 ? field_byte_6 : _GEN_1851; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2012 = 8'h5c == total_offset_6 ? field_byte_6 : _GEN_1852; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2013 = 8'h5d == total_offset_6 ? field_byte_6 : _GEN_1853; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2014 = 8'h5e == total_offset_6 ? field_byte_6 : _GEN_1854; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2015 = 8'h5f == total_offset_6 ? field_byte_6 : _GEN_1855; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2016 = 8'h60 == total_offset_6 ? field_byte_6 : _GEN_1856; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2017 = 8'h61 == total_offset_6 ? field_byte_6 : _GEN_1857; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2018 = 8'h62 == total_offset_6 ? field_byte_6 : _GEN_1858; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2019 = 8'h63 == total_offset_6 ? field_byte_6 : _GEN_1859; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2020 = 8'h64 == total_offset_6 ? field_byte_6 : _GEN_1860; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2021 = 8'h65 == total_offset_6 ? field_byte_6 : _GEN_1861; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2022 = 8'h66 == total_offset_6 ? field_byte_6 : _GEN_1862; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2023 = 8'h67 == total_offset_6 ? field_byte_6 : _GEN_1863; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2024 = 8'h68 == total_offset_6 ? field_byte_6 : _GEN_1864; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2025 = 8'h69 == total_offset_6 ? field_byte_6 : _GEN_1865; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2026 = 8'h6a == total_offset_6 ? field_byte_6 : _GEN_1866; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2027 = 8'h6b == total_offset_6 ? field_byte_6 : _GEN_1867; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2028 = 8'h6c == total_offset_6 ? field_byte_6 : _GEN_1868; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2029 = 8'h6d == total_offset_6 ? field_byte_6 : _GEN_1869; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2030 = 8'h6e == total_offset_6 ? field_byte_6 : _GEN_1870; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2031 = 8'h6f == total_offset_6 ? field_byte_6 : _GEN_1871; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2032 = 8'h70 == total_offset_6 ? field_byte_6 : _GEN_1872; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2033 = 8'h71 == total_offset_6 ? field_byte_6 : _GEN_1873; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2034 = 8'h72 == total_offset_6 ? field_byte_6 : _GEN_1874; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2035 = 8'h73 == total_offset_6 ? field_byte_6 : _GEN_1875; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2036 = 8'h74 == total_offset_6 ? field_byte_6 : _GEN_1876; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2037 = 8'h75 == total_offset_6 ? field_byte_6 : _GEN_1877; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2038 = 8'h76 == total_offset_6 ? field_byte_6 : _GEN_1878; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2039 = 8'h77 == total_offset_6 ? field_byte_6 : _GEN_1879; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2040 = 8'h78 == total_offset_6 ? field_byte_6 : _GEN_1880; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2041 = 8'h79 == total_offset_6 ? field_byte_6 : _GEN_1881; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2042 = 8'h7a == total_offset_6 ? field_byte_6 : _GEN_1882; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2043 = 8'h7b == total_offset_6 ? field_byte_6 : _GEN_1883; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2044 = 8'h7c == total_offset_6 ? field_byte_6 : _GEN_1884; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2045 = 8'h7d == total_offset_6 ? field_byte_6 : _GEN_1885; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2046 = 8'h7e == total_offset_6 ? field_byte_6 : _GEN_1886; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2047 = 8'h7f == total_offset_6 ? field_byte_6 : _GEN_1887; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2048 = 8'h80 == total_offset_6 ? field_byte_6 : _GEN_1888; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2049 = 8'h81 == total_offset_6 ? field_byte_6 : _GEN_1889; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2050 = 8'h82 == total_offset_6 ? field_byte_6 : _GEN_1890; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2051 = 8'h83 == total_offset_6 ? field_byte_6 : _GEN_1891; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2052 = 8'h84 == total_offset_6 ? field_byte_6 : _GEN_1892; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2053 = 8'h85 == total_offset_6 ? field_byte_6 : _GEN_1893; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2054 = 8'h86 == total_offset_6 ? field_byte_6 : _GEN_1894; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2055 = 8'h87 == total_offset_6 ? field_byte_6 : _GEN_1895; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2056 = 8'h88 == total_offset_6 ? field_byte_6 : _GEN_1896; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2057 = 8'h89 == total_offset_6 ? field_byte_6 : _GEN_1897; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2058 = 8'h8a == total_offset_6 ? field_byte_6 : _GEN_1898; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2059 = 8'h8b == total_offset_6 ? field_byte_6 : _GEN_1899; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2060 = 8'h8c == total_offset_6 ? field_byte_6 : _GEN_1900; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2061 = 8'h8d == total_offset_6 ? field_byte_6 : _GEN_1901; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2062 = 8'h8e == total_offset_6 ? field_byte_6 : _GEN_1902; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2063 = 8'h8f == total_offset_6 ? field_byte_6 : _GEN_1903; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2064 = 8'h90 == total_offset_6 ? field_byte_6 : _GEN_1904; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2065 = 8'h91 == total_offset_6 ? field_byte_6 : _GEN_1905; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2066 = 8'h92 == total_offset_6 ? field_byte_6 : _GEN_1906; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2067 = 8'h93 == total_offset_6 ? field_byte_6 : _GEN_1907; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2068 = 8'h94 == total_offset_6 ? field_byte_6 : _GEN_1908; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2069 = 8'h95 == total_offset_6 ? field_byte_6 : _GEN_1909; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2070 = 8'h96 == total_offset_6 ? field_byte_6 : _GEN_1910; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2071 = 8'h97 == total_offset_6 ? field_byte_6 : _GEN_1911; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2072 = 8'h98 == total_offset_6 ? field_byte_6 : _GEN_1912; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2073 = 8'h99 == total_offset_6 ? field_byte_6 : _GEN_1913; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2074 = 8'h9a == total_offset_6 ? field_byte_6 : _GEN_1914; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2075 = 8'h9b == total_offset_6 ? field_byte_6 : _GEN_1915; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2076 = 8'h9c == total_offset_6 ? field_byte_6 : _GEN_1916; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2077 = 8'h9d == total_offset_6 ? field_byte_6 : _GEN_1917; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2078 = 8'h9e == total_offset_6 ? field_byte_6 : _GEN_1918; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2079 = 8'h9f == total_offset_6 ? field_byte_6 : _GEN_1919; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2080 = 8'h6 < length_0 ? _GEN_1920 : _GEN_1760; // @[executor.scala 308:60]
  wire [7:0] _GEN_2081 = 8'h6 < length_0 ? _GEN_1921 : _GEN_1761; // @[executor.scala 308:60]
  wire [7:0] _GEN_2082 = 8'h6 < length_0 ? _GEN_1922 : _GEN_1762; // @[executor.scala 308:60]
  wire [7:0] _GEN_2083 = 8'h6 < length_0 ? _GEN_1923 : _GEN_1763; // @[executor.scala 308:60]
  wire [7:0] _GEN_2084 = 8'h6 < length_0 ? _GEN_1924 : _GEN_1764; // @[executor.scala 308:60]
  wire [7:0] _GEN_2085 = 8'h6 < length_0 ? _GEN_1925 : _GEN_1765; // @[executor.scala 308:60]
  wire [7:0] _GEN_2086 = 8'h6 < length_0 ? _GEN_1926 : _GEN_1766; // @[executor.scala 308:60]
  wire [7:0] _GEN_2087 = 8'h6 < length_0 ? _GEN_1927 : _GEN_1767; // @[executor.scala 308:60]
  wire [7:0] _GEN_2088 = 8'h6 < length_0 ? _GEN_1928 : _GEN_1768; // @[executor.scala 308:60]
  wire [7:0] _GEN_2089 = 8'h6 < length_0 ? _GEN_1929 : _GEN_1769; // @[executor.scala 308:60]
  wire [7:0] _GEN_2090 = 8'h6 < length_0 ? _GEN_1930 : _GEN_1770; // @[executor.scala 308:60]
  wire [7:0] _GEN_2091 = 8'h6 < length_0 ? _GEN_1931 : _GEN_1771; // @[executor.scala 308:60]
  wire [7:0] _GEN_2092 = 8'h6 < length_0 ? _GEN_1932 : _GEN_1772; // @[executor.scala 308:60]
  wire [7:0] _GEN_2093 = 8'h6 < length_0 ? _GEN_1933 : _GEN_1773; // @[executor.scala 308:60]
  wire [7:0] _GEN_2094 = 8'h6 < length_0 ? _GEN_1934 : _GEN_1774; // @[executor.scala 308:60]
  wire [7:0] _GEN_2095 = 8'h6 < length_0 ? _GEN_1935 : _GEN_1775; // @[executor.scala 308:60]
  wire [7:0] _GEN_2096 = 8'h6 < length_0 ? _GEN_1936 : _GEN_1776; // @[executor.scala 308:60]
  wire [7:0] _GEN_2097 = 8'h6 < length_0 ? _GEN_1937 : _GEN_1777; // @[executor.scala 308:60]
  wire [7:0] _GEN_2098 = 8'h6 < length_0 ? _GEN_1938 : _GEN_1778; // @[executor.scala 308:60]
  wire [7:0] _GEN_2099 = 8'h6 < length_0 ? _GEN_1939 : _GEN_1779; // @[executor.scala 308:60]
  wire [7:0] _GEN_2100 = 8'h6 < length_0 ? _GEN_1940 : _GEN_1780; // @[executor.scala 308:60]
  wire [7:0] _GEN_2101 = 8'h6 < length_0 ? _GEN_1941 : _GEN_1781; // @[executor.scala 308:60]
  wire [7:0] _GEN_2102 = 8'h6 < length_0 ? _GEN_1942 : _GEN_1782; // @[executor.scala 308:60]
  wire [7:0] _GEN_2103 = 8'h6 < length_0 ? _GEN_1943 : _GEN_1783; // @[executor.scala 308:60]
  wire [7:0] _GEN_2104 = 8'h6 < length_0 ? _GEN_1944 : _GEN_1784; // @[executor.scala 308:60]
  wire [7:0] _GEN_2105 = 8'h6 < length_0 ? _GEN_1945 : _GEN_1785; // @[executor.scala 308:60]
  wire [7:0] _GEN_2106 = 8'h6 < length_0 ? _GEN_1946 : _GEN_1786; // @[executor.scala 308:60]
  wire [7:0] _GEN_2107 = 8'h6 < length_0 ? _GEN_1947 : _GEN_1787; // @[executor.scala 308:60]
  wire [7:0] _GEN_2108 = 8'h6 < length_0 ? _GEN_1948 : _GEN_1788; // @[executor.scala 308:60]
  wire [7:0] _GEN_2109 = 8'h6 < length_0 ? _GEN_1949 : _GEN_1789; // @[executor.scala 308:60]
  wire [7:0] _GEN_2110 = 8'h6 < length_0 ? _GEN_1950 : _GEN_1790; // @[executor.scala 308:60]
  wire [7:0] _GEN_2111 = 8'h6 < length_0 ? _GEN_1951 : _GEN_1791; // @[executor.scala 308:60]
  wire [7:0] _GEN_2112 = 8'h6 < length_0 ? _GEN_1952 : _GEN_1792; // @[executor.scala 308:60]
  wire [7:0] _GEN_2113 = 8'h6 < length_0 ? _GEN_1953 : _GEN_1793; // @[executor.scala 308:60]
  wire [7:0] _GEN_2114 = 8'h6 < length_0 ? _GEN_1954 : _GEN_1794; // @[executor.scala 308:60]
  wire [7:0] _GEN_2115 = 8'h6 < length_0 ? _GEN_1955 : _GEN_1795; // @[executor.scala 308:60]
  wire [7:0] _GEN_2116 = 8'h6 < length_0 ? _GEN_1956 : _GEN_1796; // @[executor.scala 308:60]
  wire [7:0] _GEN_2117 = 8'h6 < length_0 ? _GEN_1957 : _GEN_1797; // @[executor.scala 308:60]
  wire [7:0] _GEN_2118 = 8'h6 < length_0 ? _GEN_1958 : _GEN_1798; // @[executor.scala 308:60]
  wire [7:0] _GEN_2119 = 8'h6 < length_0 ? _GEN_1959 : _GEN_1799; // @[executor.scala 308:60]
  wire [7:0] _GEN_2120 = 8'h6 < length_0 ? _GEN_1960 : _GEN_1800; // @[executor.scala 308:60]
  wire [7:0] _GEN_2121 = 8'h6 < length_0 ? _GEN_1961 : _GEN_1801; // @[executor.scala 308:60]
  wire [7:0] _GEN_2122 = 8'h6 < length_0 ? _GEN_1962 : _GEN_1802; // @[executor.scala 308:60]
  wire [7:0] _GEN_2123 = 8'h6 < length_0 ? _GEN_1963 : _GEN_1803; // @[executor.scala 308:60]
  wire [7:0] _GEN_2124 = 8'h6 < length_0 ? _GEN_1964 : _GEN_1804; // @[executor.scala 308:60]
  wire [7:0] _GEN_2125 = 8'h6 < length_0 ? _GEN_1965 : _GEN_1805; // @[executor.scala 308:60]
  wire [7:0] _GEN_2126 = 8'h6 < length_0 ? _GEN_1966 : _GEN_1806; // @[executor.scala 308:60]
  wire [7:0] _GEN_2127 = 8'h6 < length_0 ? _GEN_1967 : _GEN_1807; // @[executor.scala 308:60]
  wire [7:0] _GEN_2128 = 8'h6 < length_0 ? _GEN_1968 : _GEN_1808; // @[executor.scala 308:60]
  wire [7:0] _GEN_2129 = 8'h6 < length_0 ? _GEN_1969 : _GEN_1809; // @[executor.scala 308:60]
  wire [7:0] _GEN_2130 = 8'h6 < length_0 ? _GEN_1970 : _GEN_1810; // @[executor.scala 308:60]
  wire [7:0] _GEN_2131 = 8'h6 < length_0 ? _GEN_1971 : _GEN_1811; // @[executor.scala 308:60]
  wire [7:0] _GEN_2132 = 8'h6 < length_0 ? _GEN_1972 : _GEN_1812; // @[executor.scala 308:60]
  wire [7:0] _GEN_2133 = 8'h6 < length_0 ? _GEN_1973 : _GEN_1813; // @[executor.scala 308:60]
  wire [7:0] _GEN_2134 = 8'h6 < length_0 ? _GEN_1974 : _GEN_1814; // @[executor.scala 308:60]
  wire [7:0] _GEN_2135 = 8'h6 < length_0 ? _GEN_1975 : _GEN_1815; // @[executor.scala 308:60]
  wire [7:0] _GEN_2136 = 8'h6 < length_0 ? _GEN_1976 : _GEN_1816; // @[executor.scala 308:60]
  wire [7:0] _GEN_2137 = 8'h6 < length_0 ? _GEN_1977 : _GEN_1817; // @[executor.scala 308:60]
  wire [7:0] _GEN_2138 = 8'h6 < length_0 ? _GEN_1978 : _GEN_1818; // @[executor.scala 308:60]
  wire [7:0] _GEN_2139 = 8'h6 < length_0 ? _GEN_1979 : _GEN_1819; // @[executor.scala 308:60]
  wire [7:0] _GEN_2140 = 8'h6 < length_0 ? _GEN_1980 : _GEN_1820; // @[executor.scala 308:60]
  wire [7:0] _GEN_2141 = 8'h6 < length_0 ? _GEN_1981 : _GEN_1821; // @[executor.scala 308:60]
  wire [7:0] _GEN_2142 = 8'h6 < length_0 ? _GEN_1982 : _GEN_1822; // @[executor.scala 308:60]
  wire [7:0] _GEN_2143 = 8'h6 < length_0 ? _GEN_1983 : _GEN_1823; // @[executor.scala 308:60]
  wire [7:0] _GEN_2144 = 8'h6 < length_0 ? _GEN_1984 : _GEN_1824; // @[executor.scala 308:60]
  wire [7:0] _GEN_2145 = 8'h6 < length_0 ? _GEN_1985 : _GEN_1825; // @[executor.scala 308:60]
  wire [7:0] _GEN_2146 = 8'h6 < length_0 ? _GEN_1986 : _GEN_1826; // @[executor.scala 308:60]
  wire [7:0] _GEN_2147 = 8'h6 < length_0 ? _GEN_1987 : _GEN_1827; // @[executor.scala 308:60]
  wire [7:0] _GEN_2148 = 8'h6 < length_0 ? _GEN_1988 : _GEN_1828; // @[executor.scala 308:60]
  wire [7:0] _GEN_2149 = 8'h6 < length_0 ? _GEN_1989 : _GEN_1829; // @[executor.scala 308:60]
  wire [7:0] _GEN_2150 = 8'h6 < length_0 ? _GEN_1990 : _GEN_1830; // @[executor.scala 308:60]
  wire [7:0] _GEN_2151 = 8'h6 < length_0 ? _GEN_1991 : _GEN_1831; // @[executor.scala 308:60]
  wire [7:0] _GEN_2152 = 8'h6 < length_0 ? _GEN_1992 : _GEN_1832; // @[executor.scala 308:60]
  wire [7:0] _GEN_2153 = 8'h6 < length_0 ? _GEN_1993 : _GEN_1833; // @[executor.scala 308:60]
  wire [7:0] _GEN_2154 = 8'h6 < length_0 ? _GEN_1994 : _GEN_1834; // @[executor.scala 308:60]
  wire [7:0] _GEN_2155 = 8'h6 < length_0 ? _GEN_1995 : _GEN_1835; // @[executor.scala 308:60]
  wire [7:0] _GEN_2156 = 8'h6 < length_0 ? _GEN_1996 : _GEN_1836; // @[executor.scala 308:60]
  wire [7:0] _GEN_2157 = 8'h6 < length_0 ? _GEN_1997 : _GEN_1837; // @[executor.scala 308:60]
  wire [7:0] _GEN_2158 = 8'h6 < length_0 ? _GEN_1998 : _GEN_1838; // @[executor.scala 308:60]
  wire [7:0] _GEN_2159 = 8'h6 < length_0 ? _GEN_1999 : _GEN_1839; // @[executor.scala 308:60]
  wire [7:0] _GEN_2160 = 8'h6 < length_0 ? _GEN_2000 : _GEN_1840; // @[executor.scala 308:60]
  wire [7:0] _GEN_2161 = 8'h6 < length_0 ? _GEN_2001 : _GEN_1841; // @[executor.scala 308:60]
  wire [7:0] _GEN_2162 = 8'h6 < length_0 ? _GEN_2002 : _GEN_1842; // @[executor.scala 308:60]
  wire [7:0] _GEN_2163 = 8'h6 < length_0 ? _GEN_2003 : _GEN_1843; // @[executor.scala 308:60]
  wire [7:0] _GEN_2164 = 8'h6 < length_0 ? _GEN_2004 : _GEN_1844; // @[executor.scala 308:60]
  wire [7:0] _GEN_2165 = 8'h6 < length_0 ? _GEN_2005 : _GEN_1845; // @[executor.scala 308:60]
  wire [7:0] _GEN_2166 = 8'h6 < length_0 ? _GEN_2006 : _GEN_1846; // @[executor.scala 308:60]
  wire [7:0] _GEN_2167 = 8'h6 < length_0 ? _GEN_2007 : _GEN_1847; // @[executor.scala 308:60]
  wire [7:0] _GEN_2168 = 8'h6 < length_0 ? _GEN_2008 : _GEN_1848; // @[executor.scala 308:60]
  wire [7:0] _GEN_2169 = 8'h6 < length_0 ? _GEN_2009 : _GEN_1849; // @[executor.scala 308:60]
  wire [7:0] _GEN_2170 = 8'h6 < length_0 ? _GEN_2010 : _GEN_1850; // @[executor.scala 308:60]
  wire [7:0] _GEN_2171 = 8'h6 < length_0 ? _GEN_2011 : _GEN_1851; // @[executor.scala 308:60]
  wire [7:0] _GEN_2172 = 8'h6 < length_0 ? _GEN_2012 : _GEN_1852; // @[executor.scala 308:60]
  wire [7:0] _GEN_2173 = 8'h6 < length_0 ? _GEN_2013 : _GEN_1853; // @[executor.scala 308:60]
  wire [7:0] _GEN_2174 = 8'h6 < length_0 ? _GEN_2014 : _GEN_1854; // @[executor.scala 308:60]
  wire [7:0] _GEN_2175 = 8'h6 < length_0 ? _GEN_2015 : _GEN_1855; // @[executor.scala 308:60]
  wire [7:0] _GEN_2176 = 8'h6 < length_0 ? _GEN_2016 : _GEN_1856; // @[executor.scala 308:60]
  wire [7:0] _GEN_2177 = 8'h6 < length_0 ? _GEN_2017 : _GEN_1857; // @[executor.scala 308:60]
  wire [7:0] _GEN_2178 = 8'h6 < length_0 ? _GEN_2018 : _GEN_1858; // @[executor.scala 308:60]
  wire [7:0] _GEN_2179 = 8'h6 < length_0 ? _GEN_2019 : _GEN_1859; // @[executor.scala 308:60]
  wire [7:0] _GEN_2180 = 8'h6 < length_0 ? _GEN_2020 : _GEN_1860; // @[executor.scala 308:60]
  wire [7:0] _GEN_2181 = 8'h6 < length_0 ? _GEN_2021 : _GEN_1861; // @[executor.scala 308:60]
  wire [7:0] _GEN_2182 = 8'h6 < length_0 ? _GEN_2022 : _GEN_1862; // @[executor.scala 308:60]
  wire [7:0] _GEN_2183 = 8'h6 < length_0 ? _GEN_2023 : _GEN_1863; // @[executor.scala 308:60]
  wire [7:0] _GEN_2184 = 8'h6 < length_0 ? _GEN_2024 : _GEN_1864; // @[executor.scala 308:60]
  wire [7:0] _GEN_2185 = 8'h6 < length_0 ? _GEN_2025 : _GEN_1865; // @[executor.scala 308:60]
  wire [7:0] _GEN_2186 = 8'h6 < length_0 ? _GEN_2026 : _GEN_1866; // @[executor.scala 308:60]
  wire [7:0] _GEN_2187 = 8'h6 < length_0 ? _GEN_2027 : _GEN_1867; // @[executor.scala 308:60]
  wire [7:0] _GEN_2188 = 8'h6 < length_0 ? _GEN_2028 : _GEN_1868; // @[executor.scala 308:60]
  wire [7:0] _GEN_2189 = 8'h6 < length_0 ? _GEN_2029 : _GEN_1869; // @[executor.scala 308:60]
  wire [7:0] _GEN_2190 = 8'h6 < length_0 ? _GEN_2030 : _GEN_1870; // @[executor.scala 308:60]
  wire [7:0] _GEN_2191 = 8'h6 < length_0 ? _GEN_2031 : _GEN_1871; // @[executor.scala 308:60]
  wire [7:0] _GEN_2192 = 8'h6 < length_0 ? _GEN_2032 : _GEN_1872; // @[executor.scala 308:60]
  wire [7:0] _GEN_2193 = 8'h6 < length_0 ? _GEN_2033 : _GEN_1873; // @[executor.scala 308:60]
  wire [7:0] _GEN_2194 = 8'h6 < length_0 ? _GEN_2034 : _GEN_1874; // @[executor.scala 308:60]
  wire [7:0] _GEN_2195 = 8'h6 < length_0 ? _GEN_2035 : _GEN_1875; // @[executor.scala 308:60]
  wire [7:0] _GEN_2196 = 8'h6 < length_0 ? _GEN_2036 : _GEN_1876; // @[executor.scala 308:60]
  wire [7:0] _GEN_2197 = 8'h6 < length_0 ? _GEN_2037 : _GEN_1877; // @[executor.scala 308:60]
  wire [7:0] _GEN_2198 = 8'h6 < length_0 ? _GEN_2038 : _GEN_1878; // @[executor.scala 308:60]
  wire [7:0] _GEN_2199 = 8'h6 < length_0 ? _GEN_2039 : _GEN_1879; // @[executor.scala 308:60]
  wire [7:0] _GEN_2200 = 8'h6 < length_0 ? _GEN_2040 : _GEN_1880; // @[executor.scala 308:60]
  wire [7:0] _GEN_2201 = 8'h6 < length_0 ? _GEN_2041 : _GEN_1881; // @[executor.scala 308:60]
  wire [7:0] _GEN_2202 = 8'h6 < length_0 ? _GEN_2042 : _GEN_1882; // @[executor.scala 308:60]
  wire [7:0] _GEN_2203 = 8'h6 < length_0 ? _GEN_2043 : _GEN_1883; // @[executor.scala 308:60]
  wire [7:0] _GEN_2204 = 8'h6 < length_0 ? _GEN_2044 : _GEN_1884; // @[executor.scala 308:60]
  wire [7:0] _GEN_2205 = 8'h6 < length_0 ? _GEN_2045 : _GEN_1885; // @[executor.scala 308:60]
  wire [7:0] _GEN_2206 = 8'h6 < length_0 ? _GEN_2046 : _GEN_1886; // @[executor.scala 308:60]
  wire [7:0] _GEN_2207 = 8'h6 < length_0 ? _GEN_2047 : _GEN_1887; // @[executor.scala 308:60]
  wire [7:0] _GEN_2208 = 8'h6 < length_0 ? _GEN_2048 : _GEN_1888; // @[executor.scala 308:60]
  wire [7:0] _GEN_2209 = 8'h6 < length_0 ? _GEN_2049 : _GEN_1889; // @[executor.scala 308:60]
  wire [7:0] _GEN_2210 = 8'h6 < length_0 ? _GEN_2050 : _GEN_1890; // @[executor.scala 308:60]
  wire [7:0] _GEN_2211 = 8'h6 < length_0 ? _GEN_2051 : _GEN_1891; // @[executor.scala 308:60]
  wire [7:0] _GEN_2212 = 8'h6 < length_0 ? _GEN_2052 : _GEN_1892; // @[executor.scala 308:60]
  wire [7:0] _GEN_2213 = 8'h6 < length_0 ? _GEN_2053 : _GEN_1893; // @[executor.scala 308:60]
  wire [7:0] _GEN_2214 = 8'h6 < length_0 ? _GEN_2054 : _GEN_1894; // @[executor.scala 308:60]
  wire [7:0] _GEN_2215 = 8'h6 < length_0 ? _GEN_2055 : _GEN_1895; // @[executor.scala 308:60]
  wire [7:0] _GEN_2216 = 8'h6 < length_0 ? _GEN_2056 : _GEN_1896; // @[executor.scala 308:60]
  wire [7:0] _GEN_2217 = 8'h6 < length_0 ? _GEN_2057 : _GEN_1897; // @[executor.scala 308:60]
  wire [7:0] _GEN_2218 = 8'h6 < length_0 ? _GEN_2058 : _GEN_1898; // @[executor.scala 308:60]
  wire [7:0] _GEN_2219 = 8'h6 < length_0 ? _GEN_2059 : _GEN_1899; // @[executor.scala 308:60]
  wire [7:0] _GEN_2220 = 8'h6 < length_0 ? _GEN_2060 : _GEN_1900; // @[executor.scala 308:60]
  wire [7:0] _GEN_2221 = 8'h6 < length_0 ? _GEN_2061 : _GEN_1901; // @[executor.scala 308:60]
  wire [7:0] _GEN_2222 = 8'h6 < length_0 ? _GEN_2062 : _GEN_1902; // @[executor.scala 308:60]
  wire [7:0] _GEN_2223 = 8'h6 < length_0 ? _GEN_2063 : _GEN_1903; // @[executor.scala 308:60]
  wire [7:0] _GEN_2224 = 8'h6 < length_0 ? _GEN_2064 : _GEN_1904; // @[executor.scala 308:60]
  wire [7:0] _GEN_2225 = 8'h6 < length_0 ? _GEN_2065 : _GEN_1905; // @[executor.scala 308:60]
  wire [7:0] _GEN_2226 = 8'h6 < length_0 ? _GEN_2066 : _GEN_1906; // @[executor.scala 308:60]
  wire [7:0] _GEN_2227 = 8'h6 < length_0 ? _GEN_2067 : _GEN_1907; // @[executor.scala 308:60]
  wire [7:0] _GEN_2228 = 8'h6 < length_0 ? _GEN_2068 : _GEN_1908; // @[executor.scala 308:60]
  wire [7:0] _GEN_2229 = 8'h6 < length_0 ? _GEN_2069 : _GEN_1909; // @[executor.scala 308:60]
  wire [7:0] _GEN_2230 = 8'h6 < length_0 ? _GEN_2070 : _GEN_1910; // @[executor.scala 308:60]
  wire [7:0] _GEN_2231 = 8'h6 < length_0 ? _GEN_2071 : _GEN_1911; // @[executor.scala 308:60]
  wire [7:0] _GEN_2232 = 8'h6 < length_0 ? _GEN_2072 : _GEN_1912; // @[executor.scala 308:60]
  wire [7:0] _GEN_2233 = 8'h6 < length_0 ? _GEN_2073 : _GEN_1913; // @[executor.scala 308:60]
  wire [7:0] _GEN_2234 = 8'h6 < length_0 ? _GEN_2074 : _GEN_1914; // @[executor.scala 308:60]
  wire [7:0] _GEN_2235 = 8'h6 < length_0 ? _GEN_2075 : _GEN_1915; // @[executor.scala 308:60]
  wire [7:0] _GEN_2236 = 8'h6 < length_0 ? _GEN_2076 : _GEN_1916; // @[executor.scala 308:60]
  wire [7:0] _GEN_2237 = 8'h6 < length_0 ? _GEN_2077 : _GEN_1917; // @[executor.scala 308:60]
  wire [7:0] _GEN_2238 = 8'h6 < length_0 ? _GEN_2078 : _GEN_1918; // @[executor.scala 308:60]
  wire [7:0] _GEN_2239 = 8'h6 < length_0 ? _GEN_2079 : _GEN_1919; // @[executor.scala 308:60]
  wire [7:0] field_byte_7 = field_0[7:0]; // @[executor.scala 305:57]
  wire [7:0] total_offset_7 = offset_0 + 8'h7; // @[executor.scala 307:57]
  wire [7:0] _GEN_2240 = 8'h0 == total_offset_7 ? field_byte_7 : _GEN_2080; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2241 = 8'h1 == total_offset_7 ? field_byte_7 : _GEN_2081; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2242 = 8'h2 == total_offset_7 ? field_byte_7 : _GEN_2082; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2243 = 8'h3 == total_offset_7 ? field_byte_7 : _GEN_2083; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2244 = 8'h4 == total_offset_7 ? field_byte_7 : _GEN_2084; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2245 = 8'h5 == total_offset_7 ? field_byte_7 : _GEN_2085; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2246 = 8'h6 == total_offset_7 ? field_byte_7 : _GEN_2086; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2247 = 8'h7 == total_offset_7 ? field_byte_7 : _GEN_2087; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2248 = 8'h8 == total_offset_7 ? field_byte_7 : _GEN_2088; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2249 = 8'h9 == total_offset_7 ? field_byte_7 : _GEN_2089; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2250 = 8'ha == total_offset_7 ? field_byte_7 : _GEN_2090; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2251 = 8'hb == total_offset_7 ? field_byte_7 : _GEN_2091; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2252 = 8'hc == total_offset_7 ? field_byte_7 : _GEN_2092; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2253 = 8'hd == total_offset_7 ? field_byte_7 : _GEN_2093; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2254 = 8'he == total_offset_7 ? field_byte_7 : _GEN_2094; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2255 = 8'hf == total_offset_7 ? field_byte_7 : _GEN_2095; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2256 = 8'h10 == total_offset_7 ? field_byte_7 : _GEN_2096; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2257 = 8'h11 == total_offset_7 ? field_byte_7 : _GEN_2097; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2258 = 8'h12 == total_offset_7 ? field_byte_7 : _GEN_2098; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2259 = 8'h13 == total_offset_7 ? field_byte_7 : _GEN_2099; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2260 = 8'h14 == total_offset_7 ? field_byte_7 : _GEN_2100; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2261 = 8'h15 == total_offset_7 ? field_byte_7 : _GEN_2101; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2262 = 8'h16 == total_offset_7 ? field_byte_7 : _GEN_2102; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2263 = 8'h17 == total_offset_7 ? field_byte_7 : _GEN_2103; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2264 = 8'h18 == total_offset_7 ? field_byte_7 : _GEN_2104; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2265 = 8'h19 == total_offset_7 ? field_byte_7 : _GEN_2105; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2266 = 8'h1a == total_offset_7 ? field_byte_7 : _GEN_2106; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2267 = 8'h1b == total_offset_7 ? field_byte_7 : _GEN_2107; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2268 = 8'h1c == total_offset_7 ? field_byte_7 : _GEN_2108; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2269 = 8'h1d == total_offset_7 ? field_byte_7 : _GEN_2109; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2270 = 8'h1e == total_offset_7 ? field_byte_7 : _GEN_2110; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2271 = 8'h1f == total_offset_7 ? field_byte_7 : _GEN_2111; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2272 = 8'h20 == total_offset_7 ? field_byte_7 : _GEN_2112; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2273 = 8'h21 == total_offset_7 ? field_byte_7 : _GEN_2113; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2274 = 8'h22 == total_offset_7 ? field_byte_7 : _GEN_2114; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2275 = 8'h23 == total_offset_7 ? field_byte_7 : _GEN_2115; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2276 = 8'h24 == total_offset_7 ? field_byte_7 : _GEN_2116; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2277 = 8'h25 == total_offset_7 ? field_byte_7 : _GEN_2117; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2278 = 8'h26 == total_offset_7 ? field_byte_7 : _GEN_2118; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2279 = 8'h27 == total_offset_7 ? field_byte_7 : _GEN_2119; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2280 = 8'h28 == total_offset_7 ? field_byte_7 : _GEN_2120; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2281 = 8'h29 == total_offset_7 ? field_byte_7 : _GEN_2121; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2282 = 8'h2a == total_offset_7 ? field_byte_7 : _GEN_2122; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2283 = 8'h2b == total_offset_7 ? field_byte_7 : _GEN_2123; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2284 = 8'h2c == total_offset_7 ? field_byte_7 : _GEN_2124; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2285 = 8'h2d == total_offset_7 ? field_byte_7 : _GEN_2125; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2286 = 8'h2e == total_offset_7 ? field_byte_7 : _GEN_2126; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2287 = 8'h2f == total_offset_7 ? field_byte_7 : _GEN_2127; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2288 = 8'h30 == total_offset_7 ? field_byte_7 : _GEN_2128; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2289 = 8'h31 == total_offset_7 ? field_byte_7 : _GEN_2129; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2290 = 8'h32 == total_offset_7 ? field_byte_7 : _GEN_2130; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2291 = 8'h33 == total_offset_7 ? field_byte_7 : _GEN_2131; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2292 = 8'h34 == total_offset_7 ? field_byte_7 : _GEN_2132; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2293 = 8'h35 == total_offset_7 ? field_byte_7 : _GEN_2133; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2294 = 8'h36 == total_offset_7 ? field_byte_7 : _GEN_2134; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2295 = 8'h37 == total_offset_7 ? field_byte_7 : _GEN_2135; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2296 = 8'h38 == total_offset_7 ? field_byte_7 : _GEN_2136; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2297 = 8'h39 == total_offset_7 ? field_byte_7 : _GEN_2137; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2298 = 8'h3a == total_offset_7 ? field_byte_7 : _GEN_2138; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2299 = 8'h3b == total_offset_7 ? field_byte_7 : _GEN_2139; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2300 = 8'h3c == total_offset_7 ? field_byte_7 : _GEN_2140; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2301 = 8'h3d == total_offset_7 ? field_byte_7 : _GEN_2141; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2302 = 8'h3e == total_offset_7 ? field_byte_7 : _GEN_2142; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2303 = 8'h3f == total_offset_7 ? field_byte_7 : _GEN_2143; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2304 = 8'h40 == total_offset_7 ? field_byte_7 : _GEN_2144; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2305 = 8'h41 == total_offset_7 ? field_byte_7 : _GEN_2145; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2306 = 8'h42 == total_offset_7 ? field_byte_7 : _GEN_2146; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2307 = 8'h43 == total_offset_7 ? field_byte_7 : _GEN_2147; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2308 = 8'h44 == total_offset_7 ? field_byte_7 : _GEN_2148; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2309 = 8'h45 == total_offset_7 ? field_byte_7 : _GEN_2149; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2310 = 8'h46 == total_offset_7 ? field_byte_7 : _GEN_2150; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2311 = 8'h47 == total_offset_7 ? field_byte_7 : _GEN_2151; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2312 = 8'h48 == total_offset_7 ? field_byte_7 : _GEN_2152; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2313 = 8'h49 == total_offset_7 ? field_byte_7 : _GEN_2153; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2314 = 8'h4a == total_offset_7 ? field_byte_7 : _GEN_2154; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2315 = 8'h4b == total_offset_7 ? field_byte_7 : _GEN_2155; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2316 = 8'h4c == total_offset_7 ? field_byte_7 : _GEN_2156; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2317 = 8'h4d == total_offset_7 ? field_byte_7 : _GEN_2157; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2318 = 8'h4e == total_offset_7 ? field_byte_7 : _GEN_2158; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2319 = 8'h4f == total_offset_7 ? field_byte_7 : _GEN_2159; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2320 = 8'h50 == total_offset_7 ? field_byte_7 : _GEN_2160; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2321 = 8'h51 == total_offset_7 ? field_byte_7 : _GEN_2161; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2322 = 8'h52 == total_offset_7 ? field_byte_7 : _GEN_2162; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2323 = 8'h53 == total_offset_7 ? field_byte_7 : _GEN_2163; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2324 = 8'h54 == total_offset_7 ? field_byte_7 : _GEN_2164; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2325 = 8'h55 == total_offset_7 ? field_byte_7 : _GEN_2165; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2326 = 8'h56 == total_offset_7 ? field_byte_7 : _GEN_2166; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2327 = 8'h57 == total_offset_7 ? field_byte_7 : _GEN_2167; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2328 = 8'h58 == total_offset_7 ? field_byte_7 : _GEN_2168; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2329 = 8'h59 == total_offset_7 ? field_byte_7 : _GEN_2169; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2330 = 8'h5a == total_offset_7 ? field_byte_7 : _GEN_2170; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2331 = 8'h5b == total_offset_7 ? field_byte_7 : _GEN_2171; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2332 = 8'h5c == total_offset_7 ? field_byte_7 : _GEN_2172; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2333 = 8'h5d == total_offset_7 ? field_byte_7 : _GEN_2173; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2334 = 8'h5e == total_offset_7 ? field_byte_7 : _GEN_2174; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2335 = 8'h5f == total_offset_7 ? field_byte_7 : _GEN_2175; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2336 = 8'h60 == total_offset_7 ? field_byte_7 : _GEN_2176; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2337 = 8'h61 == total_offset_7 ? field_byte_7 : _GEN_2177; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2338 = 8'h62 == total_offset_7 ? field_byte_7 : _GEN_2178; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2339 = 8'h63 == total_offset_7 ? field_byte_7 : _GEN_2179; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2340 = 8'h64 == total_offset_7 ? field_byte_7 : _GEN_2180; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2341 = 8'h65 == total_offset_7 ? field_byte_7 : _GEN_2181; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2342 = 8'h66 == total_offset_7 ? field_byte_7 : _GEN_2182; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2343 = 8'h67 == total_offset_7 ? field_byte_7 : _GEN_2183; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2344 = 8'h68 == total_offset_7 ? field_byte_7 : _GEN_2184; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2345 = 8'h69 == total_offset_7 ? field_byte_7 : _GEN_2185; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2346 = 8'h6a == total_offset_7 ? field_byte_7 : _GEN_2186; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2347 = 8'h6b == total_offset_7 ? field_byte_7 : _GEN_2187; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2348 = 8'h6c == total_offset_7 ? field_byte_7 : _GEN_2188; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2349 = 8'h6d == total_offset_7 ? field_byte_7 : _GEN_2189; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2350 = 8'h6e == total_offset_7 ? field_byte_7 : _GEN_2190; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2351 = 8'h6f == total_offset_7 ? field_byte_7 : _GEN_2191; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2352 = 8'h70 == total_offset_7 ? field_byte_7 : _GEN_2192; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2353 = 8'h71 == total_offset_7 ? field_byte_7 : _GEN_2193; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2354 = 8'h72 == total_offset_7 ? field_byte_7 : _GEN_2194; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2355 = 8'h73 == total_offset_7 ? field_byte_7 : _GEN_2195; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2356 = 8'h74 == total_offset_7 ? field_byte_7 : _GEN_2196; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2357 = 8'h75 == total_offset_7 ? field_byte_7 : _GEN_2197; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2358 = 8'h76 == total_offset_7 ? field_byte_7 : _GEN_2198; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2359 = 8'h77 == total_offset_7 ? field_byte_7 : _GEN_2199; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2360 = 8'h78 == total_offset_7 ? field_byte_7 : _GEN_2200; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2361 = 8'h79 == total_offset_7 ? field_byte_7 : _GEN_2201; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2362 = 8'h7a == total_offset_7 ? field_byte_7 : _GEN_2202; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2363 = 8'h7b == total_offset_7 ? field_byte_7 : _GEN_2203; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2364 = 8'h7c == total_offset_7 ? field_byte_7 : _GEN_2204; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2365 = 8'h7d == total_offset_7 ? field_byte_7 : _GEN_2205; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2366 = 8'h7e == total_offset_7 ? field_byte_7 : _GEN_2206; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2367 = 8'h7f == total_offset_7 ? field_byte_7 : _GEN_2207; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2368 = 8'h80 == total_offset_7 ? field_byte_7 : _GEN_2208; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2369 = 8'h81 == total_offset_7 ? field_byte_7 : _GEN_2209; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2370 = 8'h82 == total_offset_7 ? field_byte_7 : _GEN_2210; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2371 = 8'h83 == total_offset_7 ? field_byte_7 : _GEN_2211; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2372 = 8'h84 == total_offset_7 ? field_byte_7 : _GEN_2212; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2373 = 8'h85 == total_offset_7 ? field_byte_7 : _GEN_2213; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2374 = 8'h86 == total_offset_7 ? field_byte_7 : _GEN_2214; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2375 = 8'h87 == total_offset_7 ? field_byte_7 : _GEN_2215; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2376 = 8'h88 == total_offset_7 ? field_byte_7 : _GEN_2216; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2377 = 8'h89 == total_offset_7 ? field_byte_7 : _GEN_2217; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2378 = 8'h8a == total_offset_7 ? field_byte_7 : _GEN_2218; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2379 = 8'h8b == total_offset_7 ? field_byte_7 : _GEN_2219; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2380 = 8'h8c == total_offset_7 ? field_byte_7 : _GEN_2220; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2381 = 8'h8d == total_offset_7 ? field_byte_7 : _GEN_2221; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2382 = 8'h8e == total_offset_7 ? field_byte_7 : _GEN_2222; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2383 = 8'h8f == total_offset_7 ? field_byte_7 : _GEN_2223; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2384 = 8'h90 == total_offset_7 ? field_byte_7 : _GEN_2224; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2385 = 8'h91 == total_offset_7 ? field_byte_7 : _GEN_2225; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2386 = 8'h92 == total_offset_7 ? field_byte_7 : _GEN_2226; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2387 = 8'h93 == total_offset_7 ? field_byte_7 : _GEN_2227; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2388 = 8'h94 == total_offset_7 ? field_byte_7 : _GEN_2228; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2389 = 8'h95 == total_offset_7 ? field_byte_7 : _GEN_2229; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2390 = 8'h96 == total_offset_7 ? field_byte_7 : _GEN_2230; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2391 = 8'h97 == total_offset_7 ? field_byte_7 : _GEN_2231; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2392 = 8'h98 == total_offset_7 ? field_byte_7 : _GEN_2232; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2393 = 8'h99 == total_offset_7 ? field_byte_7 : _GEN_2233; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2394 = 8'h9a == total_offset_7 ? field_byte_7 : _GEN_2234; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2395 = 8'h9b == total_offset_7 ? field_byte_7 : _GEN_2235; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2396 = 8'h9c == total_offset_7 ? field_byte_7 : _GEN_2236; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2397 = 8'h9d == total_offset_7 ? field_byte_7 : _GEN_2237; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2398 = 8'h9e == total_offset_7 ? field_byte_7 : _GEN_2238; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2399 = 8'h9f == total_offset_7 ? field_byte_7 : _GEN_2239; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2400 = 8'h7 < length_0 ? _GEN_2240 : _GEN_2080; // @[executor.scala 308:60]
  wire [7:0] _GEN_2401 = 8'h7 < length_0 ? _GEN_2241 : _GEN_2081; // @[executor.scala 308:60]
  wire [7:0] _GEN_2402 = 8'h7 < length_0 ? _GEN_2242 : _GEN_2082; // @[executor.scala 308:60]
  wire [7:0] _GEN_2403 = 8'h7 < length_0 ? _GEN_2243 : _GEN_2083; // @[executor.scala 308:60]
  wire [7:0] _GEN_2404 = 8'h7 < length_0 ? _GEN_2244 : _GEN_2084; // @[executor.scala 308:60]
  wire [7:0] _GEN_2405 = 8'h7 < length_0 ? _GEN_2245 : _GEN_2085; // @[executor.scala 308:60]
  wire [7:0] _GEN_2406 = 8'h7 < length_0 ? _GEN_2246 : _GEN_2086; // @[executor.scala 308:60]
  wire [7:0] _GEN_2407 = 8'h7 < length_0 ? _GEN_2247 : _GEN_2087; // @[executor.scala 308:60]
  wire [7:0] _GEN_2408 = 8'h7 < length_0 ? _GEN_2248 : _GEN_2088; // @[executor.scala 308:60]
  wire [7:0] _GEN_2409 = 8'h7 < length_0 ? _GEN_2249 : _GEN_2089; // @[executor.scala 308:60]
  wire [7:0] _GEN_2410 = 8'h7 < length_0 ? _GEN_2250 : _GEN_2090; // @[executor.scala 308:60]
  wire [7:0] _GEN_2411 = 8'h7 < length_0 ? _GEN_2251 : _GEN_2091; // @[executor.scala 308:60]
  wire [7:0] _GEN_2412 = 8'h7 < length_0 ? _GEN_2252 : _GEN_2092; // @[executor.scala 308:60]
  wire [7:0] _GEN_2413 = 8'h7 < length_0 ? _GEN_2253 : _GEN_2093; // @[executor.scala 308:60]
  wire [7:0] _GEN_2414 = 8'h7 < length_0 ? _GEN_2254 : _GEN_2094; // @[executor.scala 308:60]
  wire [7:0] _GEN_2415 = 8'h7 < length_0 ? _GEN_2255 : _GEN_2095; // @[executor.scala 308:60]
  wire [7:0] _GEN_2416 = 8'h7 < length_0 ? _GEN_2256 : _GEN_2096; // @[executor.scala 308:60]
  wire [7:0] _GEN_2417 = 8'h7 < length_0 ? _GEN_2257 : _GEN_2097; // @[executor.scala 308:60]
  wire [7:0] _GEN_2418 = 8'h7 < length_0 ? _GEN_2258 : _GEN_2098; // @[executor.scala 308:60]
  wire [7:0] _GEN_2419 = 8'h7 < length_0 ? _GEN_2259 : _GEN_2099; // @[executor.scala 308:60]
  wire [7:0] _GEN_2420 = 8'h7 < length_0 ? _GEN_2260 : _GEN_2100; // @[executor.scala 308:60]
  wire [7:0] _GEN_2421 = 8'h7 < length_0 ? _GEN_2261 : _GEN_2101; // @[executor.scala 308:60]
  wire [7:0] _GEN_2422 = 8'h7 < length_0 ? _GEN_2262 : _GEN_2102; // @[executor.scala 308:60]
  wire [7:0] _GEN_2423 = 8'h7 < length_0 ? _GEN_2263 : _GEN_2103; // @[executor.scala 308:60]
  wire [7:0] _GEN_2424 = 8'h7 < length_0 ? _GEN_2264 : _GEN_2104; // @[executor.scala 308:60]
  wire [7:0] _GEN_2425 = 8'h7 < length_0 ? _GEN_2265 : _GEN_2105; // @[executor.scala 308:60]
  wire [7:0] _GEN_2426 = 8'h7 < length_0 ? _GEN_2266 : _GEN_2106; // @[executor.scala 308:60]
  wire [7:0] _GEN_2427 = 8'h7 < length_0 ? _GEN_2267 : _GEN_2107; // @[executor.scala 308:60]
  wire [7:0] _GEN_2428 = 8'h7 < length_0 ? _GEN_2268 : _GEN_2108; // @[executor.scala 308:60]
  wire [7:0] _GEN_2429 = 8'h7 < length_0 ? _GEN_2269 : _GEN_2109; // @[executor.scala 308:60]
  wire [7:0] _GEN_2430 = 8'h7 < length_0 ? _GEN_2270 : _GEN_2110; // @[executor.scala 308:60]
  wire [7:0] _GEN_2431 = 8'h7 < length_0 ? _GEN_2271 : _GEN_2111; // @[executor.scala 308:60]
  wire [7:0] _GEN_2432 = 8'h7 < length_0 ? _GEN_2272 : _GEN_2112; // @[executor.scala 308:60]
  wire [7:0] _GEN_2433 = 8'h7 < length_0 ? _GEN_2273 : _GEN_2113; // @[executor.scala 308:60]
  wire [7:0] _GEN_2434 = 8'h7 < length_0 ? _GEN_2274 : _GEN_2114; // @[executor.scala 308:60]
  wire [7:0] _GEN_2435 = 8'h7 < length_0 ? _GEN_2275 : _GEN_2115; // @[executor.scala 308:60]
  wire [7:0] _GEN_2436 = 8'h7 < length_0 ? _GEN_2276 : _GEN_2116; // @[executor.scala 308:60]
  wire [7:0] _GEN_2437 = 8'h7 < length_0 ? _GEN_2277 : _GEN_2117; // @[executor.scala 308:60]
  wire [7:0] _GEN_2438 = 8'h7 < length_0 ? _GEN_2278 : _GEN_2118; // @[executor.scala 308:60]
  wire [7:0] _GEN_2439 = 8'h7 < length_0 ? _GEN_2279 : _GEN_2119; // @[executor.scala 308:60]
  wire [7:0] _GEN_2440 = 8'h7 < length_0 ? _GEN_2280 : _GEN_2120; // @[executor.scala 308:60]
  wire [7:0] _GEN_2441 = 8'h7 < length_0 ? _GEN_2281 : _GEN_2121; // @[executor.scala 308:60]
  wire [7:0] _GEN_2442 = 8'h7 < length_0 ? _GEN_2282 : _GEN_2122; // @[executor.scala 308:60]
  wire [7:0] _GEN_2443 = 8'h7 < length_0 ? _GEN_2283 : _GEN_2123; // @[executor.scala 308:60]
  wire [7:0] _GEN_2444 = 8'h7 < length_0 ? _GEN_2284 : _GEN_2124; // @[executor.scala 308:60]
  wire [7:0] _GEN_2445 = 8'h7 < length_0 ? _GEN_2285 : _GEN_2125; // @[executor.scala 308:60]
  wire [7:0] _GEN_2446 = 8'h7 < length_0 ? _GEN_2286 : _GEN_2126; // @[executor.scala 308:60]
  wire [7:0] _GEN_2447 = 8'h7 < length_0 ? _GEN_2287 : _GEN_2127; // @[executor.scala 308:60]
  wire [7:0] _GEN_2448 = 8'h7 < length_0 ? _GEN_2288 : _GEN_2128; // @[executor.scala 308:60]
  wire [7:0] _GEN_2449 = 8'h7 < length_0 ? _GEN_2289 : _GEN_2129; // @[executor.scala 308:60]
  wire [7:0] _GEN_2450 = 8'h7 < length_0 ? _GEN_2290 : _GEN_2130; // @[executor.scala 308:60]
  wire [7:0] _GEN_2451 = 8'h7 < length_0 ? _GEN_2291 : _GEN_2131; // @[executor.scala 308:60]
  wire [7:0] _GEN_2452 = 8'h7 < length_0 ? _GEN_2292 : _GEN_2132; // @[executor.scala 308:60]
  wire [7:0] _GEN_2453 = 8'h7 < length_0 ? _GEN_2293 : _GEN_2133; // @[executor.scala 308:60]
  wire [7:0] _GEN_2454 = 8'h7 < length_0 ? _GEN_2294 : _GEN_2134; // @[executor.scala 308:60]
  wire [7:0] _GEN_2455 = 8'h7 < length_0 ? _GEN_2295 : _GEN_2135; // @[executor.scala 308:60]
  wire [7:0] _GEN_2456 = 8'h7 < length_0 ? _GEN_2296 : _GEN_2136; // @[executor.scala 308:60]
  wire [7:0] _GEN_2457 = 8'h7 < length_0 ? _GEN_2297 : _GEN_2137; // @[executor.scala 308:60]
  wire [7:0] _GEN_2458 = 8'h7 < length_0 ? _GEN_2298 : _GEN_2138; // @[executor.scala 308:60]
  wire [7:0] _GEN_2459 = 8'h7 < length_0 ? _GEN_2299 : _GEN_2139; // @[executor.scala 308:60]
  wire [7:0] _GEN_2460 = 8'h7 < length_0 ? _GEN_2300 : _GEN_2140; // @[executor.scala 308:60]
  wire [7:0] _GEN_2461 = 8'h7 < length_0 ? _GEN_2301 : _GEN_2141; // @[executor.scala 308:60]
  wire [7:0] _GEN_2462 = 8'h7 < length_0 ? _GEN_2302 : _GEN_2142; // @[executor.scala 308:60]
  wire [7:0] _GEN_2463 = 8'h7 < length_0 ? _GEN_2303 : _GEN_2143; // @[executor.scala 308:60]
  wire [7:0] _GEN_2464 = 8'h7 < length_0 ? _GEN_2304 : _GEN_2144; // @[executor.scala 308:60]
  wire [7:0] _GEN_2465 = 8'h7 < length_0 ? _GEN_2305 : _GEN_2145; // @[executor.scala 308:60]
  wire [7:0] _GEN_2466 = 8'h7 < length_0 ? _GEN_2306 : _GEN_2146; // @[executor.scala 308:60]
  wire [7:0] _GEN_2467 = 8'h7 < length_0 ? _GEN_2307 : _GEN_2147; // @[executor.scala 308:60]
  wire [7:0] _GEN_2468 = 8'h7 < length_0 ? _GEN_2308 : _GEN_2148; // @[executor.scala 308:60]
  wire [7:0] _GEN_2469 = 8'h7 < length_0 ? _GEN_2309 : _GEN_2149; // @[executor.scala 308:60]
  wire [7:0] _GEN_2470 = 8'h7 < length_0 ? _GEN_2310 : _GEN_2150; // @[executor.scala 308:60]
  wire [7:0] _GEN_2471 = 8'h7 < length_0 ? _GEN_2311 : _GEN_2151; // @[executor.scala 308:60]
  wire [7:0] _GEN_2472 = 8'h7 < length_0 ? _GEN_2312 : _GEN_2152; // @[executor.scala 308:60]
  wire [7:0] _GEN_2473 = 8'h7 < length_0 ? _GEN_2313 : _GEN_2153; // @[executor.scala 308:60]
  wire [7:0] _GEN_2474 = 8'h7 < length_0 ? _GEN_2314 : _GEN_2154; // @[executor.scala 308:60]
  wire [7:0] _GEN_2475 = 8'h7 < length_0 ? _GEN_2315 : _GEN_2155; // @[executor.scala 308:60]
  wire [7:0] _GEN_2476 = 8'h7 < length_0 ? _GEN_2316 : _GEN_2156; // @[executor.scala 308:60]
  wire [7:0] _GEN_2477 = 8'h7 < length_0 ? _GEN_2317 : _GEN_2157; // @[executor.scala 308:60]
  wire [7:0] _GEN_2478 = 8'h7 < length_0 ? _GEN_2318 : _GEN_2158; // @[executor.scala 308:60]
  wire [7:0] _GEN_2479 = 8'h7 < length_0 ? _GEN_2319 : _GEN_2159; // @[executor.scala 308:60]
  wire [7:0] _GEN_2480 = 8'h7 < length_0 ? _GEN_2320 : _GEN_2160; // @[executor.scala 308:60]
  wire [7:0] _GEN_2481 = 8'h7 < length_0 ? _GEN_2321 : _GEN_2161; // @[executor.scala 308:60]
  wire [7:0] _GEN_2482 = 8'h7 < length_0 ? _GEN_2322 : _GEN_2162; // @[executor.scala 308:60]
  wire [7:0] _GEN_2483 = 8'h7 < length_0 ? _GEN_2323 : _GEN_2163; // @[executor.scala 308:60]
  wire [7:0] _GEN_2484 = 8'h7 < length_0 ? _GEN_2324 : _GEN_2164; // @[executor.scala 308:60]
  wire [7:0] _GEN_2485 = 8'h7 < length_0 ? _GEN_2325 : _GEN_2165; // @[executor.scala 308:60]
  wire [7:0] _GEN_2486 = 8'h7 < length_0 ? _GEN_2326 : _GEN_2166; // @[executor.scala 308:60]
  wire [7:0] _GEN_2487 = 8'h7 < length_0 ? _GEN_2327 : _GEN_2167; // @[executor.scala 308:60]
  wire [7:0] _GEN_2488 = 8'h7 < length_0 ? _GEN_2328 : _GEN_2168; // @[executor.scala 308:60]
  wire [7:0] _GEN_2489 = 8'h7 < length_0 ? _GEN_2329 : _GEN_2169; // @[executor.scala 308:60]
  wire [7:0] _GEN_2490 = 8'h7 < length_0 ? _GEN_2330 : _GEN_2170; // @[executor.scala 308:60]
  wire [7:0] _GEN_2491 = 8'h7 < length_0 ? _GEN_2331 : _GEN_2171; // @[executor.scala 308:60]
  wire [7:0] _GEN_2492 = 8'h7 < length_0 ? _GEN_2332 : _GEN_2172; // @[executor.scala 308:60]
  wire [7:0] _GEN_2493 = 8'h7 < length_0 ? _GEN_2333 : _GEN_2173; // @[executor.scala 308:60]
  wire [7:0] _GEN_2494 = 8'h7 < length_0 ? _GEN_2334 : _GEN_2174; // @[executor.scala 308:60]
  wire [7:0] _GEN_2495 = 8'h7 < length_0 ? _GEN_2335 : _GEN_2175; // @[executor.scala 308:60]
  wire [7:0] _GEN_2496 = 8'h7 < length_0 ? _GEN_2336 : _GEN_2176; // @[executor.scala 308:60]
  wire [7:0] _GEN_2497 = 8'h7 < length_0 ? _GEN_2337 : _GEN_2177; // @[executor.scala 308:60]
  wire [7:0] _GEN_2498 = 8'h7 < length_0 ? _GEN_2338 : _GEN_2178; // @[executor.scala 308:60]
  wire [7:0] _GEN_2499 = 8'h7 < length_0 ? _GEN_2339 : _GEN_2179; // @[executor.scala 308:60]
  wire [7:0] _GEN_2500 = 8'h7 < length_0 ? _GEN_2340 : _GEN_2180; // @[executor.scala 308:60]
  wire [7:0] _GEN_2501 = 8'h7 < length_0 ? _GEN_2341 : _GEN_2181; // @[executor.scala 308:60]
  wire [7:0] _GEN_2502 = 8'h7 < length_0 ? _GEN_2342 : _GEN_2182; // @[executor.scala 308:60]
  wire [7:0] _GEN_2503 = 8'h7 < length_0 ? _GEN_2343 : _GEN_2183; // @[executor.scala 308:60]
  wire [7:0] _GEN_2504 = 8'h7 < length_0 ? _GEN_2344 : _GEN_2184; // @[executor.scala 308:60]
  wire [7:0] _GEN_2505 = 8'h7 < length_0 ? _GEN_2345 : _GEN_2185; // @[executor.scala 308:60]
  wire [7:0] _GEN_2506 = 8'h7 < length_0 ? _GEN_2346 : _GEN_2186; // @[executor.scala 308:60]
  wire [7:0] _GEN_2507 = 8'h7 < length_0 ? _GEN_2347 : _GEN_2187; // @[executor.scala 308:60]
  wire [7:0] _GEN_2508 = 8'h7 < length_0 ? _GEN_2348 : _GEN_2188; // @[executor.scala 308:60]
  wire [7:0] _GEN_2509 = 8'h7 < length_0 ? _GEN_2349 : _GEN_2189; // @[executor.scala 308:60]
  wire [7:0] _GEN_2510 = 8'h7 < length_0 ? _GEN_2350 : _GEN_2190; // @[executor.scala 308:60]
  wire [7:0] _GEN_2511 = 8'h7 < length_0 ? _GEN_2351 : _GEN_2191; // @[executor.scala 308:60]
  wire [7:0] _GEN_2512 = 8'h7 < length_0 ? _GEN_2352 : _GEN_2192; // @[executor.scala 308:60]
  wire [7:0] _GEN_2513 = 8'h7 < length_0 ? _GEN_2353 : _GEN_2193; // @[executor.scala 308:60]
  wire [7:0] _GEN_2514 = 8'h7 < length_0 ? _GEN_2354 : _GEN_2194; // @[executor.scala 308:60]
  wire [7:0] _GEN_2515 = 8'h7 < length_0 ? _GEN_2355 : _GEN_2195; // @[executor.scala 308:60]
  wire [7:0] _GEN_2516 = 8'h7 < length_0 ? _GEN_2356 : _GEN_2196; // @[executor.scala 308:60]
  wire [7:0] _GEN_2517 = 8'h7 < length_0 ? _GEN_2357 : _GEN_2197; // @[executor.scala 308:60]
  wire [7:0] _GEN_2518 = 8'h7 < length_0 ? _GEN_2358 : _GEN_2198; // @[executor.scala 308:60]
  wire [7:0] _GEN_2519 = 8'h7 < length_0 ? _GEN_2359 : _GEN_2199; // @[executor.scala 308:60]
  wire [7:0] _GEN_2520 = 8'h7 < length_0 ? _GEN_2360 : _GEN_2200; // @[executor.scala 308:60]
  wire [7:0] _GEN_2521 = 8'h7 < length_0 ? _GEN_2361 : _GEN_2201; // @[executor.scala 308:60]
  wire [7:0] _GEN_2522 = 8'h7 < length_0 ? _GEN_2362 : _GEN_2202; // @[executor.scala 308:60]
  wire [7:0] _GEN_2523 = 8'h7 < length_0 ? _GEN_2363 : _GEN_2203; // @[executor.scala 308:60]
  wire [7:0] _GEN_2524 = 8'h7 < length_0 ? _GEN_2364 : _GEN_2204; // @[executor.scala 308:60]
  wire [7:0] _GEN_2525 = 8'h7 < length_0 ? _GEN_2365 : _GEN_2205; // @[executor.scala 308:60]
  wire [7:0] _GEN_2526 = 8'h7 < length_0 ? _GEN_2366 : _GEN_2206; // @[executor.scala 308:60]
  wire [7:0] _GEN_2527 = 8'h7 < length_0 ? _GEN_2367 : _GEN_2207; // @[executor.scala 308:60]
  wire [7:0] _GEN_2528 = 8'h7 < length_0 ? _GEN_2368 : _GEN_2208; // @[executor.scala 308:60]
  wire [7:0] _GEN_2529 = 8'h7 < length_0 ? _GEN_2369 : _GEN_2209; // @[executor.scala 308:60]
  wire [7:0] _GEN_2530 = 8'h7 < length_0 ? _GEN_2370 : _GEN_2210; // @[executor.scala 308:60]
  wire [7:0] _GEN_2531 = 8'h7 < length_0 ? _GEN_2371 : _GEN_2211; // @[executor.scala 308:60]
  wire [7:0] _GEN_2532 = 8'h7 < length_0 ? _GEN_2372 : _GEN_2212; // @[executor.scala 308:60]
  wire [7:0] _GEN_2533 = 8'h7 < length_0 ? _GEN_2373 : _GEN_2213; // @[executor.scala 308:60]
  wire [7:0] _GEN_2534 = 8'h7 < length_0 ? _GEN_2374 : _GEN_2214; // @[executor.scala 308:60]
  wire [7:0] _GEN_2535 = 8'h7 < length_0 ? _GEN_2375 : _GEN_2215; // @[executor.scala 308:60]
  wire [7:0] _GEN_2536 = 8'h7 < length_0 ? _GEN_2376 : _GEN_2216; // @[executor.scala 308:60]
  wire [7:0] _GEN_2537 = 8'h7 < length_0 ? _GEN_2377 : _GEN_2217; // @[executor.scala 308:60]
  wire [7:0] _GEN_2538 = 8'h7 < length_0 ? _GEN_2378 : _GEN_2218; // @[executor.scala 308:60]
  wire [7:0] _GEN_2539 = 8'h7 < length_0 ? _GEN_2379 : _GEN_2219; // @[executor.scala 308:60]
  wire [7:0] _GEN_2540 = 8'h7 < length_0 ? _GEN_2380 : _GEN_2220; // @[executor.scala 308:60]
  wire [7:0] _GEN_2541 = 8'h7 < length_0 ? _GEN_2381 : _GEN_2221; // @[executor.scala 308:60]
  wire [7:0] _GEN_2542 = 8'h7 < length_0 ? _GEN_2382 : _GEN_2222; // @[executor.scala 308:60]
  wire [7:0] _GEN_2543 = 8'h7 < length_0 ? _GEN_2383 : _GEN_2223; // @[executor.scala 308:60]
  wire [7:0] _GEN_2544 = 8'h7 < length_0 ? _GEN_2384 : _GEN_2224; // @[executor.scala 308:60]
  wire [7:0] _GEN_2545 = 8'h7 < length_0 ? _GEN_2385 : _GEN_2225; // @[executor.scala 308:60]
  wire [7:0] _GEN_2546 = 8'h7 < length_0 ? _GEN_2386 : _GEN_2226; // @[executor.scala 308:60]
  wire [7:0] _GEN_2547 = 8'h7 < length_0 ? _GEN_2387 : _GEN_2227; // @[executor.scala 308:60]
  wire [7:0] _GEN_2548 = 8'h7 < length_0 ? _GEN_2388 : _GEN_2228; // @[executor.scala 308:60]
  wire [7:0] _GEN_2549 = 8'h7 < length_0 ? _GEN_2389 : _GEN_2229; // @[executor.scala 308:60]
  wire [7:0] _GEN_2550 = 8'h7 < length_0 ? _GEN_2390 : _GEN_2230; // @[executor.scala 308:60]
  wire [7:0] _GEN_2551 = 8'h7 < length_0 ? _GEN_2391 : _GEN_2231; // @[executor.scala 308:60]
  wire [7:0] _GEN_2552 = 8'h7 < length_0 ? _GEN_2392 : _GEN_2232; // @[executor.scala 308:60]
  wire [7:0] _GEN_2553 = 8'h7 < length_0 ? _GEN_2393 : _GEN_2233; // @[executor.scala 308:60]
  wire [7:0] _GEN_2554 = 8'h7 < length_0 ? _GEN_2394 : _GEN_2234; // @[executor.scala 308:60]
  wire [7:0] _GEN_2555 = 8'h7 < length_0 ? _GEN_2395 : _GEN_2235; // @[executor.scala 308:60]
  wire [7:0] _GEN_2556 = 8'h7 < length_0 ? _GEN_2396 : _GEN_2236; // @[executor.scala 308:60]
  wire [7:0] _GEN_2557 = 8'h7 < length_0 ? _GEN_2397 : _GEN_2237; // @[executor.scala 308:60]
  wire [7:0] _GEN_2558 = 8'h7 < length_0 ? _GEN_2398 : _GEN_2238; // @[executor.scala 308:60]
  wire [7:0] _GEN_2559 = 8'h7 < length_0 ? _GEN_2399 : _GEN_2239; // @[executor.scala 308:60]
  wire [3:0] _GEN_2560 = length_0 == 8'h0 ? field_0[13:10] : phv_next_processor_id; // @[executor.scala 300:71 executor.scala 301:55 executor.scala 286:25]
  wire  _GEN_2561 = length_0 == 8'h0 ? field_0[0] : phv_next_config_id; // @[executor.scala 300:71 executor.scala 302:55 executor.scala 286:25]
  wire [7:0] _GEN_2562 = length_0 == 8'h0 ? phv_data_0 : _GEN_2400; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2563 = length_0 == 8'h0 ? phv_data_1 : _GEN_2401; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2564 = length_0 == 8'h0 ? phv_data_2 : _GEN_2402; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2565 = length_0 == 8'h0 ? phv_data_3 : _GEN_2403; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2566 = length_0 == 8'h0 ? phv_data_4 : _GEN_2404; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2567 = length_0 == 8'h0 ? phv_data_5 : _GEN_2405; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2568 = length_0 == 8'h0 ? phv_data_6 : _GEN_2406; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2569 = length_0 == 8'h0 ? phv_data_7 : _GEN_2407; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2570 = length_0 == 8'h0 ? phv_data_8 : _GEN_2408; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2571 = length_0 == 8'h0 ? phv_data_9 : _GEN_2409; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2572 = length_0 == 8'h0 ? phv_data_10 : _GEN_2410; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2573 = length_0 == 8'h0 ? phv_data_11 : _GEN_2411; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2574 = length_0 == 8'h0 ? phv_data_12 : _GEN_2412; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2575 = length_0 == 8'h0 ? phv_data_13 : _GEN_2413; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2576 = length_0 == 8'h0 ? phv_data_14 : _GEN_2414; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2577 = length_0 == 8'h0 ? phv_data_15 : _GEN_2415; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2578 = length_0 == 8'h0 ? phv_data_16 : _GEN_2416; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2579 = length_0 == 8'h0 ? phv_data_17 : _GEN_2417; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2580 = length_0 == 8'h0 ? phv_data_18 : _GEN_2418; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2581 = length_0 == 8'h0 ? phv_data_19 : _GEN_2419; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2582 = length_0 == 8'h0 ? phv_data_20 : _GEN_2420; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2583 = length_0 == 8'h0 ? phv_data_21 : _GEN_2421; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2584 = length_0 == 8'h0 ? phv_data_22 : _GEN_2422; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2585 = length_0 == 8'h0 ? phv_data_23 : _GEN_2423; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2586 = length_0 == 8'h0 ? phv_data_24 : _GEN_2424; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2587 = length_0 == 8'h0 ? phv_data_25 : _GEN_2425; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2588 = length_0 == 8'h0 ? phv_data_26 : _GEN_2426; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2589 = length_0 == 8'h0 ? phv_data_27 : _GEN_2427; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2590 = length_0 == 8'h0 ? phv_data_28 : _GEN_2428; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2591 = length_0 == 8'h0 ? phv_data_29 : _GEN_2429; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2592 = length_0 == 8'h0 ? phv_data_30 : _GEN_2430; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2593 = length_0 == 8'h0 ? phv_data_31 : _GEN_2431; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2594 = length_0 == 8'h0 ? phv_data_32 : _GEN_2432; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2595 = length_0 == 8'h0 ? phv_data_33 : _GEN_2433; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2596 = length_0 == 8'h0 ? phv_data_34 : _GEN_2434; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2597 = length_0 == 8'h0 ? phv_data_35 : _GEN_2435; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2598 = length_0 == 8'h0 ? phv_data_36 : _GEN_2436; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2599 = length_0 == 8'h0 ? phv_data_37 : _GEN_2437; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2600 = length_0 == 8'h0 ? phv_data_38 : _GEN_2438; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2601 = length_0 == 8'h0 ? phv_data_39 : _GEN_2439; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2602 = length_0 == 8'h0 ? phv_data_40 : _GEN_2440; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2603 = length_0 == 8'h0 ? phv_data_41 : _GEN_2441; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2604 = length_0 == 8'h0 ? phv_data_42 : _GEN_2442; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2605 = length_0 == 8'h0 ? phv_data_43 : _GEN_2443; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2606 = length_0 == 8'h0 ? phv_data_44 : _GEN_2444; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2607 = length_0 == 8'h0 ? phv_data_45 : _GEN_2445; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2608 = length_0 == 8'h0 ? phv_data_46 : _GEN_2446; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2609 = length_0 == 8'h0 ? phv_data_47 : _GEN_2447; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2610 = length_0 == 8'h0 ? phv_data_48 : _GEN_2448; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2611 = length_0 == 8'h0 ? phv_data_49 : _GEN_2449; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2612 = length_0 == 8'h0 ? phv_data_50 : _GEN_2450; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2613 = length_0 == 8'h0 ? phv_data_51 : _GEN_2451; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2614 = length_0 == 8'h0 ? phv_data_52 : _GEN_2452; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2615 = length_0 == 8'h0 ? phv_data_53 : _GEN_2453; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2616 = length_0 == 8'h0 ? phv_data_54 : _GEN_2454; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2617 = length_0 == 8'h0 ? phv_data_55 : _GEN_2455; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2618 = length_0 == 8'h0 ? phv_data_56 : _GEN_2456; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2619 = length_0 == 8'h0 ? phv_data_57 : _GEN_2457; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2620 = length_0 == 8'h0 ? phv_data_58 : _GEN_2458; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2621 = length_0 == 8'h0 ? phv_data_59 : _GEN_2459; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2622 = length_0 == 8'h0 ? phv_data_60 : _GEN_2460; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2623 = length_0 == 8'h0 ? phv_data_61 : _GEN_2461; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2624 = length_0 == 8'h0 ? phv_data_62 : _GEN_2462; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2625 = length_0 == 8'h0 ? phv_data_63 : _GEN_2463; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2626 = length_0 == 8'h0 ? phv_data_64 : _GEN_2464; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2627 = length_0 == 8'h0 ? phv_data_65 : _GEN_2465; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2628 = length_0 == 8'h0 ? phv_data_66 : _GEN_2466; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2629 = length_0 == 8'h0 ? phv_data_67 : _GEN_2467; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2630 = length_0 == 8'h0 ? phv_data_68 : _GEN_2468; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2631 = length_0 == 8'h0 ? phv_data_69 : _GEN_2469; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2632 = length_0 == 8'h0 ? phv_data_70 : _GEN_2470; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2633 = length_0 == 8'h0 ? phv_data_71 : _GEN_2471; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2634 = length_0 == 8'h0 ? phv_data_72 : _GEN_2472; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2635 = length_0 == 8'h0 ? phv_data_73 : _GEN_2473; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2636 = length_0 == 8'h0 ? phv_data_74 : _GEN_2474; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2637 = length_0 == 8'h0 ? phv_data_75 : _GEN_2475; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2638 = length_0 == 8'h0 ? phv_data_76 : _GEN_2476; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2639 = length_0 == 8'h0 ? phv_data_77 : _GEN_2477; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2640 = length_0 == 8'h0 ? phv_data_78 : _GEN_2478; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2641 = length_0 == 8'h0 ? phv_data_79 : _GEN_2479; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2642 = length_0 == 8'h0 ? phv_data_80 : _GEN_2480; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2643 = length_0 == 8'h0 ? phv_data_81 : _GEN_2481; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2644 = length_0 == 8'h0 ? phv_data_82 : _GEN_2482; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2645 = length_0 == 8'h0 ? phv_data_83 : _GEN_2483; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2646 = length_0 == 8'h0 ? phv_data_84 : _GEN_2484; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2647 = length_0 == 8'h0 ? phv_data_85 : _GEN_2485; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2648 = length_0 == 8'h0 ? phv_data_86 : _GEN_2486; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2649 = length_0 == 8'h0 ? phv_data_87 : _GEN_2487; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2650 = length_0 == 8'h0 ? phv_data_88 : _GEN_2488; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2651 = length_0 == 8'h0 ? phv_data_89 : _GEN_2489; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2652 = length_0 == 8'h0 ? phv_data_90 : _GEN_2490; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2653 = length_0 == 8'h0 ? phv_data_91 : _GEN_2491; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2654 = length_0 == 8'h0 ? phv_data_92 : _GEN_2492; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2655 = length_0 == 8'h0 ? phv_data_93 : _GEN_2493; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2656 = length_0 == 8'h0 ? phv_data_94 : _GEN_2494; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2657 = length_0 == 8'h0 ? phv_data_95 : _GEN_2495; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2658 = length_0 == 8'h0 ? phv_data_96 : _GEN_2496; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2659 = length_0 == 8'h0 ? phv_data_97 : _GEN_2497; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2660 = length_0 == 8'h0 ? phv_data_98 : _GEN_2498; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2661 = length_0 == 8'h0 ? phv_data_99 : _GEN_2499; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2662 = length_0 == 8'h0 ? phv_data_100 : _GEN_2500; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2663 = length_0 == 8'h0 ? phv_data_101 : _GEN_2501; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2664 = length_0 == 8'h0 ? phv_data_102 : _GEN_2502; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2665 = length_0 == 8'h0 ? phv_data_103 : _GEN_2503; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2666 = length_0 == 8'h0 ? phv_data_104 : _GEN_2504; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2667 = length_0 == 8'h0 ? phv_data_105 : _GEN_2505; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2668 = length_0 == 8'h0 ? phv_data_106 : _GEN_2506; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2669 = length_0 == 8'h0 ? phv_data_107 : _GEN_2507; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2670 = length_0 == 8'h0 ? phv_data_108 : _GEN_2508; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2671 = length_0 == 8'h0 ? phv_data_109 : _GEN_2509; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2672 = length_0 == 8'h0 ? phv_data_110 : _GEN_2510; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2673 = length_0 == 8'h0 ? phv_data_111 : _GEN_2511; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2674 = length_0 == 8'h0 ? phv_data_112 : _GEN_2512; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2675 = length_0 == 8'h0 ? phv_data_113 : _GEN_2513; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2676 = length_0 == 8'h0 ? phv_data_114 : _GEN_2514; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2677 = length_0 == 8'h0 ? phv_data_115 : _GEN_2515; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2678 = length_0 == 8'h0 ? phv_data_116 : _GEN_2516; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2679 = length_0 == 8'h0 ? phv_data_117 : _GEN_2517; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2680 = length_0 == 8'h0 ? phv_data_118 : _GEN_2518; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2681 = length_0 == 8'h0 ? phv_data_119 : _GEN_2519; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2682 = length_0 == 8'h0 ? phv_data_120 : _GEN_2520; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2683 = length_0 == 8'h0 ? phv_data_121 : _GEN_2521; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2684 = length_0 == 8'h0 ? phv_data_122 : _GEN_2522; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2685 = length_0 == 8'h0 ? phv_data_123 : _GEN_2523; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2686 = length_0 == 8'h0 ? phv_data_124 : _GEN_2524; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2687 = length_0 == 8'h0 ? phv_data_125 : _GEN_2525; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2688 = length_0 == 8'h0 ? phv_data_126 : _GEN_2526; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2689 = length_0 == 8'h0 ? phv_data_127 : _GEN_2527; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2690 = length_0 == 8'h0 ? phv_data_128 : _GEN_2528; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2691 = length_0 == 8'h0 ? phv_data_129 : _GEN_2529; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2692 = length_0 == 8'h0 ? phv_data_130 : _GEN_2530; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2693 = length_0 == 8'h0 ? phv_data_131 : _GEN_2531; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2694 = length_0 == 8'h0 ? phv_data_132 : _GEN_2532; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2695 = length_0 == 8'h0 ? phv_data_133 : _GEN_2533; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2696 = length_0 == 8'h0 ? phv_data_134 : _GEN_2534; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2697 = length_0 == 8'h0 ? phv_data_135 : _GEN_2535; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2698 = length_0 == 8'h0 ? phv_data_136 : _GEN_2536; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2699 = length_0 == 8'h0 ? phv_data_137 : _GEN_2537; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2700 = length_0 == 8'h0 ? phv_data_138 : _GEN_2538; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2701 = length_0 == 8'h0 ? phv_data_139 : _GEN_2539; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2702 = length_0 == 8'h0 ? phv_data_140 : _GEN_2540; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2703 = length_0 == 8'h0 ? phv_data_141 : _GEN_2541; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2704 = length_0 == 8'h0 ? phv_data_142 : _GEN_2542; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2705 = length_0 == 8'h0 ? phv_data_143 : _GEN_2543; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2706 = length_0 == 8'h0 ? phv_data_144 : _GEN_2544; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2707 = length_0 == 8'h0 ? phv_data_145 : _GEN_2545; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2708 = length_0 == 8'h0 ? phv_data_146 : _GEN_2546; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2709 = length_0 == 8'h0 ? phv_data_147 : _GEN_2547; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2710 = length_0 == 8'h0 ? phv_data_148 : _GEN_2548; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2711 = length_0 == 8'h0 ? phv_data_149 : _GEN_2549; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2712 = length_0 == 8'h0 ? phv_data_150 : _GEN_2550; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2713 = length_0 == 8'h0 ? phv_data_151 : _GEN_2551; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2714 = length_0 == 8'h0 ? phv_data_152 : _GEN_2552; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2715 = length_0 == 8'h0 ? phv_data_153 : _GEN_2553; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2716 = length_0 == 8'h0 ? phv_data_154 : _GEN_2554; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2717 = length_0 == 8'h0 ? phv_data_155 : _GEN_2555; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2718 = length_0 == 8'h0 ? phv_data_156 : _GEN_2556; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2719 = length_0 == 8'h0 ? phv_data_157 : _GEN_2557; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2720 = length_0 == 8'h0 ? phv_data_158 : _GEN_2558; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] _GEN_2721 = length_0 == 8'h0 ? phv_data_159 : _GEN_2559; // @[executor.scala 300:71 executor.scala 286:25]
  wire [7:0] field_byte_8 = field_1[63:56]; // @[executor.scala 305:57]
  wire [8:0] _total_offset_T_8 = {{1'd0}, offset_1}; // @[executor.scala 307:57]
  wire [7:0] total_offset_8 = _total_offset_T_8[7:0]; // @[executor.scala 307:57]
  wire [7:0] _GEN_2722 = 8'h0 == total_offset_8 ? field_byte_8 : _GEN_2562; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2723 = 8'h1 == total_offset_8 ? field_byte_8 : _GEN_2563; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2724 = 8'h2 == total_offset_8 ? field_byte_8 : _GEN_2564; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2725 = 8'h3 == total_offset_8 ? field_byte_8 : _GEN_2565; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2726 = 8'h4 == total_offset_8 ? field_byte_8 : _GEN_2566; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2727 = 8'h5 == total_offset_8 ? field_byte_8 : _GEN_2567; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2728 = 8'h6 == total_offset_8 ? field_byte_8 : _GEN_2568; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2729 = 8'h7 == total_offset_8 ? field_byte_8 : _GEN_2569; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2730 = 8'h8 == total_offset_8 ? field_byte_8 : _GEN_2570; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2731 = 8'h9 == total_offset_8 ? field_byte_8 : _GEN_2571; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2732 = 8'ha == total_offset_8 ? field_byte_8 : _GEN_2572; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2733 = 8'hb == total_offset_8 ? field_byte_8 : _GEN_2573; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2734 = 8'hc == total_offset_8 ? field_byte_8 : _GEN_2574; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2735 = 8'hd == total_offset_8 ? field_byte_8 : _GEN_2575; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2736 = 8'he == total_offset_8 ? field_byte_8 : _GEN_2576; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2737 = 8'hf == total_offset_8 ? field_byte_8 : _GEN_2577; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2738 = 8'h10 == total_offset_8 ? field_byte_8 : _GEN_2578; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2739 = 8'h11 == total_offset_8 ? field_byte_8 : _GEN_2579; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2740 = 8'h12 == total_offset_8 ? field_byte_8 : _GEN_2580; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2741 = 8'h13 == total_offset_8 ? field_byte_8 : _GEN_2581; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2742 = 8'h14 == total_offset_8 ? field_byte_8 : _GEN_2582; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2743 = 8'h15 == total_offset_8 ? field_byte_8 : _GEN_2583; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2744 = 8'h16 == total_offset_8 ? field_byte_8 : _GEN_2584; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2745 = 8'h17 == total_offset_8 ? field_byte_8 : _GEN_2585; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2746 = 8'h18 == total_offset_8 ? field_byte_8 : _GEN_2586; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2747 = 8'h19 == total_offset_8 ? field_byte_8 : _GEN_2587; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2748 = 8'h1a == total_offset_8 ? field_byte_8 : _GEN_2588; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2749 = 8'h1b == total_offset_8 ? field_byte_8 : _GEN_2589; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2750 = 8'h1c == total_offset_8 ? field_byte_8 : _GEN_2590; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2751 = 8'h1d == total_offset_8 ? field_byte_8 : _GEN_2591; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2752 = 8'h1e == total_offset_8 ? field_byte_8 : _GEN_2592; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2753 = 8'h1f == total_offset_8 ? field_byte_8 : _GEN_2593; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2754 = 8'h20 == total_offset_8 ? field_byte_8 : _GEN_2594; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2755 = 8'h21 == total_offset_8 ? field_byte_8 : _GEN_2595; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2756 = 8'h22 == total_offset_8 ? field_byte_8 : _GEN_2596; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2757 = 8'h23 == total_offset_8 ? field_byte_8 : _GEN_2597; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2758 = 8'h24 == total_offset_8 ? field_byte_8 : _GEN_2598; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2759 = 8'h25 == total_offset_8 ? field_byte_8 : _GEN_2599; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2760 = 8'h26 == total_offset_8 ? field_byte_8 : _GEN_2600; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2761 = 8'h27 == total_offset_8 ? field_byte_8 : _GEN_2601; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2762 = 8'h28 == total_offset_8 ? field_byte_8 : _GEN_2602; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2763 = 8'h29 == total_offset_8 ? field_byte_8 : _GEN_2603; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2764 = 8'h2a == total_offset_8 ? field_byte_8 : _GEN_2604; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2765 = 8'h2b == total_offset_8 ? field_byte_8 : _GEN_2605; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2766 = 8'h2c == total_offset_8 ? field_byte_8 : _GEN_2606; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2767 = 8'h2d == total_offset_8 ? field_byte_8 : _GEN_2607; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2768 = 8'h2e == total_offset_8 ? field_byte_8 : _GEN_2608; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2769 = 8'h2f == total_offset_8 ? field_byte_8 : _GEN_2609; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2770 = 8'h30 == total_offset_8 ? field_byte_8 : _GEN_2610; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2771 = 8'h31 == total_offset_8 ? field_byte_8 : _GEN_2611; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2772 = 8'h32 == total_offset_8 ? field_byte_8 : _GEN_2612; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2773 = 8'h33 == total_offset_8 ? field_byte_8 : _GEN_2613; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2774 = 8'h34 == total_offset_8 ? field_byte_8 : _GEN_2614; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2775 = 8'h35 == total_offset_8 ? field_byte_8 : _GEN_2615; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2776 = 8'h36 == total_offset_8 ? field_byte_8 : _GEN_2616; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2777 = 8'h37 == total_offset_8 ? field_byte_8 : _GEN_2617; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2778 = 8'h38 == total_offset_8 ? field_byte_8 : _GEN_2618; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2779 = 8'h39 == total_offset_8 ? field_byte_8 : _GEN_2619; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2780 = 8'h3a == total_offset_8 ? field_byte_8 : _GEN_2620; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2781 = 8'h3b == total_offset_8 ? field_byte_8 : _GEN_2621; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2782 = 8'h3c == total_offset_8 ? field_byte_8 : _GEN_2622; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2783 = 8'h3d == total_offset_8 ? field_byte_8 : _GEN_2623; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2784 = 8'h3e == total_offset_8 ? field_byte_8 : _GEN_2624; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2785 = 8'h3f == total_offset_8 ? field_byte_8 : _GEN_2625; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2786 = 8'h40 == total_offset_8 ? field_byte_8 : _GEN_2626; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2787 = 8'h41 == total_offset_8 ? field_byte_8 : _GEN_2627; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2788 = 8'h42 == total_offset_8 ? field_byte_8 : _GEN_2628; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2789 = 8'h43 == total_offset_8 ? field_byte_8 : _GEN_2629; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2790 = 8'h44 == total_offset_8 ? field_byte_8 : _GEN_2630; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2791 = 8'h45 == total_offset_8 ? field_byte_8 : _GEN_2631; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2792 = 8'h46 == total_offset_8 ? field_byte_8 : _GEN_2632; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2793 = 8'h47 == total_offset_8 ? field_byte_8 : _GEN_2633; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2794 = 8'h48 == total_offset_8 ? field_byte_8 : _GEN_2634; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2795 = 8'h49 == total_offset_8 ? field_byte_8 : _GEN_2635; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2796 = 8'h4a == total_offset_8 ? field_byte_8 : _GEN_2636; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2797 = 8'h4b == total_offset_8 ? field_byte_8 : _GEN_2637; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2798 = 8'h4c == total_offset_8 ? field_byte_8 : _GEN_2638; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2799 = 8'h4d == total_offset_8 ? field_byte_8 : _GEN_2639; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2800 = 8'h4e == total_offset_8 ? field_byte_8 : _GEN_2640; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2801 = 8'h4f == total_offset_8 ? field_byte_8 : _GEN_2641; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2802 = 8'h50 == total_offset_8 ? field_byte_8 : _GEN_2642; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2803 = 8'h51 == total_offset_8 ? field_byte_8 : _GEN_2643; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2804 = 8'h52 == total_offset_8 ? field_byte_8 : _GEN_2644; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2805 = 8'h53 == total_offset_8 ? field_byte_8 : _GEN_2645; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2806 = 8'h54 == total_offset_8 ? field_byte_8 : _GEN_2646; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2807 = 8'h55 == total_offset_8 ? field_byte_8 : _GEN_2647; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2808 = 8'h56 == total_offset_8 ? field_byte_8 : _GEN_2648; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2809 = 8'h57 == total_offset_8 ? field_byte_8 : _GEN_2649; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2810 = 8'h58 == total_offset_8 ? field_byte_8 : _GEN_2650; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2811 = 8'h59 == total_offset_8 ? field_byte_8 : _GEN_2651; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2812 = 8'h5a == total_offset_8 ? field_byte_8 : _GEN_2652; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2813 = 8'h5b == total_offset_8 ? field_byte_8 : _GEN_2653; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2814 = 8'h5c == total_offset_8 ? field_byte_8 : _GEN_2654; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2815 = 8'h5d == total_offset_8 ? field_byte_8 : _GEN_2655; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2816 = 8'h5e == total_offset_8 ? field_byte_8 : _GEN_2656; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2817 = 8'h5f == total_offset_8 ? field_byte_8 : _GEN_2657; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2818 = 8'h60 == total_offset_8 ? field_byte_8 : _GEN_2658; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2819 = 8'h61 == total_offset_8 ? field_byte_8 : _GEN_2659; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2820 = 8'h62 == total_offset_8 ? field_byte_8 : _GEN_2660; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2821 = 8'h63 == total_offset_8 ? field_byte_8 : _GEN_2661; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2822 = 8'h64 == total_offset_8 ? field_byte_8 : _GEN_2662; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2823 = 8'h65 == total_offset_8 ? field_byte_8 : _GEN_2663; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2824 = 8'h66 == total_offset_8 ? field_byte_8 : _GEN_2664; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2825 = 8'h67 == total_offset_8 ? field_byte_8 : _GEN_2665; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2826 = 8'h68 == total_offset_8 ? field_byte_8 : _GEN_2666; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2827 = 8'h69 == total_offset_8 ? field_byte_8 : _GEN_2667; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2828 = 8'h6a == total_offset_8 ? field_byte_8 : _GEN_2668; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2829 = 8'h6b == total_offset_8 ? field_byte_8 : _GEN_2669; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2830 = 8'h6c == total_offset_8 ? field_byte_8 : _GEN_2670; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2831 = 8'h6d == total_offset_8 ? field_byte_8 : _GEN_2671; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2832 = 8'h6e == total_offset_8 ? field_byte_8 : _GEN_2672; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2833 = 8'h6f == total_offset_8 ? field_byte_8 : _GEN_2673; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2834 = 8'h70 == total_offset_8 ? field_byte_8 : _GEN_2674; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2835 = 8'h71 == total_offset_8 ? field_byte_8 : _GEN_2675; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2836 = 8'h72 == total_offset_8 ? field_byte_8 : _GEN_2676; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2837 = 8'h73 == total_offset_8 ? field_byte_8 : _GEN_2677; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2838 = 8'h74 == total_offset_8 ? field_byte_8 : _GEN_2678; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2839 = 8'h75 == total_offset_8 ? field_byte_8 : _GEN_2679; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2840 = 8'h76 == total_offset_8 ? field_byte_8 : _GEN_2680; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2841 = 8'h77 == total_offset_8 ? field_byte_8 : _GEN_2681; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2842 = 8'h78 == total_offset_8 ? field_byte_8 : _GEN_2682; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2843 = 8'h79 == total_offset_8 ? field_byte_8 : _GEN_2683; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2844 = 8'h7a == total_offset_8 ? field_byte_8 : _GEN_2684; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2845 = 8'h7b == total_offset_8 ? field_byte_8 : _GEN_2685; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2846 = 8'h7c == total_offset_8 ? field_byte_8 : _GEN_2686; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2847 = 8'h7d == total_offset_8 ? field_byte_8 : _GEN_2687; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2848 = 8'h7e == total_offset_8 ? field_byte_8 : _GEN_2688; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2849 = 8'h7f == total_offset_8 ? field_byte_8 : _GEN_2689; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2850 = 8'h80 == total_offset_8 ? field_byte_8 : _GEN_2690; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2851 = 8'h81 == total_offset_8 ? field_byte_8 : _GEN_2691; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2852 = 8'h82 == total_offset_8 ? field_byte_8 : _GEN_2692; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2853 = 8'h83 == total_offset_8 ? field_byte_8 : _GEN_2693; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2854 = 8'h84 == total_offset_8 ? field_byte_8 : _GEN_2694; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2855 = 8'h85 == total_offset_8 ? field_byte_8 : _GEN_2695; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2856 = 8'h86 == total_offset_8 ? field_byte_8 : _GEN_2696; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2857 = 8'h87 == total_offset_8 ? field_byte_8 : _GEN_2697; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2858 = 8'h88 == total_offset_8 ? field_byte_8 : _GEN_2698; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2859 = 8'h89 == total_offset_8 ? field_byte_8 : _GEN_2699; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2860 = 8'h8a == total_offset_8 ? field_byte_8 : _GEN_2700; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2861 = 8'h8b == total_offset_8 ? field_byte_8 : _GEN_2701; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2862 = 8'h8c == total_offset_8 ? field_byte_8 : _GEN_2702; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2863 = 8'h8d == total_offset_8 ? field_byte_8 : _GEN_2703; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2864 = 8'h8e == total_offset_8 ? field_byte_8 : _GEN_2704; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2865 = 8'h8f == total_offset_8 ? field_byte_8 : _GEN_2705; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2866 = 8'h90 == total_offset_8 ? field_byte_8 : _GEN_2706; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2867 = 8'h91 == total_offset_8 ? field_byte_8 : _GEN_2707; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2868 = 8'h92 == total_offset_8 ? field_byte_8 : _GEN_2708; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2869 = 8'h93 == total_offset_8 ? field_byte_8 : _GEN_2709; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2870 = 8'h94 == total_offset_8 ? field_byte_8 : _GEN_2710; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2871 = 8'h95 == total_offset_8 ? field_byte_8 : _GEN_2711; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2872 = 8'h96 == total_offset_8 ? field_byte_8 : _GEN_2712; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2873 = 8'h97 == total_offset_8 ? field_byte_8 : _GEN_2713; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2874 = 8'h98 == total_offset_8 ? field_byte_8 : _GEN_2714; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2875 = 8'h99 == total_offset_8 ? field_byte_8 : _GEN_2715; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2876 = 8'h9a == total_offset_8 ? field_byte_8 : _GEN_2716; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2877 = 8'h9b == total_offset_8 ? field_byte_8 : _GEN_2717; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2878 = 8'h9c == total_offset_8 ? field_byte_8 : _GEN_2718; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2879 = 8'h9d == total_offset_8 ? field_byte_8 : _GEN_2719; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2880 = 8'h9e == total_offset_8 ? field_byte_8 : _GEN_2720; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2881 = 8'h9f == total_offset_8 ? field_byte_8 : _GEN_2721; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_2882 = 8'h0 < length_1 ? _GEN_2722 : _GEN_2562; // @[executor.scala 308:60]
  wire [7:0] _GEN_2883 = 8'h0 < length_1 ? _GEN_2723 : _GEN_2563; // @[executor.scala 308:60]
  wire [7:0] _GEN_2884 = 8'h0 < length_1 ? _GEN_2724 : _GEN_2564; // @[executor.scala 308:60]
  wire [7:0] _GEN_2885 = 8'h0 < length_1 ? _GEN_2725 : _GEN_2565; // @[executor.scala 308:60]
  wire [7:0] _GEN_2886 = 8'h0 < length_1 ? _GEN_2726 : _GEN_2566; // @[executor.scala 308:60]
  wire [7:0] _GEN_2887 = 8'h0 < length_1 ? _GEN_2727 : _GEN_2567; // @[executor.scala 308:60]
  wire [7:0] _GEN_2888 = 8'h0 < length_1 ? _GEN_2728 : _GEN_2568; // @[executor.scala 308:60]
  wire [7:0] _GEN_2889 = 8'h0 < length_1 ? _GEN_2729 : _GEN_2569; // @[executor.scala 308:60]
  wire [7:0] _GEN_2890 = 8'h0 < length_1 ? _GEN_2730 : _GEN_2570; // @[executor.scala 308:60]
  wire [7:0] _GEN_2891 = 8'h0 < length_1 ? _GEN_2731 : _GEN_2571; // @[executor.scala 308:60]
  wire [7:0] _GEN_2892 = 8'h0 < length_1 ? _GEN_2732 : _GEN_2572; // @[executor.scala 308:60]
  wire [7:0] _GEN_2893 = 8'h0 < length_1 ? _GEN_2733 : _GEN_2573; // @[executor.scala 308:60]
  wire [7:0] _GEN_2894 = 8'h0 < length_1 ? _GEN_2734 : _GEN_2574; // @[executor.scala 308:60]
  wire [7:0] _GEN_2895 = 8'h0 < length_1 ? _GEN_2735 : _GEN_2575; // @[executor.scala 308:60]
  wire [7:0] _GEN_2896 = 8'h0 < length_1 ? _GEN_2736 : _GEN_2576; // @[executor.scala 308:60]
  wire [7:0] _GEN_2897 = 8'h0 < length_1 ? _GEN_2737 : _GEN_2577; // @[executor.scala 308:60]
  wire [7:0] _GEN_2898 = 8'h0 < length_1 ? _GEN_2738 : _GEN_2578; // @[executor.scala 308:60]
  wire [7:0] _GEN_2899 = 8'h0 < length_1 ? _GEN_2739 : _GEN_2579; // @[executor.scala 308:60]
  wire [7:0] _GEN_2900 = 8'h0 < length_1 ? _GEN_2740 : _GEN_2580; // @[executor.scala 308:60]
  wire [7:0] _GEN_2901 = 8'h0 < length_1 ? _GEN_2741 : _GEN_2581; // @[executor.scala 308:60]
  wire [7:0] _GEN_2902 = 8'h0 < length_1 ? _GEN_2742 : _GEN_2582; // @[executor.scala 308:60]
  wire [7:0] _GEN_2903 = 8'h0 < length_1 ? _GEN_2743 : _GEN_2583; // @[executor.scala 308:60]
  wire [7:0] _GEN_2904 = 8'h0 < length_1 ? _GEN_2744 : _GEN_2584; // @[executor.scala 308:60]
  wire [7:0] _GEN_2905 = 8'h0 < length_1 ? _GEN_2745 : _GEN_2585; // @[executor.scala 308:60]
  wire [7:0] _GEN_2906 = 8'h0 < length_1 ? _GEN_2746 : _GEN_2586; // @[executor.scala 308:60]
  wire [7:0] _GEN_2907 = 8'h0 < length_1 ? _GEN_2747 : _GEN_2587; // @[executor.scala 308:60]
  wire [7:0] _GEN_2908 = 8'h0 < length_1 ? _GEN_2748 : _GEN_2588; // @[executor.scala 308:60]
  wire [7:0] _GEN_2909 = 8'h0 < length_1 ? _GEN_2749 : _GEN_2589; // @[executor.scala 308:60]
  wire [7:0] _GEN_2910 = 8'h0 < length_1 ? _GEN_2750 : _GEN_2590; // @[executor.scala 308:60]
  wire [7:0] _GEN_2911 = 8'h0 < length_1 ? _GEN_2751 : _GEN_2591; // @[executor.scala 308:60]
  wire [7:0] _GEN_2912 = 8'h0 < length_1 ? _GEN_2752 : _GEN_2592; // @[executor.scala 308:60]
  wire [7:0] _GEN_2913 = 8'h0 < length_1 ? _GEN_2753 : _GEN_2593; // @[executor.scala 308:60]
  wire [7:0] _GEN_2914 = 8'h0 < length_1 ? _GEN_2754 : _GEN_2594; // @[executor.scala 308:60]
  wire [7:0] _GEN_2915 = 8'h0 < length_1 ? _GEN_2755 : _GEN_2595; // @[executor.scala 308:60]
  wire [7:0] _GEN_2916 = 8'h0 < length_1 ? _GEN_2756 : _GEN_2596; // @[executor.scala 308:60]
  wire [7:0] _GEN_2917 = 8'h0 < length_1 ? _GEN_2757 : _GEN_2597; // @[executor.scala 308:60]
  wire [7:0] _GEN_2918 = 8'h0 < length_1 ? _GEN_2758 : _GEN_2598; // @[executor.scala 308:60]
  wire [7:0] _GEN_2919 = 8'h0 < length_1 ? _GEN_2759 : _GEN_2599; // @[executor.scala 308:60]
  wire [7:0] _GEN_2920 = 8'h0 < length_1 ? _GEN_2760 : _GEN_2600; // @[executor.scala 308:60]
  wire [7:0] _GEN_2921 = 8'h0 < length_1 ? _GEN_2761 : _GEN_2601; // @[executor.scala 308:60]
  wire [7:0] _GEN_2922 = 8'h0 < length_1 ? _GEN_2762 : _GEN_2602; // @[executor.scala 308:60]
  wire [7:0] _GEN_2923 = 8'h0 < length_1 ? _GEN_2763 : _GEN_2603; // @[executor.scala 308:60]
  wire [7:0] _GEN_2924 = 8'h0 < length_1 ? _GEN_2764 : _GEN_2604; // @[executor.scala 308:60]
  wire [7:0] _GEN_2925 = 8'h0 < length_1 ? _GEN_2765 : _GEN_2605; // @[executor.scala 308:60]
  wire [7:0] _GEN_2926 = 8'h0 < length_1 ? _GEN_2766 : _GEN_2606; // @[executor.scala 308:60]
  wire [7:0] _GEN_2927 = 8'h0 < length_1 ? _GEN_2767 : _GEN_2607; // @[executor.scala 308:60]
  wire [7:0] _GEN_2928 = 8'h0 < length_1 ? _GEN_2768 : _GEN_2608; // @[executor.scala 308:60]
  wire [7:0] _GEN_2929 = 8'h0 < length_1 ? _GEN_2769 : _GEN_2609; // @[executor.scala 308:60]
  wire [7:0] _GEN_2930 = 8'h0 < length_1 ? _GEN_2770 : _GEN_2610; // @[executor.scala 308:60]
  wire [7:0] _GEN_2931 = 8'h0 < length_1 ? _GEN_2771 : _GEN_2611; // @[executor.scala 308:60]
  wire [7:0] _GEN_2932 = 8'h0 < length_1 ? _GEN_2772 : _GEN_2612; // @[executor.scala 308:60]
  wire [7:0] _GEN_2933 = 8'h0 < length_1 ? _GEN_2773 : _GEN_2613; // @[executor.scala 308:60]
  wire [7:0] _GEN_2934 = 8'h0 < length_1 ? _GEN_2774 : _GEN_2614; // @[executor.scala 308:60]
  wire [7:0] _GEN_2935 = 8'h0 < length_1 ? _GEN_2775 : _GEN_2615; // @[executor.scala 308:60]
  wire [7:0] _GEN_2936 = 8'h0 < length_1 ? _GEN_2776 : _GEN_2616; // @[executor.scala 308:60]
  wire [7:0] _GEN_2937 = 8'h0 < length_1 ? _GEN_2777 : _GEN_2617; // @[executor.scala 308:60]
  wire [7:0] _GEN_2938 = 8'h0 < length_1 ? _GEN_2778 : _GEN_2618; // @[executor.scala 308:60]
  wire [7:0] _GEN_2939 = 8'h0 < length_1 ? _GEN_2779 : _GEN_2619; // @[executor.scala 308:60]
  wire [7:0] _GEN_2940 = 8'h0 < length_1 ? _GEN_2780 : _GEN_2620; // @[executor.scala 308:60]
  wire [7:0] _GEN_2941 = 8'h0 < length_1 ? _GEN_2781 : _GEN_2621; // @[executor.scala 308:60]
  wire [7:0] _GEN_2942 = 8'h0 < length_1 ? _GEN_2782 : _GEN_2622; // @[executor.scala 308:60]
  wire [7:0] _GEN_2943 = 8'h0 < length_1 ? _GEN_2783 : _GEN_2623; // @[executor.scala 308:60]
  wire [7:0] _GEN_2944 = 8'h0 < length_1 ? _GEN_2784 : _GEN_2624; // @[executor.scala 308:60]
  wire [7:0] _GEN_2945 = 8'h0 < length_1 ? _GEN_2785 : _GEN_2625; // @[executor.scala 308:60]
  wire [7:0] _GEN_2946 = 8'h0 < length_1 ? _GEN_2786 : _GEN_2626; // @[executor.scala 308:60]
  wire [7:0] _GEN_2947 = 8'h0 < length_1 ? _GEN_2787 : _GEN_2627; // @[executor.scala 308:60]
  wire [7:0] _GEN_2948 = 8'h0 < length_1 ? _GEN_2788 : _GEN_2628; // @[executor.scala 308:60]
  wire [7:0] _GEN_2949 = 8'h0 < length_1 ? _GEN_2789 : _GEN_2629; // @[executor.scala 308:60]
  wire [7:0] _GEN_2950 = 8'h0 < length_1 ? _GEN_2790 : _GEN_2630; // @[executor.scala 308:60]
  wire [7:0] _GEN_2951 = 8'h0 < length_1 ? _GEN_2791 : _GEN_2631; // @[executor.scala 308:60]
  wire [7:0] _GEN_2952 = 8'h0 < length_1 ? _GEN_2792 : _GEN_2632; // @[executor.scala 308:60]
  wire [7:0] _GEN_2953 = 8'h0 < length_1 ? _GEN_2793 : _GEN_2633; // @[executor.scala 308:60]
  wire [7:0] _GEN_2954 = 8'h0 < length_1 ? _GEN_2794 : _GEN_2634; // @[executor.scala 308:60]
  wire [7:0] _GEN_2955 = 8'h0 < length_1 ? _GEN_2795 : _GEN_2635; // @[executor.scala 308:60]
  wire [7:0] _GEN_2956 = 8'h0 < length_1 ? _GEN_2796 : _GEN_2636; // @[executor.scala 308:60]
  wire [7:0] _GEN_2957 = 8'h0 < length_1 ? _GEN_2797 : _GEN_2637; // @[executor.scala 308:60]
  wire [7:0] _GEN_2958 = 8'h0 < length_1 ? _GEN_2798 : _GEN_2638; // @[executor.scala 308:60]
  wire [7:0] _GEN_2959 = 8'h0 < length_1 ? _GEN_2799 : _GEN_2639; // @[executor.scala 308:60]
  wire [7:0] _GEN_2960 = 8'h0 < length_1 ? _GEN_2800 : _GEN_2640; // @[executor.scala 308:60]
  wire [7:0] _GEN_2961 = 8'h0 < length_1 ? _GEN_2801 : _GEN_2641; // @[executor.scala 308:60]
  wire [7:0] _GEN_2962 = 8'h0 < length_1 ? _GEN_2802 : _GEN_2642; // @[executor.scala 308:60]
  wire [7:0] _GEN_2963 = 8'h0 < length_1 ? _GEN_2803 : _GEN_2643; // @[executor.scala 308:60]
  wire [7:0] _GEN_2964 = 8'h0 < length_1 ? _GEN_2804 : _GEN_2644; // @[executor.scala 308:60]
  wire [7:0] _GEN_2965 = 8'h0 < length_1 ? _GEN_2805 : _GEN_2645; // @[executor.scala 308:60]
  wire [7:0] _GEN_2966 = 8'h0 < length_1 ? _GEN_2806 : _GEN_2646; // @[executor.scala 308:60]
  wire [7:0] _GEN_2967 = 8'h0 < length_1 ? _GEN_2807 : _GEN_2647; // @[executor.scala 308:60]
  wire [7:0] _GEN_2968 = 8'h0 < length_1 ? _GEN_2808 : _GEN_2648; // @[executor.scala 308:60]
  wire [7:0] _GEN_2969 = 8'h0 < length_1 ? _GEN_2809 : _GEN_2649; // @[executor.scala 308:60]
  wire [7:0] _GEN_2970 = 8'h0 < length_1 ? _GEN_2810 : _GEN_2650; // @[executor.scala 308:60]
  wire [7:0] _GEN_2971 = 8'h0 < length_1 ? _GEN_2811 : _GEN_2651; // @[executor.scala 308:60]
  wire [7:0] _GEN_2972 = 8'h0 < length_1 ? _GEN_2812 : _GEN_2652; // @[executor.scala 308:60]
  wire [7:0] _GEN_2973 = 8'h0 < length_1 ? _GEN_2813 : _GEN_2653; // @[executor.scala 308:60]
  wire [7:0] _GEN_2974 = 8'h0 < length_1 ? _GEN_2814 : _GEN_2654; // @[executor.scala 308:60]
  wire [7:0] _GEN_2975 = 8'h0 < length_1 ? _GEN_2815 : _GEN_2655; // @[executor.scala 308:60]
  wire [7:0] _GEN_2976 = 8'h0 < length_1 ? _GEN_2816 : _GEN_2656; // @[executor.scala 308:60]
  wire [7:0] _GEN_2977 = 8'h0 < length_1 ? _GEN_2817 : _GEN_2657; // @[executor.scala 308:60]
  wire [7:0] _GEN_2978 = 8'h0 < length_1 ? _GEN_2818 : _GEN_2658; // @[executor.scala 308:60]
  wire [7:0] _GEN_2979 = 8'h0 < length_1 ? _GEN_2819 : _GEN_2659; // @[executor.scala 308:60]
  wire [7:0] _GEN_2980 = 8'h0 < length_1 ? _GEN_2820 : _GEN_2660; // @[executor.scala 308:60]
  wire [7:0] _GEN_2981 = 8'h0 < length_1 ? _GEN_2821 : _GEN_2661; // @[executor.scala 308:60]
  wire [7:0] _GEN_2982 = 8'h0 < length_1 ? _GEN_2822 : _GEN_2662; // @[executor.scala 308:60]
  wire [7:0] _GEN_2983 = 8'h0 < length_1 ? _GEN_2823 : _GEN_2663; // @[executor.scala 308:60]
  wire [7:0] _GEN_2984 = 8'h0 < length_1 ? _GEN_2824 : _GEN_2664; // @[executor.scala 308:60]
  wire [7:0] _GEN_2985 = 8'h0 < length_1 ? _GEN_2825 : _GEN_2665; // @[executor.scala 308:60]
  wire [7:0] _GEN_2986 = 8'h0 < length_1 ? _GEN_2826 : _GEN_2666; // @[executor.scala 308:60]
  wire [7:0] _GEN_2987 = 8'h0 < length_1 ? _GEN_2827 : _GEN_2667; // @[executor.scala 308:60]
  wire [7:0] _GEN_2988 = 8'h0 < length_1 ? _GEN_2828 : _GEN_2668; // @[executor.scala 308:60]
  wire [7:0] _GEN_2989 = 8'h0 < length_1 ? _GEN_2829 : _GEN_2669; // @[executor.scala 308:60]
  wire [7:0] _GEN_2990 = 8'h0 < length_1 ? _GEN_2830 : _GEN_2670; // @[executor.scala 308:60]
  wire [7:0] _GEN_2991 = 8'h0 < length_1 ? _GEN_2831 : _GEN_2671; // @[executor.scala 308:60]
  wire [7:0] _GEN_2992 = 8'h0 < length_1 ? _GEN_2832 : _GEN_2672; // @[executor.scala 308:60]
  wire [7:0] _GEN_2993 = 8'h0 < length_1 ? _GEN_2833 : _GEN_2673; // @[executor.scala 308:60]
  wire [7:0] _GEN_2994 = 8'h0 < length_1 ? _GEN_2834 : _GEN_2674; // @[executor.scala 308:60]
  wire [7:0] _GEN_2995 = 8'h0 < length_1 ? _GEN_2835 : _GEN_2675; // @[executor.scala 308:60]
  wire [7:0] _GEN_2996 = 8'h0 < length_1 ? _GEN_2836 : _GEN_2676; // @[executor.scala 308:60]
  wire [7:0] _GEN_2997 = 8'h0 < length_1 ? _GEN_2837 : _GEN_2677; // @[executor.scala 308:60]
  wire [7:0] _GEN_2998 = 8'h0 < length_1 ? _GEN_2838 : _GEN_2678; // @[executor.scala 308:60]
  wire [7:0] _GEN_2999 = 8'h0 < length_1 ? _GEN_2839 : _GEN_2679; // @[executor.scala 308:60]
  wire [7:0] _GEN_3000 = 8'h0 < length_1 ? _GEN_2840 : _GEN_2680; // @[executor.scala 308:60]
  wire [7:0] _GEN_3001 = 8'h0 < length_1 ? _GEN_2841 : _GEN_2681; // @[executor.scala 308:60]
  wire [7:0] _GEN_3002 = 8'h0 < length_1 ? _GEN_2842 : _GEN_2682; // @[executor.scala 308:60]
  wire [7:0] _GEN_3003 = 8'h0 < length_1 ? _GEN_2843 : _GEN_2683; // @[executor.scala 308:60]
  wire [7:0] _GEN_3004 = 8'h0 < length_1 ? _GEN_2844 : _GEN_2684; // @[executor.scala 308:60]
  wire [7:0] _GEN_3005 = 8'h0 < length_1 ? _GEN_2845 : _GEN_2685; // @[executor.scala 308:60]
  wire [7:0] _GEN_3006 = 8'h0 < length_1 ? _GEN_2846 : _GEN_2686; // @[executor.scala 308:60]
  wire [7:0] _GEN_3007 = 8'h0 < length_1 ? _GEN_2847 : _GEN_2687; // @[executor.scala 308:60]
  wire [7:0] _GEN_3008 = 8'h0 < length_1 ? _GEN_2848 : _GEN_2688; // @[executor.scala 308:60]
  wire [7:0] _GEN_3009 = 8'h0 < length_1 ? _GEN_2849 : _GEN_2689; // @[executor.scala 308:60]
  wire [7:0] _GEN_3010 = 8'h0 < length_1 ? _GEN_2850 : _GEN_2690; // @[executor.scala 308:60]
  wire [7:0] _GEN_3011 = 8'h0 < length_1 ? _GEN_2851 : _GEN_2691; // @[executor.scala 308:60]
  wire [7:0] _GEN_3012 = 8'h0 < length_1 ? _GEN_2852 : _GEN_2692; // @[executor.scala 308:60]
  wire [7:0] _GEN_3013 = 8'h0 < length_1 ? _GEN_2853 : _GEN_2693; // @[executor.scala 308:60]
  wire [7:0] _GEN_3014 = 8'h0 < length_1 ? _GEN_2854 : _GEN_2694; // @[executor.scala 308:60]
  wire [7:0] _GEN_3015 = 8'h0 < length_1 ? _GEN_2855 : _GEN_2695; // @[executor.scala 308:60]
  wire [7:0] _GEN_3016 = 8'h0 < length_1 ? _GEN_2856 : _GEN_2696; // @[executor.scala 308:60]
  wire [7:0] _GEN_3017 = 8'h0 < length_1 ? _GEN_2857 : _GEN_2697; // @[executor.scala 308:60]
  wire [7:0] _GEN_3018 = 8'h0 < length_1 ? _GEN_2858 : _GEN_2698; // @[executor.scala 308:60]
  wire [7:0] _GEN_3019 = 8'h0 < length_1 ? _GEN_2859 : _GEN_2699; // @[executor.scala 308:60]
  wire [7:0] _GEN_3020 = 8'h0 < length_1 ? _GEN_2860 : _GEN_2700; // @[executor.scala 308:60]
  wire [7:0] _GEN_3021 = 8'h0 < length_1 ? _GEN_2861 : _GEN_2701; // @[executor.scala 308:60]
  wire [7:0] _GEN_3022 = 8'h0 < length_1 ? _GEN_2862 : _GEN_2702; // @[executor.scala 308:60]
  wire [7:0] _GEN_3023 = 8'h0 < length_1 ? _GEN_2863 : _GEN_2703; // @[executor.scala 308:60]
  wire [7:0] _GEN_3024 = 8'h0 < length_1 ? _GEN_2864 : _GEN_2704; // @[executor.scala 308:60]
  wire [7:0] _GEN_3025 = 8'h0 < length_1 ? _GEN_2865 : _GEN_2705; // @[executor.scala 308:60]
  wire [7:0] _GEN_3026 = 8'h0 < length_1 ? _GEN_2866 : _GEN_2706; // @[executor.scala 308:60]
  wire [7:0] _GEN_3027 = 8'h0 < length_1 ? _GEN_2867 : _GEN_2707; // @[executor.scala 308:60]
  wire [7:0] _GEN_3028 = 8'h0 < length_1 ? _GEN_2868 : _GEN_2708; // @[executor.scala 308:60]
  wire [7:0] _GEN_3029 = 8'h0 < length_1 ? _GEN_2869 : _GEN_2709; // @[executor.scala 308:60]
  wire [7:0] _GEN_3030 = 8'h0 < length_1 ? _GEN_2870 : _GEN_2710; // @[executor.scala 308:60]
  wire [7:0] _GEN_3031 = 8'h0 < length_1 ? _GEN_2871 : _GEN_2711; // @[executor.scala 308:60]
  wire [7:0] _GEN_3032 = 8'h0 < length_1 ? _GEN_2872 : _GEN_2712; // @[executor.scala 308:60]
  wire [7:0] _GEN_3033 = 8'h0 < length_1 ? _GEN_2873 : _GEN_2713; // @[executor.scala 308:60]
  wire [7:0] _GEN_3034 = 8'h0 < length_1 ? _GEN_2874 : _GEN_2714; // @[executor.scala 308:60]
  wire [7:0] _GEN_3035 = 8'h0 < length_1 ? _GEN_2875 : _GEN_2715; // @[executor.scala 308:60]
  wire [7:0] _GEN_3036 = 8'h0 < length_1 ? _GEN_2876 : _GEN_2716; // @[executor.scala 308:60]
  wire [7:0] _GEN_3037 = 8'h0 < length_1 ? _GEN_2877 : _GEN_2717; // @[executor.scala 308:60]
  wire [7:0] _GEN_3038 = 8'h0 < length_1 ? _GEN_2878 : _GEN_2718; // @[executor.scala 308:60]
  wire [7:0] _GEN_3039 = 8'h0 < length_1 ? _GEN_2879 : _GEN_2719; // @[executor.scala 308:60]
  wire [7:0] _GEN_3040 = 8'h0 < length_1 ? _GEN_2880 : _GEN_2720; // @[executor.scala 308:60]
  wire [7:0] _GEN_3041 = 8'h0 < length_1 ? _GEN_2881 : _GEN_2721; // @[executor.scala 308:60]
  wire [7:0] field_byte_9 = field_1[55:48]; // @[executor.scala 305:57]
  wire [7:0] total_offset_9 = offset_1 + 8'h1; // @[executor.scala 307:57]
  wire [7:0] _GEN_3042 = 8'h0 == total_offset_9 ? field_byte_9 : _GEN_2882; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3043 = 8'h1 == total_offset_9 ? field_byte_9 : _GEN_2883; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3044 = 8'h2 == total_offset_9 ? field_byte_9 : _GEN_2884; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3045 = 8'h3 == total_offset_9 ? field_byte_9 : _GEN_2885; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3046 = 8'h4 == total_offset_9 ? field_byte_9 : _GEN_2886; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3047 = 8'h5 == total_offset_9 ? field_byte_9 : _GEN_2887; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3048 = 8'h6 == total_offset_9 ? field_byte_9 : _GEN_2888; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3049 = 8'h7 == total_offset_9 ? field_byte_9 : _GEN_2889; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3050 = 8'h8 == total_offset_9 ? field_byte_9 : _GEN_2890; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3051 = 8'h9 == total_offset_9 ? field_byte_9 : _GEN_2891; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3052 = 8'ha == total_offset_9 ? field_byte_9 : _GEN_2892; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3053 = 8'hb == total_offset_9 ? field_byte_9 : _GEN_2893; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3054 = 8'hc == total_offset_9 ? field_byte_9 : _GEN_2894; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3055 = 8'hd == total_offset_9 ? field_byte_9 : _GEN_2895; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3056 = 8'he == total_offset_9 ? field_byte_9 : _GEN_2896; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3057 = 8'hf == total_offset_9 ? field_byte_9 : _GEN_2897; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3058 = 8'h10 == total_offset_9 ? field_byte_9 : _GEN_2898; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3059 = 8'h11 == total_offset_9 ? field_byte_9 : _GEN_2899; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3060 = 8'h12 == total_offset_9 ? field_byte_9 : _GEN_2900; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3061 = 8'h13 == total_offset_9 ? field_byte_9 : _GEN_2901; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3062 = 8'h14 == total_offset_9 ? field_byte_9 : _GEN_2902; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3063 = 8'h15 == total_offset_9 ? field_byte_9 : _GEN_2903; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3064 = 8'h16 == total_offset_9 ? field_byte_9 : _GEN_2904; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3065 = 8'h17 == total_offset_9 ? field_byte_9 : _GEN_2905; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3066 = 8'h18 == total_offset_9 ? field_byte_9 : _GEN_2906; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3067 = 8'h19 == total_offset_9 ? field_byte_9 : _GEN_2907; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3068 = 8'h1a == total_offset_9 ? field_byte_9 : _GEN_2908; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3069 = 8'h1b == total_offset_9 ? field_byte_9 : _GEN_2909; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3070 = 8'h1c == total_offset_9 ? field_byte_9 : _GEN_2910; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3071 = 8'h1d == total_offset_9 ? field_byte_9 : _GEN_2911; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3072 = 8'h1e == total_offset_9 ? field_byte_9 : _GEN_2912; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3073 = 8'h1f == total_offset_9 ? field_byte_9 : _GEN_2913; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3074 = 8'h20 == total_offset_9 ? field_byte_9 : _GEN_2914; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3075 = 8'h21 == total_offset_9 ? field_byte_9 : _GEN_2915; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3076 = 8'h22 == total_offset_9 ? field_byte_9 : _GEN_2916; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3077 = 8'h23 == total_offset_9 ? field_byte_9 : _GEN_2917; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3078 = 8'h24 == total_offset_9 ? field_byte_9 : _GEN_2918; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3079 = 8'h25 == total_offset_9 ? field_byte_9 : _GEN_2919; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3080 = 8'h26 == total_offset_9 ? field_byte_9 : _GEN_2920; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3081 = 8'h27 == total_offset_9 ? field_byte_9 : _GEN_2921; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3082 = 8'h28 == total_offset_9 ? field_byte_9 : _GEN_2922; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3083 = 8'h29 == total_offset_9 ? field_byte_9 : _GEN_2923; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3084 = 8'h2a == total_offset_9 ? field_byte_9 : _GEN_2924; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3085 = 8'h2b == total_offset_9 ? field_byte_9 : _GEN_2925; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3086 = 8'h2c == total_offset_9 ? field_byte_9 : _GEN_2926; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3087 = 8'h2d == total_offset_9 ? field_byte_9 : _GEN_2927; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3088 = 8'h2e == total_offset_9 ? field_byte_9 : _GEN_2928; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3089 = 8'h2f == total_offset_9 ? field_byte_9 : _GEN_2929; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3090 = 8'h30 == total_offset_9 ? field_byte_9 : _GEN_2930; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3091 = 8'h31 == total_offset_9 ? field_byte_9 : _GEN_2931; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3092 = 8'h32 == total_offset_9 ? field_byte_9 : _GEN_2932; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3093 = 8'h33 == total_offset_9 ? field_byte_9 : _GEN_2933; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3094 = 8'h34 == total_offset_9 ? field_byte_9 : _GEN_2934; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3095 = 8'h35 == total_offset_9 ? field_byte_9 : _GEN_2935; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3096 = 8'h36 == total_offset_9 ? field_byte_9 : _GEN_2936; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3097 = 8'h37 == total_offset_9 ? field_byte_9 : _GEN_2937; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3098 = 8'h38 == total_offset_9 ? field_byte_9 : _GEN_2938; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3099 = 8'h39 == total_offset_9 ? field_byte_9 : _GEN_2939; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3100 = 8'h3a == total_offset_9 ? field_byte_9 : _GEN_2940; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3101 = 8'h3b == total_offset_9 ? field_byte_9 : _GEN_2941; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3102 = 8'h3c == total_offset_9 ? field_byte_9 : _GEN_2942; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3103 = 8'h3d == total_offset_9 ? field_byte_9 : _GEN_2943; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3104 = 8'h3e == total_offset_9 ? field_byte_9 : _GEN_2944; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3105 = 8'h3f == total_offset_9 ? field_byte_9 : _GEN_2945; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3106 = 8'h40 == total_offset_9 ? field_byte_9 : _GEN_2946; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3107 = 8'h41 == total_offset_9 ? field_byte_9 : _GEN_2947; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3108 = 8'h42 == total_offset_9 ? field_byte_9 : _GEN_2948; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3109 = 8'h43 == total_offset_9 ? field_byte_9 : _GEN_2949; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3110 = 8'h44 == total_offset_9 ? field_byte_9 : _GEN_2950; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3111 = 8'h45 == total_offset_9 ? field_byte_9 : _GEN_2951; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3112 = 8'h46 == total_offset_9 ? field_byte_9 : _GEN_2952; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3113 = 8'h47 == total_offset_9 ? field_byte_9 : _GEN_2953; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3114 = 8'h48 == total_offset_9 ? field_byte_9 : _GEN_2954; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3115 = 8'h49 == total_offset_9 ? field_byte_9 : _GEN_2955; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3116 = 8'h4a == total_offset_9 ? field_byte_9 : _GEN_2956; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3117 = 8'h4b == total_offset_9 ? field_byte_9 : _GEN_2957; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3118 = 8'h4c == total_offset_9 ? field_byte_9 : _GEN_2958; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3119 = 8'h4d == total_offset_9 ? field_byte_9 : _GEN_2959; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3120 = 8'h4e == total_offset_9 ? field_byte_9 : _GEN_2960; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3121 = 8'h4f == total_offset_9 ? field_byte_9 : _GEN_2961; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3122 = 8'h50 == total_offset_9 ? field_byte_9 : _GEN_2962; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3123 = 8'h51 == total_offset_9 ? field_byte_9 : _GEN_2963; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3124 = 8'h52 == total_offset_9 ? field_byte_9 : _GEN_2964; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3125 = 8'h53 == total_offset_9 ? field_byte_9 : _GEN_2965; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3126 = 8'h54 == total_offset_9 ? field_byte_9 : _GEN_2966; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3127 = 8'h55 == total_offset_9 ? field_byte_9 : _GEN_2967; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3128 = 8'h56 == total_offset_9 ? field_byte_9 : _GEN_2968; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3129 = 8'h57 == total_offset_9 ? field_byte_9 : _GEN_2969; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3130 = 8'h58 == total_offset_9 ? field_byte_9 : _GEN_2970; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3131 = 8'h59 == total_offset_9 ? field_byte_9 : _GEN_2971; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3132 = 8'h5a == total_offset_9 ? field_byte_9 : _GEN_2972; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3133 = 8'h5b == total_offset_9 ? field_byte_9 : _GEN_2973; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3134 = 8'h5c == total_offset_9 ? field_byte_9 : _GEN_2974; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3135 = 8'h5d == total_offset_9 ? field_byte_9 : _GEN_2975; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3136 = 8'h5e == total_offset_9 ? field_byte_9 : _GEN_2976; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3137 = 8'h5f == total_offset_9 ? field_byte_9 : _GEN_2977; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3138 = 8'h60 == total_offset_9 ? field_byte_9 : _GEN_2978; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3139 = 8'h61 == total_offset_9 ? field_byte_9 : _GEN_2979; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3140 = 8'h62 == total_offset_9 ? field_byte_9 : _GEN_2980; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3141 = 8'h63 == total_offset_9 ? field_byte_9 : _GEN_2981; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3142 = 8'h64 == total_offset_9 ? field_byte_9 : _GEN_2982; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3143 = 8'h65 == total_offset_9 ? field_byte_9 : _GEN_2983; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3144 = 8'h66 == total_offset_9 ? field_byte_9 : _GEN_2984; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3145 = 8'h67 == total_offset_9 ? field_byte_9 : _GEN_2985; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3146 = 8'h68 == total_offset_9 ? field_byte_9 : _GEN_2986; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3147 = 8'h69 == total_offset_9 ? field_byte_9 : _GEN_2987; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3148 = 8'h6a == total_offset_9 ? field_byte_9 : _GEN_2988; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3149 = 8'h6b == total_offset_9 ? field_byte_9 : _GEN_2989; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3150 = 8'h6c == total_offset_9 ? field_byte_9 : _GEN_2990; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3151 = 8'h6d == total_offset_9 ? field_byte_9 : _GEN_2991; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3152 = 8'h6e == total_offset_9 ? field_byte_9 : _GEN_2992; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3153 = 8'h6f == total_offset_9 ? field_byte_9 : _GEN_2993; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3154 = 8'h70 == total_offset_9 ? field_byte_9 : _GEN_2994; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3155 = 8'h71 == total_offset_9 ? field_byte_9 : _GEN_2995; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3156 = 8'h72 == total_offset_9 ? field_byte_9 : _GEN_2996; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3157 = 8'h73 == total_offset_9 ? field_byte_9 : _GEN_2997; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3158 = 8'h74 == total_offset_9 ? field_byte_9 : _GEN_2998; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3159 = 8'h75 == total_offset_9 ? field_byte_9 : _GEN_2999; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3160 = 8'h76 == total_offset_9 ? field_byte_9 : _GEN_3000; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3161 = 8'h77 == total_offset_9 ? field_byte_9 : _GEN_3001; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3162 = 8'h78 == total_offset_9 ? field_byte_9 : _GEN_3002; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3163 = 8'h79 == total_offset_9 ? field_byte_9 : _GEN_3003; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3164 = 8'h7a == total_offset_9 ? field_byte_9 : _GEN_3004; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3165 = 8'h7b == total_offset_9 ? field_byte_9 : _GEN_3005; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3166 = 8'h7c == total_offset_9 ? field_byte_9 : _GEN_3006; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3167 = 8'h7d == total_offset_9 ? field_byte_9 : _GEN_3007; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3168 = 8'h7e == total_offset_9 ? field_byte_9 : _GEN_3008; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3169 = 8'h7f == total_offset_9 ? field_byte_9 : _GEN_3009; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3170 = 8'h80 == total_offset_9 ? field_byte_9 : _GEN_3010; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3171 = 8'h81 == total_offset_9 ? field_byte_9 : _GEN_3011; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3172 = 8'h82 == total_offset_9 ? field_byte_9 : _GEN_3012; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3173 = 8'h83 == total_offset_9 ? field_byte_9 : _GEN_3013; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3174 = 8'h84 == total_offset_9 ? field_byte_9 : _GEN_3014; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3175 = 8'h85 == total_offset_9 ? field_byte_9 : _GEN_3015; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3176 = 8'h86 == total_offset_9 ? field_byte_9 : _GEN_3016; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3177 = 8'h87 == total_offset_9 ? field_byte_9 : _GEN_3017; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3178 = 8'h88 == total_offset_9 ? field_byte_9 : _GEN_3018; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3179 = 8'h89 == total_offset_9 ? field_byte_9 : _GEN_3019; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3180 = 8'h8a == total_offset_9 ? field_byte_9 : _GEN_3020; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3181 = 8'h8b == total_offset_9 ? field_byte_9 : _GEN_3021; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3182 = 8'h8c == total_offset_9 ? field_byte_9 : _GEN_3022; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3183 = 8'h8d == total_offset_9 ? field_byte_9 : _GEN_3023; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3184 = 8'h8e == total_offset_9 ? field_byte_9 : _GEN_3024; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3185 = 8'h8f == total_offset_9 ? field_byte_9 : _GEN_3025; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3186 = 8'h90 == total_offset_9 ? field_byte_9 : _GEN_3026; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3187 = 8'h91 == total_offset_9 ? field_byte_9 : _GEN_3027; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3188 = 8'h92 == total_offset_9 ? field_byte_9 : _GEN_3028; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3189 = 8'h93 == total_offset_9 ? field_byte_9 : _GEN_3029; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3190 = 8'h94 == total_offset_9 ? field_byte_9 : _GEN_3030; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3191 = 8'h95 == total_offset_9 ? field_byte_9 : _GEN_3031; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3192 = 8'h96 == total_offset_9 ? field_byte_9 : _GEN_3032; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3193 = 8'h97 == total_offset_9 ? field_byte_9 : _GEN_3033; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3194 = 8'h98 == total_offset_9 ? field_byte_9 : _GEN_3034; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3195 = 8'h99 == total_offset_9 ? field_byte_9 : _GEN_3035; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3196 = 8'h9a == total_offset_9 ? field_byte_9 : _GEN_3036; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3197 = 8'h9b == total_offset_9 ? field_byte_9 : _GEN_3037; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3198 = 8'h9c == total_offset_9 ? field_byte_9 : _GEN_3038; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3199 = 8'h9d == total_offset_9 ? field_byte_9 : _GEN_3039; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3200 = 8'h9e == total_offset_9 ? field_byte_9 : _GEN_3040; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3201 = 8'h9f == total_offset_9 ? field_byte_9 : _GEN_3041; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3202 = 8'h1 < length_1 ? _GEN_3042 : _GEN_2882; // @[executor.scala 308:60]
  wire [7:0] _GEN_3203 = 8'h1 < length_1 ? _GEN_3043 : _GEN_2883; // @[executor.scala 308:60]
  wire [7:0] _GEN_3204 = 8'h1 < length_1 ? _GEN_3044 : _GEN_2884; // @[executor.scala 308:60]
  wire [7:0] _GEN_3205 = 8'h1 < length_1 ? _GEN_3045 : _GEN_2885; // @[executor.scala 308:60]
  wire [7:0] _GEN_3206 = 8'h1 < length_1 ? _GEN_3046 : _GEN_2886; // @[executor.scala 308:60]
  wire [7:0] _GEN_3207 = 8'h1 < length_1 ? _GEN_3047 : _GEN_2887; // @[executor.scala 308:60]
  wire [7:0] _GEN_3208 = 8'h1 < length_1 ? _GEN_3048 : _GEN_2888; // @[executor.scala 308:60]
  wire [7:0] _GEN_3209 = 8'h1 < length_1 ? _GEN_3049 : _GEN_2889; // @[executor.scala 308:60]
  wire [7:0] _GEN_3210 = 8'h1 < length_1 ? _GEN_3050 : _GEN_2890; // @[executor.scala 308:60]
  wire [7:0] _GEN_3211 = 8'h1 < length_1 ? _GEN_3051 : _GEN_2891; // @[executor.scala 308:60]
  wire [7:0] _GEN_3212 = 8'h1 < length_1 ? _GEN_3052 : _GEN_2892; // @[executor.scala 308:60]
  wire [7:0] _GEN_3213 = 8'h1 < length_1 ? _GEN_3053 : _GEN_2893; // @[executor.scala 308:60]
  wire [7:0] _GEN_3214 = 8'h1 < length_1 ? _GEN_3054 : _GEN_2894; // @[executor.scala 308:60]
  wire [7:0] _GEN_3215 = 8'h1 < length_1 ? _GEN_3055 : _GEN_2895; // @[executor.scala 308:60]
  wire [7:0] _GEN_3216 = 8'h1 < length_1 ? _GEN_3056 : _GEN_2896; // @[executor.scala 308:60]
  wire [7:0] _GEN_3217 = 8'h1 < length_1 ? _GEN_3057 : _GEN_2897; // @[executor.scala 308:60]
  wire [7:0] _GEN_3218 = 8'h1 < length_1 ? _GEN_3058 : _GEN_2898; // @[executor.scala 308:60]
  wire [7:0] _GEN_3219 = 8'h1 < length_1 ? _GEN_3059 : _GEN_2899; // @[executor.scala 308:60]
  wire [7:0] _GEN_3220 = 8'h1 < length_1 ? _GEN_3060 : _GEN_2900; // @[executor.scala 308:60]
  wire [7:0] _GEN_3221 = 8'h1 < length_1 ? _GEN_3061 : _GEN_2901; // @[executor.scala 308:60]
  wire [7:0] _GEN_3222 = 8'h1 < length_1 ? _GEN_3062 : _GEN_2902; // @[executor.scala 308:60]
  wire [7:0] _GEN_3223 = 8'h1 < length_1 ? _GEN_3063 : _GEN_2903; // @[executor.scala 308:60]
  wire [7:0] _GEN_3224 = 8'h1 < length_1 ? _GEN_3064 : _GEN_2904; // @[executor.scala 308:60]
  wire [7:0] _GEN_3225 = 8'h1 < length_1 ? _GEN_3065 : _GEN_2905; // @[executor.scala 308:60]
  wire [7:0] _GEN_3226 = 8'h1 < length_1 ? _GEN_3066 : _GEN_2906; // @[executor.scala 308:60]
  wire [7:0] _GEN_3227 = 8'h1 < length_1 ? _GEN_3067 : _GEN_2907; // @[executor.scala 308:60]
  wire [7:0] _GEN_3228 = 8'h1 < length_1 ? _GEN_3068 : _GEN_2908; // @[executor.scala 308:60]
  wire [7:0] _GEN_3229 = 8'h1 < length_1 ? _GEN_3069 : _GEN_2909; // @[executor.scala 308:60]
  wire [7:0] _GEN_3230 = 8'h1 < length_1 ? _GEN_3070 : _GEN_2910; // @[executor.scala 308:60]
  wire [7:0] _GEN_3231 = 8'h1 < length_1 ? _GEN_3071 : _GEN_2911; // @[executor.scala 308:60]
  wire [7:0] _GEN_3232 = 8'h1 < length_1 ? _GEN_3072 : _GEN_2912; // @[executor.scala 308:60]
  wire [7:0] _GEN_3233 = 8'h1 < length_1 ? _GEN_3073 : _GEN_2913; // @[executor.scala 308:60]
  wire [7:0] _GEN_3234 = 8'h1 < length_1 ? _GEN_3074 : _GEN_2914; // @[executor.scala 308:60]
  wire [7:0] _GEN_3235 = 8'h1 < length_1 ? _GEN_3075 : _GEN_2915; // @[executor.scala 308:60]
  wire [7:0] _GEN_3236 = 8'h1 < length_1 ? _GEN_3076 : _GEN_2916; // @[executor.scala 308:60]
  wire [7:0] _GEN_3237 = 8'h1 < length_1 ? _GEN_3077 : _GEN_2917; // @[executor.scala 308:60]
  wire [7:0] _GEN_3238 = 8'h1 < length_1 ? _GEN_3078 : _GEN_2918; // @[executor.scala 308:60]
  wire [7:0] _GEN_3239 = 8'h1 < length_1 ? _GEN_3079 : _GEN_2919; // @[executor.scala 308:60]
  wire [7:0] _GEN_3240 = 8'h1 < length_1 ? _GEN_3080 : _GEN_2920; // @[executor.scala 308:60]
  wire [7:0] _GEN_3241 = 8'h1 < length_1 ? _GEN_3081 : _GEN_2921; // @[executor.scala 308:60]
  wire [7:0] _GEN_3242 = 8'h1 < length_1 ? _GEN_3082 : _GEN_2922; // @[executor.scala 308:60]
  wire [7:0] _GEN_3243 = 8'h1 < length_1 ? _GEN_3083 : _GEN_2923; // @[executor.scala 308:60]
  wire [7:0] _GEN_3244 = 8'h1 < length_1 ? _GEN_3084 : _GEN_2924; // @[executor.scala 308:60]
  wire [7:0] _GEN_3245 = 8'h1 < length_1 ? _GEN_3085 : _GEN_2925; // @[executor.scala 308:60]
  wire [7:0] _GEN_3246 = 8'h1 < length_1 ? _GEN_3086 : _GEN_2926; // @[executor.scala 308:60]
  wire [7:0] _GEN_3247 = 8'h1 < length_1 ? _GEN_3087 : _GEN_2927; // @[executor.scala 308:60]
  wire [7:0] _GEN_3248 = 8'h1 < length_1 ? _GEN_3088 : _GEN_2928; // @[executor.scala 308:60]
  wire [7:0] _GEN_3249 = 8'h1 < length_1 ? _GEN_3089 : _GEN_2929; // @[executor.scala 308:60]
  wire [7:0] _GEN_3250 = 8'h1 < length_1 ? _GEN_3090 : _GEN_2930; // @[executor.scala 308:60]
  wire [7:0] _GEN_3251 = 8'h1 < length_1 ? _GEN_3091 : _GEN_2931; // @[executor.scala 308:60]
  wire [7:0] _GEN_3252 = 8'h1 < length_1 ? _GEN_3092 : _GEN_2932; // @[executor.scala 308:60]
  wire [7:0] _GEN_3253 = 8'h1 < length_1 ? _GEN_3093 : _GEN_2933; // @[executor.scala 308:60]
  wire [7:0] _GEN_3254 = 8'h1 < length_1 ? _GEN_3094 : _GEN_2934; // @[executor.scala 308:60]
  wire [7:0] _GEN_3255 = 8'h1 < length_1 ? _GEN_3095 : _GEN_2935; // @[executor.scala 308:60]
  wire [7:0] _GEN_3256 = 8'h1 < length_1 ? _GEN_3096 : _GEN_2936; // @[executor.scala 308:60]
  wire [7:0] _GEN_3257 = 8'h1 < length_1 ? _GEN_3097 : _GEN_2937; // @[executor.scala 308:60]
  wire [7:0] _GEN_3258 = 8'h1 < length_1 ? _GEN_3098 : _GEN_2938; // @[executor.scala 308:60]
  wire [7:0] _GEN_3259 = 8'h1 < length_1 ? _GEN_3099 : _GEN_2939; // @[executor.scala 308:60]
  wire [7:0] _GEN_3260 = 8'h1 < length_1 ? _GEN_3100 : _GEN_2940; // @[executor.scala 308:60]
  wire [7:0] _GEN_3261 = 8'h1 < length_1 ? _GEN_3101 : _GEN_2941; // @[executor.scala 308:60]
  wire [7:0] _GEN_3262 = 8'h1 < length_1 ? _GEN_3102 : _GEN_2942; // @[executor.scala 308:60]
  wire [7:0] _GEN_3263 = 8'h1 < length_1 ? _GEN_3103 : _GEN_2943; // @[executor.scala 308:60]
  wire [7:0] _GEN_3264 = 8'h1 < length_1 ? _GEN_3104 : _GEN_2944; // @[executor.scala 308:60]
  wire [7:0] _GEN_3265 = 8'h1 < length_1 ? _GEN_3105 : _GEN_2945; // @[executor.scala 308:60]
  wire [7:0] _GEN_3266 = 8'h1 < length_1 ? _GEN_3106 : _GEN_2946; // @[executor.scala 308:60]
  wire [7:0] _GEN_3267 = 8'h1 < length_1 ? _GEN_3107 : _GEN_2947; // @[executor.scala 308:60]
  wire [7:0] _GEN_3268 = 8'h1 < length_1 ? _GEN_3108 : _GEN_2948; // @[executor.scala 308:60]
  wire [7:0] _GEN_3269 = 8'h1 < length_1 ? _GEN_3109 : _GEN_2949; // @[executor.scala 308:60]
  wire [7:0] _GEN_3270 = 8'h1 < length_1 ? _GEN_3110 : _GEN_2950; // @[executor.scala 308:60]
  wire [7:0] _GEN_3271 = 8'h1 < length_1 ? _GEN_3111 : _GEN_2951; // @[executor.scala 308:60]
  wire [7:0] _GEN_3272 = 8'h1 < length_1 ? _GEN_3112 : _GEN_2952; // @[executor.scala 308:60]
  wire [7:0] _GEN_3273 = 8'h1 < length_1 ? _GEN_3113 : _GEN_2953; // @[executor.scala 308:60]
  wire [7:0] _GEN_3274 = 8'h1 < length_1 ? _GEN_3114 : _GEN_2954; // @[executor.scala 308:60]
  wire [7:0] _GEN_3275 = 8'h1 < length_1 ? _GEN_3115 : _GEN_2955; // @[executor.scala 308:60]
  wire [7:0] _GEN_3276 = 8'h1 < length_1 ? _GEN_3116 : _GEN_2956; // @[executor.scala 308:60]
  wire [7:0] _GEN_3277 = 8'h1 < length_1 ? _GEN_3117 : _GEN_2957; // @[executor.scala 308:60]
  wire [7:0] _GEN_3278 = 8'h1 < length_1 ? _GEN_3118 : _GEN_2958; // @[executor.scala 308:60]
  wire [7:0] _GEN_3279 = 8'h1 < length_1 ? _GEN_3119 : _GEN_2959; // @[executor.scala 308:60]
  wire [7:0] _GEN_3280 = 8'h1 < length_1 ? _GEN_3120 : _GEN_2960; // @[executor.scala 308:60]
  wire [7:0] _GEN_3281 = 8'h1 < length_1 ? _GEN_3121 : _GEN_2961; // @[executor.scala 308:60]
  wire [7:0] _GEN_3282 = 8'h1 < length_1 ? _GEN_3122 : _GEN_2962; // @[executor.scala 308:60]
  wire [7:0] _GEN_3283 = 8'h1 < length_1 ? _GEN_3123 : _GEN_2963; // @[executor.scala 308:60]
  wire [7:0] _GEN_3284 = 8'h1 < length_1 ? _GEN_3124 : _GEN_2964; // @[executor.scala 308:60]
  wire [7:0] _GEN_3285 = 8'h1 < length_1 ? _GEN_3125 : _GEN_2965; // @[executor.scala 308:60]
  wire [7:0] _GEN_3286 = 8'h1 < length_1 ? _GEN_3126 : _GEN_2966; // @[executor.scala 308:60]
  wire [7:0] _GEN_3287 = 8'h1 < length_1 ? _GEN_3127 : _GEN_2967; // @[executor.scala 308:60]
  wire [7:0] _GEN_3288 = 8'h1 < length_1 ? _GEN_3128 : _GEN_2968; // @[executor.scala 308:60]
  wire [7:0] _GEN_3289 = 8'h1 < length_1 ? _GEN_3129 : _GEN_2969; // @[executor.scala 308:60]
  wire [7:0] _GEN_3290 = 8'h1 < length_1 ? _GEN_3130 : _GEN_2970; // @[executor.scala 308:60]
  wire [7:0] _GEN_3291 = 8'h1 < length_1 ? _GEN_3131 : _GEN_2971; // @[executor.scala 308:60]
  wire [7:0] _GEN_3292 = 8'h1 < length_1 ? _GEN_3132 : _GEN_2972; // @[executor.scala 308:60]
  wire [7:0] _GEN_3293 = 8'h1 < length_1 ? _GEN_3133 : _GEN_2973; // @[executor.scala 308:60]
  wire [7:0] _GEN_3294 = 8'h1 < length_1 ? _GEN_3134 : _GEN_2974; // @[executor.scala 308:60]
  wire [7:0] _GEN_3295 = 8'h1 < length_1 ? _GEN_3135 : _GEN_2975; // @[executor.scala 308:60]
  wire [7:0] _GEN_3296 = 8'h1 < length_1 ? _GEN_3136 : _GEN_2976; // @[executor.scala 308:60]
  wire [7:0] _GEN_3297 = 8'h1 < length_1 ? _GEN_3137 : _GEN_2977; // @[executor.scala 308:60]
  wire [7:0] _GEN_3298 = 8'h1 < length_1 ? _GEN_3138 : _GEN_2978; // @[executor.scala 308:60]
  wire [7:0] _GEN_3299 = 8'h1 < length_1 ? _GEN_3139 : _GEN_2979; // @[executor.scala 308:60]
  wire [7:0] _GEN_3300 = 8'h1 < length_1 ? _GEN_3140 : _GEN_2980; // @[executor.scala 308:60]
  wire [7:0] _GEN_3301 = 8'h1 < length_1 ? _GEN_3141 : _GEN_2981; // @[executor.scala 308:60]
  wire [7:0] _GEN_3302 = 8'h1 < length_1 ? _GEN_3142 : _GEN_2982; // @[executor.scala 308:60]
  wire [7:0] _GEN_3303 = 8'h1 < length_1 ? _GEN_3143 : _GEN_2983; // @[executor.scala 308:60]
  wire [7:0] _GEN_3304 = 8'h1 < length_1 ? _GEN_3144 : _GEN_2984; // @[executor.scala 308:60]
  wire [7:0] _GEN_3305 = 8'h1 < length_1 ? _GEN_3145 : _GEN_2985; // @[executor.scala 308:60]
  wire [7:0] _GEN_3306 = 8'h1 < length_1 ? _GEN_3146 : _GEN_2986; // @[executor.scala 308:60]
  wire [7:0] _GEN_3307 = 8'h1 < length_1 ? _GEN_3147 : _GEN_2987; // @[executor.scala 308:60]
  wire [7:0] _GEN_3308 = 8'h1 < length_1 ? _GEN_3148 : _GEN_2988; // @[executor.scala 308:60]
  wire [7:0] _GEN_3309 = 8'h1 < length_1 ? _GEN_3149 : _GEN_2989; // @[executor.scala 308:60]
  wire [7:0] _GEN_3310 = 8'h1 < length_1 ? _GEN_3150 : _GEN_2990; // @[executor.scala 308:60]
  wire [7:0] _GEN_3311 = 8'h1 < length_1 ? _GEN_3151 : _GEN_2991; // @[executor.scala 308:60]
  wire [7:0] _GEN_3312 = 8'h1 < length_1 ? _GEN_3152 : _GEN_2992; // @[executor.scala 308:60]
  wire [7:0] _GEN_3313 = 8'h1 < length_1 ? _GEN_3153 : _GEN_2993; // @[executor.scala 308:60]
  wire [7:0] _GEN_3314 = 8'h1 < length_1 ? _GEN_3154 : _GEN_2994; // @[executor.scala 308:60]
  wire [7:0] _GEN_3315 = 8'h1 < length_1 ? _GEN_3155 : _GEN_2995; // @[executor.scala 308:60]
  wire [7:0] _GEN_3316 = 8'h1 < length_1 ? _GEN_3156 : _GEN_2996; // @[executor.scala 308:60]
  wire [7:0] _GEN_3317 = 8'h1 < length_1 ? _GEN_3157 : _GEN_2997; // @[executor.scala 308:60]
  wire [7:0] _GEN_3318 = 8'h1 < length_1 ? _GEN_3158 : _GEN_2998; // @[executor.scala 308:60]
  wire [7:0] _GEN_3319 = 8'h1 < length_1 ? _GEN_3159 : _GEN_2999; // @[executor.scala 308:60]
  wire [7:0] _GEN_3320 = 8'h1 < length_1 ? _GEN_3160 : _GEN_3000; // @[executor.scala 308:60]
  wire [7:0] _GEN_3321 = 8'h1 < length_1 ? _GEN_3161 : _GEN_3001; // @[executor.scala 308:60]
  wire [7:0] _GEN_3322 = 8'h1 < length_1 ? _GEN_3162 : _GEN_3002; // @[executor.scala 308:60]
  wire [7:0] _GEN_3323 = 8'h1 < length_1 ? _GEN_3163 : _GEN_3003; // @[executor.scala 308:60]
  wire [7:0] _GEN_3324 = 8'h1 < length_1 ? _GEN_3164 : _GEN_3004; // @[executor.scala 308:60]
  wire [7:0] _GEN_3325 = 8'h1 < length_1 ? _GEN_3165 : _GEN_3005; // @[executor.scala 308:60]
  wire [7:0] _GEN_3326 = 8'h1 < length_1 ? _GEN_3166 : _GEN_3006; // @[executor.scala 308:60]
  wire [7:0] _GEN_3327 = 8'h1 < length_1 ? _GEN_3167 : _GEN_3007; // @[executor.scala 308:60]
  wire [7:0] _GEN_3328 = 8'h1 < length_1 ? _GEN_3168 : _GEN_3008; // @[executor.scala 308:60]
  wire [7:0] _GEN_3329 = 8'h1 < length_1 ? _GEN_3169 : _GEN_3009; // @[executor.scala 308:60]
  wire [7:0] _GEN_3330 = 8'h1 < length_1 ? _GEN_3170 : _GEN_3010; // @[executor.scala 308:60]
  wire [7:0] _GEN_3331 = 8'h1 < length_1 ? _GEN_3171 : _GEN_3011; // @[executor.scala 308:60]
  wire [7:0] _GEN_3332 = 8'h1 < length_1 ? _GEN_3172 : _GEN_3012; // @[executor.scala 308:60]
  wire [7:0] _GEN_3333 = 8'h1 < length_1 ? _GEN_3173 : _GEN_3013; // @[executor.scala 308:60]
  wire [7:0] _GEN_3334 = 8'h1 < length_1 ? _GEN_3174 : _GEN_3014; // @[executor.scala 308:60]
  wire [7:0] _GEN_3335 = 8'h1 < length_1 ? _GEN_3175 : _GEN_3015; // @[executor.scala 308:60]
  wire [7:0] _GEN_3336 = 8'h1 < length_1 ? _GEN_3176 : _GEN_3016; // @[executor.scala 308:60]
  wire [7:0] _GEN_3337 = 8'h1 < length_1 ? _GEN_3177 : _GEN_3017; // @[executor.scala 308:60]
  wire [7:0] _GEN_3338 = 8'h1 < length_1 ? _GEN_3178 : _GEN_3018; // @[executor.scala 308:60]
  wire [7:0] _GEN_3339 = 8'h1 < length_1 ? _GEN_3179 : _GEN_3019; // @[executor.scala 308:60]
  wire [7:0] _GEN_3340 = 8'h1 < length_1 ? _GEN_3180 : _GEN_3020; // @[executor.scala 308:60]
  wire [7:0] _GEN_3341 = 8'h1 < length_1 ? _GEN_3181 : _GEN_3021; // @[executor.scala 308:60]
  wire [7:0] _GEN_3342 = 8'h1 < length_1 ? _GEN_3182 : _GEN_3022; // @[executor.scala 308:60]
  wire [7:0] _GEN_3343 = 8'h1 < length_1 ? _GEN_3183 : _GEN_3023; // @[executor.scala 308:60]
  wire [7:0] _GEN_3344 = 8'h1 < length_1 ? _GEN_3184 : _GEN_3024; // @[executor.scala 308:60]
  wire [7:0] _GEN_3345 = 8'h1 < length_1 ? _GEN_3185 : _GEN_3025; // @[executor.scala 308:60]
  wire [7:0] _GEN_3346 = 8'h1 < length_1 ? _GEN_3186 : _GEN_3026; // @[executor.scala 308:60]
  wire [7:0] _GEN_3347 = 8'h1 < length_1 ? _GEN_3187 : _GEN_3027; // @[executor.scala 308:60]
  wire [7:0] _GEN_3348 = 8'h1 < length_1 ? _GEN_3188 : _GEN_3028; // @[executor.scala 308:60]
  wire [7:0] _GEN_3349 = 8'h1 < length_1 ? _GEN_3189 : _GEN_3029; // @[executor.scala 308:60]
  wire [7:0] _GEN_3350 = 8'h1 < length_1 ? _GEN_3190 : _GEN_3030; // @[executor.scala 308:60]
  wire [7:0] _GEN_3351 = 8'h1 < length_1 ? _GEN_3191 : _GEN_3031; // @[executor.scala 308:60]
  wire [7:0] _GEN_3352 = 8'h1 < length_1 ? _GEN_3192 : _GEN_3032; // @[executor.scala 308:60]
  wire [7:0] _GEN_3353 = 8'h1 < length_1 ? _GEN_3193 : _GEN_3033; // @[executor.scala 308:60]
  wire [7:0] _GEN_3354 = 8'h1 < length_1 ? _GEN_3194 : _GEN_3034; // @[executor.scala 308:60]
  wire [7:0] _GEN_3355 = 8'h1 < length_1 ? _GEN_3195 : _GEN_3035; // @[executor.scala 308:60]
  wire [7:0] _GEN_3356 = 8'h1 < length_1 ? _GEN_3196 : _GEN_3036; // @[executor.scala 308:60]
  wire [7:0] _GEN_3357 = 8'h1 < length_1 ? _GEN_3197 : _GEN_3037; // @[executor.scala 308:60]
  wire [7:0] _GEN_3358 = 8'h1 < length_1 ? _GEN_3198 : _GEN_3038; // @[executor.scala 308:60]
  wire [7:0] _GEN_3359 = 8'h1 < length_1 ? _GEN_3199 : _GEN_3039; // @[executor.scala 308:60]
  wire [7:0] _GEN_3360 = 8'h1 < length_1 ? _GEN_3200 : _GEN_3040; // @[executor.scala 308:60]
  wire [7:0] _GEN_3361 = 8'h1 < length_1 ? _GEN_3201 : _GEN_3041; // @[executor.scala 308:60]
  wire [7:0] field_byte_10 = field_1[47:40]; // @[executor.scala 305:57]
  wire [7:0] total_offset_10 = offset_1 + 8'h2; // @[executor.scala 307:57]
  wire [7:0] _GEN_3362 = 8'h0 == total_offset_10 ? field_byte_10 : _GEN_3202; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3363 = 8'h1 == total_offset_10 ? field_byte_10 : _GEN_3203; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3364 = 8'h2 == total_offset_10 ? field_byte_10 : _GEN_3204; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3365 = 8'h3 == total_offset_10 ? field_byte_10 : _GEN_3205; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3366 = 8'h4 == total_offset_10 ? field_byte_10 : _GEN_3206; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3367 = 8'h5 == total_offset_10 ? field_byte_10 : _GEN_3207; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3368 = 8'h6 == total_offset_10 ? field_byte_10 : _GEN_3208; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3369 = 8'h7 == total_offset_10 ? field_byte_10 : _GEN_3209; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3370 = 8'h8 == total_offset_10 ? field_byte_10 : _GEN_3210; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3371 = 8'h9 == total_offset_10 ? field_byte_10 : _GEN_3211; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3372 = 8'ha == total_offset_10 ? field_byte_10 : _GEN_3212; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3373 = 8'hb == total_offset_10 ? field_byte_10 : _GEN_3213; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3374 = 8'hc == total_offset_10 ? field_byte_10 : _GEN_3214; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3375 = 8'hd == total_offset_10 ? field_byte_10 : _GEN_3215; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3376 = 8'he == total_offset_10 ? field_byte_10 : _GEN_3216; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3377 = 8'hf == total_offset_10 ? field_byte_10 : _GEN_3217; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3378 = 8'h10 == total_offset_10 ? field_byte_10 : _GEN_3218; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3379 = 8'h11 == total_offset_10 ? field_byte_10 : _GEN_3219; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3380 = 8'h12 == total_offset_10 ? field_byte_10 : _GEN_3220; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3381 = 8'h13 == total_offset_10 ? field_byte_10 : _GEN_3221; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3382 = 8'h14 == total_offset_10 ? field_byte_10 : _GEN_3222; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3383 = 8'h15 == total_offset_10 ? field_byte_10 : _GEN_3223; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3384 = 8'h16 == total_offset_10 ? field_byte_10 : _GEN_3224; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3385 = 8'h17 == total_offset_10 ? field_byte_10 : _GEN_3225; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3386 = 8'h18 == total_offset_10 ? field_byte_10 : _GEN_3226; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3387 = 8'h19 == total_offset_10 ? field_byte_10 : _GEN_3227; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3388 = 8'h1a == total_offset_10 ? field_byte_10 : _GEN_3228; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3389 = 8'h1b == total_offset_10 ? field_byte_10 : _GEN_3229; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3390 = 8'h1c == total_offset_10 ? field_byte_10 : _GEN_3230; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3391 = 8'h1d == total_offset_10 ? field_byte_10 : _GEN_3231; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3392 = 8'h1e == total_offset_10 ? field_byte_10 : _GEN_3232; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3393 = 8'h1f == total_offset_10 ? field_byte_10 : _GEN_3233; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3394 = 8'h20 == total_offset_10 ? field_byte_10 : _GEN_3234; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3395 = 8'h21 == total_offset_10 ? field_byte_10 : _GEN_3235; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3396 = 8'h22 == total_offset_10 ? field_byte_10 : _GEN_3236; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3397 = 8'h23 == total_offset_10 ? field_byte_10 : _GEN_3237; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3398 = 8'h24 == total_offset_10 ? field_byte_10 : _GEN_3238; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3399 = 8'h25 == total_offset_10 ? field_byte_10 : _GEN_3239; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3400 = 8'h26 == total_offset_10 ? field_byte_10 : _GEN_3240; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3401 = 8'h27 == total_offset_10 ? field_byte_10 : _GEN_3241; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3402 = 8'h28 == total_offset_10 ? field_byte_10 : _GEN_3242; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3403 = 8'h29 == total_offset_10 ? field_byte_10 : _GEN_3243; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3404 = 8'h2a == total_offset_10 ? field_byte_10 : _GEN_3244; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3405 = 8'h2b == total_offset_10 ? field_byte_10 : _GEN_3245; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3406 = 8'h2c == total_offset_10 ? field_byte_10 : _GEN_3246; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3407 = 8'h2d == total_offset_10 ? field_byte_10 : _GEN_3247; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3408 = 8'h2e == total_offset_10 ? field_byte_10 : _GEN_3248; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3409 = 8'h2f == total_offset_10 ? field_byte_10 : _GEN_3249; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3410 = 8'h30 == total_offset_10 ? field_byte_10 : _GEN_3250; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3411 = 8'h31 == total_offset_10 ? field_byte_10 : _GEN_3251; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3412 = 8'h32 == total_offset_10 ? field_byte_10 : _GEN_3252; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3413 = 8'h33 == total_offset_10 ? field_byte_10 : _GEN_3253; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3414 = 8'h34 == total_offset_10 ? field_byte_10 : _GEN_3254; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3415 = 8'h35 == total_offset_10 ? field_byte_10 : _GEN_3255; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3416 = 8'h36 == total_offset_10 ? field_byte_10 : _GEN_3256; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3417 = 8'h37 == total_offset_10 ? field_byte_10 : _GEN_3257; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3418 = 8'h38 == total_offset_10 ? field_byte_10 : _GEN_3258; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3419 = 8'h39 == total_offset_10 ? field_byte_10 : _GEN_3259; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3420 = 8'h3a == total_offset_10 ? field_byte_10 : _GEN_3260; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3421 = 8'h3b == total_offset_10 ? field_byte_10 : _GEN_3261; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3422 = 8'h3c == total_offset_10 ? field_byte_10 : _GEN_3262; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3423 = 8'h3d == total_offset_10 ? field_byte_10 : _GEN_3263; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3424 = 8'h3e == total_offset_10 ? field_byte_10 : _GEN_3264; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3425 = 8'h3f == total_offset_10 ? field_byte_10 : _GEN_3265; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3426 = 8'h40 == total_offset_10 ? field_byte_10 : _GEN_3266; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3427 = 8'h41 == total_offset_10 ? field_byte_10 : _GEN_3267; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3428 = 8'h42 == total_offset_10 ? field_byte_10 : _GEN_3268; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3429 = 8'h43 == total_offset_10 ? field_byte_10 : _GEN_3269; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3430 = 8'h44 == total_offset_10 ? field_byte_10 : _GEN_3270; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3431 = 8'h45 == total_offset_10 ? field_byte_10 : _GEN_3271; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3432 = 8'h46 == total_offset_10 ? field_byte_10 : _GEN_3272; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3433 = 8'h47 == total_offset_10 ? field_byte_10 : _GEN_3273; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3434 = 8'h48 == total_offset_10 ? field_byte_10 : _GEN_3274; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3435 = 8'h49 == total_offset_10 ? field_byte_10 : _GEN_3275; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3436 = 8'h4a == total_offset_10 ? field_byte_10 : _GEN_3276; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3437 = 8'h4b == total_offset_10 ? field_byte_10 : _GEN_3277; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3438 = 8'h4c == total_offset_10 ? field_byte_10 : _GEN_3278; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3439 = 8'h4d == total_offset_10 ? field_byte_10 : _GEN_3279; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3440 = 8'h4e == total_offset_10 ? field_byte_10 : _GEN_3280; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3441 = 8'h4f == total_offset_10 ? field_byte_10 : _GEN_3281; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3442 = 8'h50 == total_offset_10 ? field_byte_10 : _GEN_3282; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3443 = 8'h51 == total_offset_10 ? field_byte_10 : _GEN_3283; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3444 = 8'h52 == total_offset_10 ? field_byte_10 : _GEN_3284; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3445 = 8'h53 == total_offset_10 ? field_byte_10 : _GEN_3285; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3446 = 8'h54 == total_offset_10 ? field_byte_10 : _GEN_3286; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3447 = 8'h55 == total_offset_10 ? field_byte_10 : _GEN_3287; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3448 = 8'h56 == total_offset_10 ? field_byte_10 : _GEN_3288; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3449 = 8'h57 == total_offset_10 ? field_byte_10 : _GEN_3289; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3450 = 8'h58 == total_offset_10 ? field_byte_10 : _GEN_3290; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3451 = 8'h59 == total_offset_10 ? field_byte_10 : _GEN_3291; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3452 = 8'h5a == total_offset_10 ? field_byte_10 : _GEN_3292; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3453 = 8'h5b == total_offset_10 ? field_byte_10 : _GEN_3293; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3454 = 8'h5c == total_offset_10 ? field_byte_10 : _GEN_3294; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3455 = 8'h5d == total_offset_10 ? field_byte_10 : _GEN_3295; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3456 = 8'h5e == total_offset_10 ? field_byte_10 : _GEN_3296; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3457 = 8'h5f == total_offset_10 ? field_byte_10 : _GEN_3297; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3458 = 8'h60 == total_offset_10 ? field_byte_10 : _GEN_3298; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3459 = 8'h61 == total_offset_10 ? field_byte_10 : _GEN_3299; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3460 = 8'h62 == total_offset_10 ? field_byte_10 : _GEN_3300; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3461 = 8'h63 == total_offset_10 ? field_byte_10 : _GEN_3301; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3462 = 8'h64 == total_offset_10 ? field_byte_10 : _GEN_3302; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3463 = 8'h65 == total_offset_10 ? field_byte_10 : _GEN_3303; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3464 = 8'h66 == total_offset_10 ? field_byte_10 : _GEN_3304; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3465 = 8'h67 == total_offset_10 ? field_byte_10 : _GEN_3305; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3466 = 8'h68 == total_offset_10 ? field_byte_10 : _GEN_3306; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3467 = 8'h69 == total_offset_10 ? field_byte_10 : _GEN_3307; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3468 = 8'h6a == total_offset_10 ? field_byte_10 : _GEN_3308; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3469 = 8'h6b == total_offset_10 ? field_byte_10 : _GEN_3309; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3470 = 8'h6c == total_offset_10 ? field_byte_10 : _GEN_3310; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3471 = 8'h6d == total_offset_10 ? field_byte_10 : _GEN_3311; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3472 = 8'h6e == total_offset_10 ? field_byte_10 : _GEN_3312; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3473 = 8'h6f == total_offset_10 ? field_byte_10 : _GEN_3313; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3474 = 8'h70 == total_offset_10 ? field_byte_10 : _GEN_3314; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3475 = 8'h71 == total_offset_10 ? field_byte_10 : _GEN_3315; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3476 = 8'h72 == total_offset_10 ? field_byte_10 : _GEN_3316; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3477 = 8'h73 == total_offset_10 ? field_byte_10 : _GEN_3317; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3478 = 8'h74 == total_offset_10 ? field_byte_10 : _GEN_3318; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3479 = 8'h75 == total_offset_10 ? field_byte_10 : _GEN_3319; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3480 = 8'h76 == total_offset_10 ? field_byte_10 : _GEN_3320; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3481 = 8'h77 == total_offset_10 ? field_byte_10 : _GEN_3321; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3482 = 8'h78 == total_offset_10 ? field_byte_10 : _GEN_3322; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3483 = 8'h79 == total_offset_10 ? field_byte_10 : _GEN_3323; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3484 = 8'h7a == total_offset_10 ? field_byte_10 : _GEN_3324; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3485 = 8'h7b == total_offset_10 ? field_byte_10 : _GEN_3325; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3486 = 8'h7c == total_offset_10 ? field_byte_10 : _GEN_3326; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3487 = 8'h7d == total_offset_10 ? field_byte_10 : _GEN_3327; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3488 = 8'h7e == total_offset_10 ? field_byte_10 : _GEN_3328; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3489 = 8'h7f == total_offset_10 ? field_byte_10 : _GEN_3329; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3490 = 8'h80 == total_offset_10 ? field_byte_10 : _GEN_3330; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3491 = 8'h81 == total_offset_10 ? field_byte_10 : _GEN_3331; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3492 = 8'h82 == total_offset_10 ? field_byte_10 : _GEN_3332; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3493 = 8'h83 == total_offset_10 ? field_byte_10 : _GEN_3333; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3494 = 8'h84 == total_offset_10 ? field_byte_10 : _GEN_3334; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3495 = 8'h85 == total_offset_10 ? field_byte_10 : _GEN_3335; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3496 = 8'h86 == total_offset_10 ? field_byte_10 : _GEN_3336; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3497 = 8'h87 == total_offset_10 ? field_byte_10 : _GEN_3337; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3498 = 8'h88 == total_offset_10 ? field_byte_10 : _GEN_3338; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3499 = 8'h89 == total_offset_10 ? field_byte_10 : _GEN_3339; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3500 = 8'h8a == total_offset_10 ? field_byte_10 : _GEN_3340; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3501 = 8'h8b == total_offset_10 ? field_byte_10 : _GEN_3341; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3502 = 8'h8c == total_offset_10 ? field_byte_10 : _GEN_3342; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3503 = 8'h8d == total_offset_10 ? field_byte_10 : _GEN_3343; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3504 = 8'h8e == total_offset_10 ? field_byte_10 : _GEN_3344; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3505 = 8'h8f == total_offset_10 ? field_byte_10 : _GEN_3345; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3506 = 8'h90 == total_offset_10 ? field_byte_10 : _GEN_3346; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3507 = 8'h91 == total_offset_10 ? field_byte_10 : _GEN_3347; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3508 = 8'h92 == total_offset_10 ? field_byte_10 : _GEN_3348; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3509 = 8'h93 == total_offset_10 ? field_byte_10 : _GEN_3349; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3510 = 8'h94 == total_offset_10 ? field_byte_10 : _GEN_3350; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3511 = 8'h95 == total_offset_10 ? field_byte_10 : _GEN_3351; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3512 = 8'h96 == total_offset_10 ? field_byte_10 : _GEN_3352; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3513 = 8'h97 == total_offset_10 ? field_byte_10 : _GEN_3353; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3514 = 8'h98 == total_offset_10 ? field_byte_10 : _GEN_3354; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3515 = 8'h99 == total_offset_10 ? field_byte_10 : _GEN_3355; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3516 = 8'h9a == total_offset_10 ? field_byte_10 : _GEN_3356; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3517 = 8'h9b == total_offset_10 ? field_byte_10 : _GEN_3357; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3518 = 8'h9c == total_offset_10 ? field_byte_10 : _GEN_3358; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3519 = 8'h9d == total_offset_10 ? field_byte_10 : _GEN_3359; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3520 = 8'h9e == total_offset_10 ? field_byte_10 : _GEN_3360; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3521 = 8'h9f == total_offset_10 ? field_byte_10 : _GEN_3361; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3522 = 8'h2 < length_1 ? _GEN_3362 : _GEN_3202; // @[executor.scala 308:60]
  wire [7:0] _GEN_3523 = 8'h2 < length_1 ? _GEN_3363 : _GEN_3203; // @[executor.scala 308:60]
  wire [7:0] _GEN_3524 = 8'h2 < length_1 ? _GEN_3364 : _GEN_3204; // @[executor.scala 308:60]
  wire [7:0] _GEN_3525 = 8'h2 < length_1 ? _GEN_3365 : _GEN_3205; // @[executor.scala 308:60]
  wire [7:0] _GEN_3526 = 8'h2 < length_1 ? _GEN_3366 : _GEN_3206; // @[executor.scala 308:60]
  wire [7:0] _GEN_3527 = 8'h2 < length_1 ? _GEN_3367 : _GEN_3207; // @[executor.scala 308:60]
  wire [7:0] _GEN_3528 = 8'h2 < length_1 ? _GEN_3368 : _GEN_3208; // @[executor.scala 308:60]
  wire [7:0] _GEN_3529 = 8'h2 < length_1 ? _GEN_3369 : _GEN_3209; // @[executor.scala 308:60]
  wire [7:0] _GEN_3530 = 8'h2 < length_1 ? _GEN_3370 : _GEN_3210; // @[executor.scala 308:60]
  wire [7:0] _GEN_3531 = 8'h2 < length_1 ? _GEN_3371 : _GEN_3211; // @[executor.scala 308:60]
  wire [7:0] _GEN_3532 = 8'h2 < length_1 ? _GEN_3372 : _GEN_3212; // @[executor.scala 308:60]
  wire [7:0] _GEN_3533 = 8'h2 < length_1 ? _GEN_3373 : _GEN_3213; // @[executor.scala 308:60]
  wire [7:0] _GEN_3534 = 8'h2 < length_1 ? _GEN_3374 : _GEN_3214; // @[executor.scala 308:60]
  wire [7:0] _GEN_3535 = 8'h2 < length_1 ? _GEN_3375 : _GEN_3215; // @[executor.scala 308:60]
  wire [7:0] _GEN_3536 = 8'h2 < length_1 ? _GEN_3376 : _GEN_3216; // @[executor.scala 308:60]
  wire [7:0] _GEN_3537 = 8'h2 < length_1 ? _GEN_3377 : _GEN_3217; // @[executor.scala 308:60]
  wire [7:0] _GEN_3538 = 8'h2 < length_1 ? _GEN_3378 : _GEN_3218; // @[executor.scala 308:60]
  wire [7:0] _GEN_3539 = 8'h2 < length_1 ? _GEN_3379 : _GEN_3219; // @[executor.scala 308:60]
  wire [7:0] _GEN_3540 = 8'h2 < length_1 ? _GEN_3380 : _GEN_3220; // @[executor.scala 308:60]
  wire [7:0] _GEN_3541 = 8'h2 < length_1 ? _GEN_3381 : _GEN_3221; // @[executor.scala 308:60]
  wire [7:0] _GEN_3542 = 8'h2 < length_1 ? _GEN_3382 : _GEN_3222; // @[executor.scala 308:60]
  wire [7:0] _GEN_3543 = 8'h2 < length_1 ? _GEN_3383 : _GEN_3223; // @[executor.scala 308:60]
  wire [7:0] _GEN_3544 = 8'h2 < length_1 ? _GEN_3384 : _GEN_3224; // @[executor.scala 308:60]
  wire [7:0] _GEN_3545 = 8'h2 < length_1 ? _GEN_3385 : _GEN_3225; // @[executor.scala 308:60]
  wire [7:0] _GEN_3546 = 8'h2 < length_1 ? _GEN_3386 : _GEN_3226; // @[executor.scala 308:60]
  wire [7:0] _GEN_3547 = 8'h2 < length_1 ? _GEN_3387 : _GEN_3227; // @[executor.scala 308:60]
  wire [7:0] _GEN_3548 = 8'h2 < length_1 ? _GEN_3388 : _GEN_3228; // @[executor.scala 308:60]
  wire [7:0] _GEN_3549 = 8'h2 < length_1 ? _GEN_3389 : _GEN_3229; // @[executor.scala 308:60]
  wire [7:0] _GEN_3550 = 8'h2 < length_1 ? _GEN_3390 : _GEN_3230; // @[executor.scala 308:60]
  wire [7:0] _GEN_3551 = 8'h2 < length_1 ? _GEN_3391 : _GEN_3231; // @[executor.scala 308:60]
  wire [7:0] _GEN_3552 = 8'h2 < length_1 ? _GEN_3392 : _GEN_3232; // @[executor.scala 308:60]
  wire [7:0] _GEN_3553 = 8'h2 < length_1 ? _GEN_3393 : _GEN_3233; // @[executor.scala 308:60]
  wire [7:0] _GEN_3554 = 8'h2 < length_1 ? _GEN_3394 : _GEN_3234; // @[executor.scala 308:60]
  wire [7:0] _GEN_3555 = 8'h2 < length_1 ? _GEN_3395 : _GEN_3235; // @[executor.scala 308:60]
  wire [7:0] _GEN_3556 = 8'h2 < length_1 ? _GEN_3396 : _GEN_3236; // @[executor.scala 308:60]
  wire [7:0] _GEN_3557 = 8'h2 < length_1 ? _GEN_3397 : _GEN_3237; // @[executor.scala 308:60]
  wire [7:0] _GEN_3558 = 8'h2 < length_1 ? _GEN_3398 : _GEN_3238; // @[executor.scala 308:60]
  wire [7:0] _GEN_3559 = 8'h2 < length_1 ? _GEN_3399 : _GEN_3239; // @[executor.scala 308:60]
  wire [7:0] _GEN_3560 = 8'h2 < length_1 ? _GEN_3400 : _GEN_3240; // @[executor.scala 308:60]
  wire [7:0] _GEN_3561 = 8'h2 < length_1 ? _GEN_3401 : _GEN_3241; // @[executor.scala 308:60]
  wire [7:0] _GEN_3562 = 8'h2 < length_1 ? _GEN_3402 : _GEN_3242; // @[executor.scala 308:60]
  wire [7:0] _GEN_3563 = 8'h2 < length_1 ? _GEN_3403 : _GEN_3243; // @[executor.scala 308:60]
  wire [7:0] _GEN_3564 = 8'h2 < length_1 ? _GEN_3404 : _GEN_3244; // @[executor.scala 308:60]
  wire [7:0] _GEN_3565 = 8'h2 < length_1 ? _GEN_3405 : _GEN_3245; // @[executor.scala 308:60]
  wire [7:0] _GEN_3566 = 8'h2 < length_1 ? _GEN_3406 : _GEN_3246; // @[executor.scala 308:60]
  wire [7:0] _GEN_3567 = 8'h2 < length_1 ? _GEN_3407 : _GEN_3247; // @[executor.scala 308:60]
  wire [7:0] _GEN_3568 = 8'h2 < length_1 ? _GEN_3408 : _GEN_3248; // @[executor.scala 308:60]
  wire [7:0] _GEN_3569 = 8'h2 < length_1 ? _GEN_3409 : _GEN_3249; // @[executor.scala 308:60]
  wire [7:0] _GEN_3570 = 8'h2 < length_1 ? _GEN_3410 : _GEN_3250; // @[executor.scala 308:60]
  wire [7:0] _GEN_3571 = 8'h2 < length_1 ? _GEN_3411 : _GEN_3251; // @[executor.scala 308:60]
  wire [7:0] _GEN_3572 = 8'h2 < length_1 ? _GEN_3412 : _GEN_3252; // @[executor.scala 308:60]
  wire [7:0] _GEN_3573 = 8'h2 < length_1 ? _GEN_3413 : _GEN_3253; // @[executor.scala 308:60]
  wire [7:0] _GEN_3574 = 8'h2 < length_1 ? _GEN_3414 : _GEN_3254; // @[executor.scala 308:60]
  wire [7:0] _GEN_3575 = 8'h2 < length_1 ? _GEN_3415 : _GEN_3255; // @[executor.scala 308:60]
  wire [7:0] _GEN_3576 = 8'h2 < length_1 ? _GEN_3416 : _GEN_3256; // @[executor.scala 308:60]
  wire [7:0] _GEN_3577 = 8'h2 < length_1 ? _GEN_3417 : _GEN_3257; // @[executor.scala 308:60]
  wire [7:0] _GEN_3578 = 8'h2 < length_1 ? _GEN_3418 : _GEN_3258; // @[executor.scala 308:60]
  wire [7:0] _GEN_3579 = 8'h2 < length_1 ? _GEN_3419 : _GEN_3259; // @[executor.scala 308:60]
  wire [7:0] _GEN_3580 = 8'h2 < length_1 ? _GEN_3420 : _GEN_3260; // @[executor.scala 308:60]
  wire [7:0] _GEN_3581 = 8'h2 < length_1 ? _GEN_3421 : _GEN_3261; // @[executor.scala 308:60]
  wire [7:0] _GEN_3582 = 8'h2 < length_1 ? _GEN_3422 : _GEN_3262; // @[executor.scala 308:60]
  wire [7:0] _GEN_3583 = 8'h2 < length_1 ? _GEN_3423 : _GEN_3263; // @[executor.scala 308:60]
  wire [7:0] _GEN_3584 = 8'h2 < length_1 ? _GEN_3424 : _GEN_3264; // @[executor.scala 308:60]
  wire [7:0] _GEN_3585 = 8'h2 < length_1 ? _GEN_3425 : _GEN_3265; // @[executor.scala 308:60]
  wire [7:0] _GEN_3586 = 8'h2 < length_1 ? _GEN_3426 : _GEN_3266; // @[executor.scala 308:60]
  wire [7:0] _GEN_3587 = 8'h2 < length_1 ? _GEN_3427 : _GEN_3267; // @[executor.scala 308:60]
  wire [7:0] _GEN_3588 = 8'h2 < length_1 ? _GEN_3428 : _GEN_3268; // @[executor.scala 308:60]
  wire [7:0] _GEN_3589 = 8'h2 < length_1 ? _GEN_3429 : _GEN_3269; // @[executor.scala 308:60]
  wire [7:0] _GEN_3590 = 8'h2 < length_1 ? _GEN_3430 : _GEN_3270; // @[executor.scala 308:60]
  wire [7:0] _GEN_3591 = 8'h2 < length_1 ? _GEN_3431 : _GEN_3271; // @[executor.scala 308:60]
  wire [7:0] _GEN_3592 = 8'h2 < length_1 ? _GEN_3432 : _GEN_3272; // @[executor.scala 308:60]
  wire [7:0] _GEN_3593 = 8'h2 < length_1 ? _GEN_3433 : _GEN_3273; // @[executor.scala 308:60]
  wire [7:0] _GEN_3594 = 8'h2 < length_1 ? _GEN_3434 : _GEN_3274; // @[executor.scala 308:60]
  wire [7:0] _GEN_3595 = 8'h2 < length_1 ? _GEN_3435 : _GEN_3275; // @[executor.scala 308:60]
  wire [7:0] _GEN_3596 = 8'h2 < length_1 ? _GEN_3436 : _GEN_3276; // @[executor.scala 308:60]
  wire [7:0] _GEN_3597 = 8'h2 < length_1 ? _GEN_3437 : _GEN_3277; // @[executor.scala 308:60]
  wire [7:0] _GEN_3598 = 8'h2 < length_1 ? _GEN_3438 : _GEN_3278; // @[executor.scala 308:60]
  wire [7:0] _GEN_3599 = 8'h2 < length_1 ? _GEN_3439 : _GEN_3279; // @[executor.scala 308:60]
  wire [7:0] _GEN_3600 = 8'h2 < length_1 ? _GEN_3440 : _GEN_3280; // @[executor.scala 308:60]
  wire [7:0] _GEN_3601 = 8'h2 < length_1 ? _GEN_3441 : _GEN_3281; // @[executor.scala 308:60]
  wire [7:0] _GEN_3602 = 8'h2 < length_1 ? _GEN_3442 : _GEN_3282; // @[executor.scala 308:60]
  wire [7:0] _GEN_3603 = 8'h2 < length_1 ? _GEN_3443 : _GEN_3283; // @[executor.scala 308:60]
  wire [7:0] _GEN_3604 = 8'h2 < length_1 ? _GEN_3444 : _GEN_3284; // @[executor.scala 308:60]
  wire [7:0] _GEN_3605 = 8'h2 < length_1 ? _GEN_3445 : _GEN_3285; // @[executor.scala 308:60]
  wire [7:0] _GEN_3606 = 8'h2 < length_1 ? _GEN_3446 : _GEN_3286; // @[executor.scala 308:60]
  wire [7:0] _GEN_3607 = 8'h2 < length_1 ? _GEN_3447 : _GEN_3287; // @[executor.scala 308:60]
  wire [7:0] _GEN_3608 = 8'h2 < length_1 ? _GEN_3448 : _GEN_3288; // @[executor.scala 308:60]
  wire [7:0] _GEN_3609 = 8'h2 < length_1 ? _GEN_3449 : _GEN_3289; // @[executor.scala 308:60]
  wire [7:0] _GEN_3610 = 8'h2 < length_1 ? _GEN_3450 : _GEN_3290; // @[executor.scala 308:60]
  wire [7:0] _GEN_3611 = 8'h2 < length_1 ? _GEN_3451 : _GEN_3291; // @[executor.scala 308:60]
  wire [7:0] _GEN_3612 = 8'h2 < length_1 ? _GEN_3452 : _GEN_3292; // @[executor.scala 308:60]
  wire [7:0] _GEN_3613 = 8'h2 < length_1 ? _GEN_3453 : _GEN_3293; // @[executor.scala 308:60]
  wire [7:0] _GEN_3614 = 8'h2 < length_1 ? _GEN_3454 : _GEN_3294; // @[executor.scala 308:60]
  wire [7:0] _GEN_3615 = 8'h2 < length_1 ? _GEN_3455 : _GEN_3295; // @[executor.scala 308:60]
  wire [7:0] _GEN_3616 = 8'h2 < length_1 ? _GEN_3456 : _GEN_3296; // @[executor.scala 308:60]
  wire [7:0] _GEN_3617 = 8'h2 < length_1 ? _GEN_3457 : _GEN_3297; // @[executor.scala 308:60]
  wire [7:0] _GEN_3618 = 8'h2 < length_1 ? _GEN_3458 : _GEN_3298; // @[executor.scala 308:60]
  wire [7:0] _GEN_3619 = 8'h2 < length_1 ? _GEN_3459 : _GEN_3299; // @[executor.scala 308:60]
  wire [7:0] _GEN_3620 = 8'h2 < length_1 ? _GEN_3460 : _GEN_3300; // @[executor.scala 308:60]
  wire [7:0] _GEN_3621 = 8'h2 < length_1 ? _GEN_3461 : _GEN_3301; // @[executor.scala 308:60]
  wire [7:0] _GEN_3622 = 8'h2 < length_1 ? _GEN_3462 : _GEN_3302; // @[executor.scala 308:60]
  wire [7:0] _GEN_3623 = 8'h2 < length_1 ? _GEN_3463 : _GEN_3303; // @[executor.scala 308:60]
  wire [7:0] _GEN_3624 = 8'h2 < length_1 ? _GEN_3464 : _GEN_3304; // @[executor.scala 308:60]
  wire [7:0] _GEN_3625 = 8'h2 < length_1 ? _GEN_3465 : _GEN_3305; // @[executor.scala 308:60]
  wire [7:0] _GEN_3626 = 8'h2 < length_1 ? _GEN_3466 : _GEN_3306; // @[executor.scala 308:60]
  wire [7:0] _GEN_3627 = 8'h2 < length_1 ? _GEN_3467 : _GEN_3307; // @[executor.scala 308:60]
  wire [7:0] _GEN_3628 = 8'h2 < length_1 ? _GEN_3468 : _GEN_3308; // @[executor.scala 308:60]
  wire [7:0] _GEN_3629 = 8'h2 < length_1 ? _GEN_3469 : _GEN_3309; // @[executor.scala 308:60]
  wire [7:0] _GEN_3630 = 8'h2 < length_1 ? _GEN_3470 : _GEN_3310; // @[executor.scala 308:60]
  wire [7:0] _GEN_3631 = 8'h2 < length_1 ? _GEN_3471 : _GEN_3311; // @[executor.scala 308:60]
  wire [7:0] _GEN_3632 = 8'h2 < length_1 ? _GEN_3472 : _GEN_3312; // @[executor.scala 308:60]
  wire [7:0] _GEN_3633 = 8'h2 < length_1 ? _GEN_3473 : _GEN_3313; // @[executor.scala 308:60]
  wire [7:0] _GEN_3634 = 8'h2 < length_1 ? _GEN_3474 : _GEN_3314; // @[executor.scala 308:60]
  wire [7:0] _GEN_3635 = 8'h2 < length_1 ? _GEN_3475 : _GEN_3315; // @[executor.scala 308:60]
  wire [7:0] _GEN_3636 = 8'h2 < length_1 ? _GEN_3476 : _GEN_3316; // @[executor.scala 308:60]
  wire [7:0] _GEN_3637 = 8'h2 < length_1 ? _GEN_3477 : _GEN_3317; // @[executor.scala 308:60]
  wire [7:0] _GEN_3638 = 8'h2 < length_1 ? _GEN_3478 : _GEN_3318; // @[executor.scala 308:60]
  wire [7:0] _GEN_3639 = 8'h2 < length_1 ? _GEN_3479 : _GEN_3319; // @[executor.scala 308:60]
  wire [7:0] _GEN_3640 = 8'h2 < length_1 ? _GEN_3480 : _GEN_3320; // @[executor.scala 308:60]
  wire [7:0] _GEN_3641 = 8'h2 < length_1 ? _GEN_3481 : _GEN_3321; // @[executor.scala 308:60]
  wire [7:0] _GEN_3642 = 8'h2 < length_1 ? _GEN_3482 : _GEN_3322; // @[executor.scala 308:60]
  wire [7:0] _GEN_3643 = 8'h2 < length_1 ? _GEN_3483 : _GEN_3323; // @[executor.scala 308:60]
  wire [7:0] _GEN_3644 = 8'h2 < length_1 ? _GEN_3484 : _GEN_3324; // @[executor.scala 308:60]
  wire [7:0] _GEN_3645 = 8'h2 < length_1 ? _GEN_3485 : _GEN_3325; // @[executor.scala 308:60]
  wire [7:0] _GEN_3646 = 8'h2 < length_1 ? _GEN_3486 : _GEN_3326; // @[executor.scala 308:60]
  wire [7:0] _GEN_3647 = 8'h2 < length_1 ? _GEN_3487 : _GEN_3327; // @[executor.scala 308:60]
  wire [7:0] _GEN_3648 = 8'h2 < length_1 ? _GEN_3488 : _GEN_3328; // @[executor.scala 308:60]
  wire [7:0] _GEN_3649 = 8'h2 < length_1 ? _GEN_3489 : _GEN_3329; // @[executor.scala 308:60]
  wire [7:0] _GEN_3650 = 8'h2 < length_1 ? _GEN_3490 : _GEN_3330; // @[executor.scala 308:60]
  wire [7:0] _GEN_3651 = 8'h2 < length_1 ? _GEN_3491 : _GEN_3331; // @[executor.scala 308:60]
  wire [7:0] _GEN_3652 = 8'h2 < length_1 ? _GEN_3492 : _GEN_3332; // @[executor.scala 308:60]
  wire [7:0] _GEN_3653 = 8'h2 < length_1 ? _GEN_3493 : _GEN_3333; // @[executor.scala 308:60]
  wire [7:0] _GEN_3654 = 8'h2 < length_1 ? _GEN_3494 : _GEN_3334; // @[executor.scala 308:60]
  wire [7:0] _GEN_3655 = 8'h2 < length_1 ? _GEN_3495 : _GEN_3335; // @[executor.scala 308:60]
  wire [7:0] _GEN_3656 = 8'h2 < length_1 ? _GEN_3496 : _GEN_3336; // @[executor.scala 308:60]
  wire [7:0] _GEN_3657 = 8'h2 < length_1 ? _GEN_3497 : _GEN_3337; // @[executor.scala 308:60]
  wire [7:0] _GEN_3658 = 8'h2 < length_1 ? _GEN_3498 : _GEN_3338; // @[executor.scala 308:60]
  wire [7:0] _GEN_3659 = 8'h2 < length_1 ? _GEN_3499 : _GEN_3339; // @[executor.scala 308:60]
  wire [7:0] _GEN_3660 = 8'h2 < length_1 ? _GEN_3500 : _GEN_3340; // @[executor.scala 308:60]
  wire [7:0] _GEN_3661 = 8'h2 < length_1 ? _GEN_3501 : _GEN_3341; // @[executor.scala 308:60]
  wire [7:0] _GEN_3662 = 8'h2 < length_1 ? _GEN_3502 : _GEN_3342; // @[executor.scala 308:60]
  wire [7:0] _GEN_3663 = 8'h2 < length_1 ? _GEN_3503 : _GEN_3343; // @[executor.scala 308:60]
  wire [7:0] _GEN_3664 = 8'h2 < length_1 ? _GEN_3504 : _GEN_3344; // @[executor.scala 308:60]
  wire [7:0] _GEN_3665 = 8'h2 < length_1 ? _GEN_3505 : _GEN_3345; // @[executor.scala 308:60]
  wire [7:0] _GEN_3666 = 8'h2 < length_1 ? _GEN_3506 : _GEN_3346; // @[executor.scala 308:60]
  wire [7:0] _GEN_3667 = 8'h2 < length_1 ? _GEN_3507 : _GEN_3347; // @[executor.scala 308:60]
  wire [7:0] _GEN_3668 = 8'h2 < length_1 ? _GEN_3508 : _GEN_3348; // @[executor.scala 308:60]
  wire [7:0] _GEN_3669 = 8'h2 < length_1 ? _GEN_3509 : _GEN_3349; // @[executor.scala 308:60]
  wire [7:0] _GEN_3670 = 8'h2 < length_1 ? _GEN_3510 : _GEN_3350; // @[executor.scala 308:60]
  wire [7:0] _GEN_3671 = 8'h2 < length_1 ? _GEN_3511 : _GEN_3351; // @[executor.scala 308:60]
  wire [7:0] _GEN_3672 = 8'h2 < length_1 ? _GEN_3512 : _GEN_3352; // @[executor.scala 308:60]
  wire [7:0] _GEN_3673 = 8'h2 < length_1 ? _GEN_3513 : _GEN_3353; // @[executor.scala 308:60]
  wire [7:0] _GEN_3674 = 8'h2 < length_1 ? _GEN_3514 : _GEN_3354; // @[executor.scala 308:60]
  wire [7:0] _GEN_3675 = 8'h2 < length_1 ? _GEN_3515 : _GEN_3355; // @[executor.scala 308:60]
  wire [7:0] _GEN_3676 = 8'h2 < length_1 ? _GEN_3516 : _GEN_3356; // @[executor.scala 308:60]
  wire [7:0] _GEN_3677 = 8'h2 < length_1 ? _GEN_3517 : _GEN_3357; // @[executor.scala 308:60]
  wire [7:0] _GEN_3678 = 8'h2 < length_1 ? _GEN_3518 : _GEN_3358; // @[executor.scala 308:60]
  wire [7:0] _GEN_3679 = 8'h2 < length_1 ? _GEN_3519 : _GEN_3359; // @[executor.scala 308:60]
  wire [7:0] _GEN_3680 = 8'h2 < length_1 ? _GEN_3520 : _GEN_3360; // @[executor.scala 308:60]
  wire [7:0] _GEN_3681 = 8'h2 < length_1 ? _GEN_3521 : _GEN_3361; // @[executor.scala 308:60]
  wire [7:0] field_byte_11 = field_1[39:32]; // @[executor.scala 305:57]
  wire [7:0] total_offset_11 = offset_1 + 8'h3; // @[executor.scala 307:57]
  wire [7:0] _GEN_3682 = 8'h0 == total_offset_11 ? field_byte_11 : _GEN_3522; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3683 = 8'h1 == total_offset_11 ? field_byte_11 : _GEN_3523; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3684 = 8'h2 == total_offset_11 ? field_byte_11 : _GEN_3524; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3685 = 8'h3 == total_offset_11 ? field_byte_11 : _GEN_3525; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3686 = 8'h4 == total_offset_11 ? field_byte_11 : _GEN_3526; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3687 = 8'h5 == total_offset_11 ? field_byte_11 : _GEN_3527; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3688 = 8'h6 == total_offset_11 ? field_byte_11 : _GEN_3528; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3689 = 8'h7 == total_offset_11 ? field_byte_11 : _GEN_3529; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3690 = 8'h8 == total_offset_11 ? field_byte_11 : _GEN_3530; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3691 = 8'h9 == total_offset_11 ? field_byte_11 : _GEN_3531; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3692 = 8'ha == total_offset_11 ? field_byte_11 : _GEN_3532; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3693 = 8'hb == total_offset_11 ? field_byte_11 : _GEN_3533; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3694 = 8'hc == total_offset_11 ? field_byte_11 : _GEN_3534; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3695 = 8'hd == total_offset_11 ? field_byte_11 : _GEN_3535; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3696 = 8'he == total_offset_11 ? field_byte_11 : _GEN_3536; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3697 = 8'hf == total_offset_11 ? field_byte_11 : _GEN_3537; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3698 = 8'h10 == total_offset_11 ? field_byte_11 : _GEN_3538; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3699 = 8'h11 == total_offset_11 ? field_byte_11 : _GEN_3539; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3700 = 8'h12 == total_offset_11 ? field_byte_11 : _GEN_3540; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3701 = 8'h13 == total_offset_11 ? field_byte_11 : _GEN_3541; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3702 = 8'h14 == total_offset_11 ? field_byte_11 : _GEN_3542; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3703 = 8'h15 == total_offset_11 ? field_byte_11 : _GEN_3543; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3704 = 8'h16 == total_offset_11 ? field_byte_11 : _GEN_3544; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3705 = 8'h17 == total_offset_11 ? field_byte_11 : _GEN_3545; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3706 = 8'h18 == total_offset_11 ? field_byte_11 : _GEN_3546; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3707 = 8'h19 == total_offset_11 ? field_byte_11 : _GEN_3547; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3708 = 8'h1a == total_offset_11 ? field_byte_11 : _GEN_3548; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3709 = 8'h1b == total_offset_11 ? field_byte_11 : _GEN_3549; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3710 = 8'h1c == total_offset_11 ? field_byte_11 : _GEN_3550; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3711 = 8'h1d == total_offset_11 ? field_byte_11 : _GEN_3551; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3712 = 8'h1e == total_offset_11 ? field_byte_11 : _GEN_3552; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3713 = 8'h1f == total_offset_11 ? field_byte_11 : _GEN_3553; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3714 = 8'h20 == total_offset_11 ? field_byte_11 : _GEN_3554; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3715 = 8'h21 == total_offset_11 ? field_byte_11 : _GEN_3555; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3716 = 8'h22 == total_offset_11 ? field_byte_11 : _GEN_3556; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3717 = 8'h23 == total_offset_11 ? field_byte_11 : _GEN_3557; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3718 = 8'h24 == total_offset_11 ? field_byte_11 : _GEN_3558; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3719 = 8'h25 == total_offset_11 ? field_byte_11 : _GEN_3559; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3720 = 8'h26 == total_offset_11 ? field_byte_11 : _GEN_3560; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3721 = 8'h27 == total_offset_11 ? field_byte_11 : _GEN_3561; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3722 = 8'h28 == total_offset_11 ? field_byte_11 : _GEN_3562; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3723 = 8'h29 == total_offset_11 ? field_byte_11 : _GEN_3563; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3724 = 8'h2a == total_offset_11 ? field_byte_11 : _GEN_3564; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3725 = 8'h2b == total_offset_11 ? field_byte_11 : _GEN_3565; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3726 = 8'h2c == total_offset_11 ? field_byte_11 : _GEN_3566; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3727 = 8'h2d == total_offset_11 ? field_byte_11 : _GEN_3567; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3728 = 8'h2e == total_offset_11 ? field_byte_11 : _GEN_3568; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3729 = 8'h2f == total_offset_11 ? field_byte_11 : _GEN_3569; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3730 = 8'h30 == total_offset_11 ? field_byte_11 : _GEN_3570; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3731 = 8'h31 == total_offset_11 ? field_byte_11 : _GEN_3571; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3732 = 8'h32 == total_offset_11 ? field_byte_11 : _GEN_3572; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3733 = 8'h33 == total_offset_11 ? field_byte_11 : _GEN_3573; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3734 = 8'h34 == total_offset_11 ? field_byte_11 : _GEN_3574; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3735 = 8'h35 == total_offset_11 ? field_byte_11 : _GEN_3575; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3736 = 8'h36 == total_offset_11 ? field_byte_11 : _GEN_3576; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3737 = 8'h37 == total_offset_11 ? field_byte_11 : _GEN_3577; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3738 = 8'h38 == total_offset_11 ? field_byte_11 : _GEN_3578; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3739 = 8'h39 == total_offset_11 ? field_byte_11 : _GEN_3579; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3740 = 8'h3a == total_offset_11 ? field_byte_11 : _GEN_3580; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3741 = 8'h3b == total_offset_11 ? field_byte_11 : _GEN_3581; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3742 = 8'h3c == total_offset_11 ? field_byte_11 : _GEN_3582; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3743 = 8'h3d == total_offset_11 ? field_byte_11 : _GEN_3583; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3744 = 8'h3e == total_offset_11 ? field_byte_11 : _GEN_3584; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3745 = 8'h3f == total_offset_11 ? field_byte_11 : _GEN_3585; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3746 = 8'h40 == total_offset_11 ? field_byte_11 : _GEN_3586; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3747 = 8'h41 == total_offset_11 ? field_byte_11 : _GEN_3587; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3748 = 8'h42 == total_offset_11 ? field_byte_11 : _GEN_3588; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3749 = 8'h43 == total_offset_11 ? field_byte_11 : _GEN_3589; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3750 = 8'h44 == total_offset_11 ? field_byte_11 : _GEN_3590; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3751 = 8'h45 == total_offset_11 ? field_byte_11 : _GEN_3591; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3752 = 8'h46 == total_offset_11 ? field_byte_11 : _GEN_3592; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3753 = 8'h47 == total_offset_11 ? field_byte_11 : _GEN_3593; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3754 = 8'h48 == total_offset_11 ? field_byte_11 : _GEN_3594; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3755 = 8'h49 == total_offset_11 ? field_byte_11 : _GEN_3595; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3756 = 8'h4a == total_offset_11 ? field_byte_11 : _GEN_3596; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3757 = 8'h4b == total_offset_11 ? field_byte_11 : _GEN_3597; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3758 = 8'h4c == total_offset_11 ? field_byte_11 : _GEN_3598; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3759 = 8'h4d == total_offset_11 ? field_byte_11 : _GEN_3599; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3760 = 8'h4e == total_offset_11 ? field_byte_11 : _GEN_3600; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3761 = 8'h4f == total_offset_11 ? field_byte_11 : _GEN_3601; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3762 = 8'h50 == total_offset_11 ? field_byte_11 : _GEN_3602; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3763 = 8'h51 == total_offset_11 ? field_byte_11 : _GEN_3603; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3764 = 8'h52 == total_offset_11 ? field_byte_11 : _GEN_3604; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3765 = 8'h53 == total_offset_11 ? field_byte_11 : _GEN_3605; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3766 = 8'h54 == total_offset_11 ? field_byte_11 : _GEN_3606; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3767 = 8'h55 == total_offset_11 ? field_byte_11 : _GEN_3607; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3768 = 8'h56 == total_offset_11 ? field_byte_11 : _GEN_3608; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3769 = 8'h57 == total_offset_11 ? field_byte_11 : _GEN_3609; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3770 = 8'h58 == total_offset_11 ? field_byte_11 : _GEN_3610; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3771 = 8'h59 == total_offset_11 ? field_byte_11 : _GEN_3611; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3772 = 8'h5a == total_offset_11 ? field_byte_11 : _GEN_3612; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3773 = 8'h5b == total_offset_11 ? field_byte_11 : _GEN_3613; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3774 = 8'h5c == total_offset_11 ? field_byte_11 : _GEN_3614; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3775 = 8'h5d == total_offset_11 ? field_byte_11 : _GEN_3615; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3776 = 8'h5e == total_offset_11 ? field_byte_11 : _GEN_3616; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3777 = 8'h5f == total_offset_11 ? field_byte_11 : _GEN_3617; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3778 = 8'h60 == total_offset_11 ? field_byte_11 : _GEN_3618; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3779 = 8'h61 == total_offset_11 ? field_byte_11 : _GEN_3619; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3780 = 8'h62 == total_offset_11 ? field_byte_11 : _GEN_3620; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3781 = 8'h63 == total_offset_11 ? field_byte_11 : _GEN_3621; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3782 = 8'h64 == total_offset_11 ? field_byte_11 : _GEN_3622; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3783 = 8'h65 == total_offset_11 ? field_byte_11 : _GEN_3623; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3784 = 8'h66 == total_offset_11 ? field_byte_11 : _GEN_3624; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3785 = 8'h67 == total_offset_11 ? field_byte_11 : _GEN_3625; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3786 = 8'h68 == total_offset_11 ? field_byte_11 : _GEN_3626; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3787 = 8'h69 == total_offset_11 ? field_byte_11 : _GEN_3627; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3788 = 8'h6a == total_offset_11 ? field_byte_11 : _GEN_3628; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3789 = 8'h6b == total_offset_11 ? field_byte_11 : _GEN_3629; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3790 = 8'h6c == total_offset_11 ? field_byte_11 : _GEN_3630; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3791 = 8'h6d == total_offset_11 ? field_byte_11 : _GEN_3631; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3792 = 8'h6e == total_offset_11 ? field_byte_11 : _GEN_3632; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3793 = 8'h6f == total_offset_11 ? field_byte_11 : _GEN_3633; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3794 = 8'h70 == total_offset_11 ? field_byte_11 : _GEN_3634; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3795 = 8'h71 == total_offset_11 ? field_byte_11 : _GEN_3635; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3796 = 8'h72 == total_offset_11 ? field_byte_11 : _GEN_3636; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3797 = 8'h73 == total_offset_11 ? field_byte_11 : _GEN_3637; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3798 = 8'h74 == total_offset_11 ? field_byte_11 : _GEN_3638; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3799 = 8'h75 == total_offset_11 ? field_byte_11 : _GEN_3639; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3800 = 8'h76 == total_offset_11 ? field_byte_11 : _GEN_3640; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3801 = 8'h77 == total_offset_11 ? field_byte_11 : _GEN_3641; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3802 = 8'h78 == total_offset_11 ? field_byte_11 : _GEN_3642; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3803 = 8'h79 == total_offset_11 ? field_byte_11 : _GEN_3643; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3804 = 8'h7a == total_offset_11 ? field_byte_11 : _GEN_3644; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3805 = 8'h7b == total_offset_11 ? field_byte_11 : _GEN_3645; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3806 = 8'h7c == total_offset_11 ? field_byte_11 : _GEN_3646; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3807 = 8'h7d == total_offset_11 ? field_byte_11 : _GEN_3647; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3808 = 8'h7e == total_offset_11 ? field_byte_11 : _GEN_3648; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3809 = 8'h7f == total_offset_11 ? field_byte_11 : _GEN_3649; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3810 = 8'h80 == total_offset_11 ? field_byte_11 : _GEN_3650; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3811 = 8'h81 == total_offset_11 ? field_byte_11 : _GEN_3651; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3812 = 8'h82 == total_offset_11 ? field_byte_11 : _GEN_3652; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3813 = 8'h83 == total_offset_11 ? field_byte_11 : _GEN_3653; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3814 = 8'h84 == total_offset_11 ? field_byte_11 : _GEN_3654; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3815 = 8'h85 == total_offset_11 ? field_byte_11 : _GEN_3655; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3816 = 8'h86 == total_offset_11 ? field_byte_11 : _GEN_3656; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3817 = 8'h87 == total_offset_11 ? field_byte_11 : _GEN_3657; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3818 = 8'h88 == total_offset_11 ? field_byte_11 : _GEN_3658; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3819 = 8'h89 == total_offset_11 ? field_byte_11 : _GEN_3659; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3820 = 8'h8a == total_offset_11 ? field_byte_11 : _GEN_3660; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3821 = 8'h8b == total_offset_11 ? field_byte_11 : _GEN_3661; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3822 = 8'h8c == total_offset_11 ? field_byte_11 : _GEN_3662; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3823 = 8'h8d == total_offset_11 ? field_byte_11 : _GEN_3663; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3824 = 8'h8e == total_offset_11 ? field_byte_11 : _GEN_3664; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3825 = 8'h8f == total_offset_11 ? field_byte_11 : _GEN_3665; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3826 = 8'h90 == total_offset_11 ? field_byte_11 : _GEN_3666; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3827 = 8'h91 == total_offset_11 ? field_byte_11 : _GEN_3667; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3828 = 8'h92 == total_offset_11 ? field_byte_11 : _GEN_3668; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3829 = 8'h93 == total_offset_11 ? field_byte_11 : _GEN_3669; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3830 = 8'h94 == total_offset_11 ? field_byte_11 : _GEN_3670; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3831 = 8'h95 == total_offset_11 ? field_byte_11 : _GEN_3671; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3832 = 8'h96 == total_offset_11 ? field_byte_11 : _GEN_3672; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3833 = 8'h97 == total_offset_11 ? field_byte_11 : _GEN_3673; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3834 = 8'h98 == total_offset_11 ? field_byte_11 : _GEN_3674; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3835 = 8'h99 == total_offset_11 ? field_byte_11 : _GEN_3675; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3836 = 8'h9a == total_offset_11 ? field_byte_11 : _GEN_3676; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3837 = 8'h9b == total_offset_11 ? field_byte_11 : _GEN_3677; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3838 = 8'h9c == total_offset_11 ? field_byte_11 : _GEN_3678; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3839 = 8'h9d == total_offset_11 ? field_byte_11 : _GEN_3679; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3840 = 8'h9e == total_offset_11 ? field_byte_11 : _GEN_3680; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3841 = 8'h9f == total_offset_11 ? field_byte_11 : _GEN_3681; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_3842 = 8'h3 < length_1 ? _GEN_3682 : _GEN_3522; // @[executor.scala 308:60]
  wire [7:0] _GEN_3843 = 8'h3 < length_1 ? _GEN_3683 : _GEN_3523; // @[executor.scala 308:60]
  wire [7:0] _GEN_3844 = 8'h3 < length_1 ? _GEN_3684 : _GEN_3524; // @[executor.scala 308:60]
  wire [7:0] _GEN_3845 = 8'h3 < length_1 ? _GEN_3685 : _GEN_3525; // @[executor.scala 308:60]
  wire [7:0] _GEN_3846 = 8'h3 < length_1 ? _GEN_3686 : _GEN_3526; // @[executor.scala 308:60]
  wire [7:0] _GEN_3847 = 8'h3 < length_1 ? _GEN_3687 : _GEN_3527; // @[executor.scala 308:60]
  wire [7:0] _GEN_3848 = 8'h3 < length_1 ? _GEN_3688 : _GEN_3528; // @[executor.scala 308:60]
  wire [7:0] _GEN_3849 = 8'h3 < length_1 ? _GEN_3689 : _GEN_3529; // @[executor.scala 308:60]
  wire [7:0] _GEN_3850 = 8'h3 < length_1 ? _GEN_3690 : _GEN_3530; // @[executor.scala 308:60]
  wire [7:0] _GEN_3851 = 8'h3 < length_1 ? _GEN_3691 : _GEN_3531; // @[executor.scala 308:60]
  wire [7:0] _GEN_3852 = 8'h3 < length_1 ? _GEN_3692 : _GEN_3532; // @[executor.scala 308:60]
  wire [7:0] _GEN_3853 = 8'h3 < length_1 ? _GEN_3693 : _GEN_3533; // @[executor.scala 308:60]
  wire [7:0] _GEN_3854 = 8'h3 < length_1 ? _GEN_3694 : _GEN_3534; // @[executor.scala 308:60]
  wire [7:0] _GEN_3855 = 8'h3 < length_1 ? _GEN_3695 : _GEN_3535; // @[executor.scala 308:60]
  wire [7:0] _GEN_3856 = 8'h3 < length_1 ? _GEN_3696 : _GEN_3536; // @[executor.scala 308:60]
  wire [7:0] _GEN_3857 = 8'h3 < length_1 ? _GEN_3697 : _GEN_3537; // @[executor.scala 308:60]
  wire [7:0] _GEN_3858 = 8'h3 < length_1 ? _GEN_3698 : _GEN_3538; // @[executor.scala 308:60]
  wire [7:0] _GEN_3859 = 8'h3 < length_1 ? _GEN_3699 : _GEN_3539; // @[executor.scala 308:60]
  wire [7:0] _GEN_3860 = 8'h3 < length_1 ? _GEN_3700 : _GEN_3540; // @[executor.scala 308:60]
  wire [7:0] _GEN_3861 = 8'h3 < length_1 ? _GEN_3701 : _GEN_3541; // @[executor.scala 308:60]
  wire [7:0] _GEN_3862 = 8'h3 < length_1 ? _GEN_3702 : _GEN_3542; // @[executor.scala 308:60]
  wire [7:0] _GEN_3863 = 8'h3 < length_1 ? _GEN_3703 : _GEN_3543; // @[executor.scala 308:60]
  wire [7:0] _GEN_3864 = 8'h3 < length_1 ? _GEN_3704 : _GEN_3544; // @[executor.scala 308:60]
  wire [7:0] _GEN_3865 = 8'h3 < length_1 ? _GEN_3705 : _GEN_3545; // @[executor.scala 308:60]
  wire [7:0] _GEN_3866 = 8'h3 < length_1 ? _GEN_3706 : _GEN_3546; // @[executor.scala 308:60]
  wire [7:0] _GEN_3867 = 8'h3 < length_1 ? _GEN_3707 : _GEN_3547; // @[executor.scala 308:60]
  wire [7:0] _GEN_3868 = 8'h3 < length_1 ? _GEN_3708 : _GEN_3548; // @[executor.scala 308:60]
  wire [7:0] _GEN_3869 = 8'h3 < length_1 ? _GEN_3709 : _GEN_3549; // @[executor.scala 308:60]
  wire [7:0] _GEN_3870 = 8'h3 < length_1 ? _GEN_3710 : _GEN_3550; // @[executor.scala 308:60]
  wire [7:0] _GEN_3871 = 8'h3 < length_1 ? _GEN_3711 : _GEN_3551; // @[executor.scala 308:60]
  wire [7:0] _GEN_3872 = 8'h3 < length_1 ? _GEN_3712 : _GEN_3552; // @[executor.scala 308:60]
  wire [7:0] _GEN_3873 = 8'h3 < length_1 ? _GEN_3713 : _GEN_3553; // @[executor.scala 308:60]
  wire [7:0] _GEN_3874 = 8'h3 < length_1 ? _GEN_3714 : _GEN_3554; // @[executor.scala 308:60]
  wire [7:0] _GEN_3875 = 8'h3 < length_1 ? _GEN_3715 : _GEN_3555; // @[executor.scala 308:60]
  wire [7:0] _GEN_3876 = 8'h3 < length_1 ? _GEN_3716 : _GEN_3556; // @[executor.scala 308:60]
  wire [7:0] _GEN_3877 = 8'h3 < length_1 ? _GEN_3717 : _GEN_3557; // @[executor.scala 308:60]
  wire [7:0] _GEN_3878 = 8'h3 < length_1 ? _GEN_3718 : _GEN_3558; // @[executor.scala 308:60]
  wire [7:0] _GEN_3879 = 8'h3 < length_1 ? _GEN_3719 : _GEN_3559; // @[executor.scala 308:60]
  wire [7:0] _GEN_3880 = 8'h3 < length_1 ? _GEN_3720 : _GEN_3560; // @[executor.scala 308:60]
  wire [7:0] _GEN_3881 = 8'h3 < length_1 ? _GEN_3721 : _GEN_3561; // @[executor.scala 308:60]
  wire [7:0] _GEN_3882 = 8'h3 < length_1 ? _GEN_3722 : _GEN_3562; // @[executor.scala 308:60]
  wire [7:0] _GEN_3883 = 8'h3 < length_1 ? _GEN_3723 : _GEN_3563; // @[executor.scala 308:60]
  wire [7:0] _GEN_3884 = 8'h3 < length_1 ? _GEN_3724 : _GEN_3564; // @[executor.scala 308:60]
  wire [7:0] _GEN_3885 = 8'h3 < length_1 ? _GEN_3725 : _GEN_3565; // @[executor.scala 308:60]
  wire [7:0] _GEN_3886 = 8'h3 < length_1 ? _GEN_3726 : _GEN_3566; // @[executor.scala 308:60]
  wire [7:0] _GEN_3887 = 8'h3 < length_1 ? _GEN_3727 : _GEN_3567; // @[executor.scala 308:60]
  wire [7:0] _GEN_3888 = 8'h3 < length_1 ? _GEN_3728 : _GEN_3568; // @[executor.scala 308:60]
  wire [7:0] _GEN_3889 = 8'h3 < length_1 ? _GEN_3729 : _GEN_3569; // @[executor.scala 308:60]
  wire [7:0] _GEN_3890 = 8'h3 < length_1 ? _GEN_3730 : _GEN_3570; // @[executor.scala 308:60]
  wire [7:0] _GEN_3891 = 8'h3 < length_1 ? _GEN_3731 : _GEN_3571; // @[executor.scala 308:60]
  wire [7:0] _GEN_3892 = 8'h3 < length_1 ? _GEN_3732 : _GEN_3572; // @[executor.scala 308:60]
  wire [7:0] _GEN_3893 = 8'h3 < length_1 ? _GEN_3733 : _GEN_3573; // @[executor.scala 308:60]
  wire [7:0] _GEN_3894 = 8'h3 < length_1 ? _GEN_3734 : _GEN_3574; // @[executor.scala 308:60]
  wire [7:0] _GEN_3895 = 8'h3 < length_1 ? _GEN_3735 : _GEN_3575; // @[executor.scala 308:60]
  wire [7:0] _GEN_3896 = 8'h3 < length_1 ? _GEN_3736 : _GEN_3576; // @[executor.scala 308:60]
  wire [7:0] _GEN_3897 = 8'h3 < length_1 ? _GEN_3737 : _GEN_3577; // @[executor.scala 308:60]
  wire [7:0] _GEN_3898 = 8'h3 < length_1 ? _GEN_3738 : _GEN_3578; // @[executor.scala 308:60]
  wire [7:0] _GEN_3899 = 8'h3 < length_1 ? _GEN_3739 : _GEN_3579; // @[executor.scala 308:60]
  wire [7:0] _GEN_3900 = 8'h3 < length_1 ? _GEN_3740 : _GEN_3580; // @[executor.scala 308:60]
  wire [7:0] _GEN_3901 = 8'h3 < length_1 ? _GEN_3741 : _GEN_3581; // @[executor.scala 308:60]
  wire [7:0] _GEN_3902 = 8'h3 < length_1 ? _GEN_3742 : _GEN_3582; // @[executor.scala 308:60]
  wire [7:0] _GEN_3903 = 8'h3 < length_1 ? _GEN_3743 : _GEN_3583; // @[executor.scala 308:60]
  wire [7:0] _GEN_3904 = 8'h3 < length_1 ? _GEN_3744 : _GEN_3584; // @[executor.scala 308:60]
  wire [7:0] _GEN_3905 = 8'h3 < length_1 ? _GEN_3745 : _GEN_3585; // @[executor.scala 308:60]
  wire [7:0] _GEN_3906 = 8'h3 < length_1 ? _GEN_3746 : _GEN_3586; // @[executor.scala 308:60]
  wire [7:0] _GEN_3907 = 8'h3 < length_1 ? _GEN_3747 : _GEN_3587; // @[executor.scala 308:60]
  wire [7:0] _GEN_3908 = 8'h3 < length_1 ? _GEN_3748 : _GEN_3588; // @[executor.scala 308:60]
  wire [7:0] _GEN_3909 = 8'h3 < length_1 ? _GEN_3749 : _GEN_3589; // @[executor.scala 308:60]
  wire [7:0] _GEN_3910 = 8'h3 < length_1 ? _GEN_3750 : _GEN_3590; // @[executor.scala 308:60]
  wire [7:0] _GEN_3911 = 8'h3 < length_1 ? _GEN_3751 : _GEN_3591; // @[executor.scala 308:60]
  wire [7:0] _GEN_3912 = 8'h3 < length_1 ? _GEN_3752 : _GEN_3592; // @[executor.scala 308:60]
  wire [7:0] _GEN_3913 = 8'h3 < length_1 ? _GEN_3753 : _GEN_3593; // @[executor.scala 308:60]
  wire [7:0] _GEN_3914 = 8'h3 < length_1 ? _GEN_3754 : _GEN_3594; // @[executor.scala 308:60]
  wire [7:0] _GEN_3915 = 8'h3 < length_1 ? _GEN_3755 : _GEN_3595; // @[executor.scala 308:60]
  wire [7:0] _GEN_3916 = 8'h3 < length_1 ? _GEN_3756 : _GEN_3596; // @[executor.scala 308:60]
  wire [7:0] _GEN_3917 = 8'h3 < length_1 ? _GEN_3757 : _GEN_3597; // @[executor.scala 308:60]
  wire [7:0] _GEN_3918 = 8'h3 < length_1 ? _GEN_3758 : _GEN_3598; // @[executor.scala 308:60]
  wire [7:0] _GEN_3919 = 8'h3 < length_1 ? _GEN_3759 : _GEN_3599; // @[executor.scala 308:60]
  wire [7:0] _GEN_3920 = 8'h3 < length_1 ? _GEN_3760 : _GEN_3600; // @[executor.scala 308:60]
  wire [7:0] _GEN_3921 = 8'h3 < length_1 ? _GEN_3761 : _GEN_3601; // @[executor.scala 308:60]
  wire [7:0] _GEN_3922 = 8'h3 < length_1 ? _GEN_3762 : _GEN_3602; // @[executor.scala 308:60]
  wire [7:0] _GEN_3923 = 8'h3 < length_1 ? _GEN_3763 : _GEN_3603; // @[executor.scala 308:60]
  wire [7:0] _GEN_3924 = 8'h3 < length_1 ? _GEN_3764 : _GEN_3604; // @[executor.scala 308:60]
  wire [7:0] _GEN_3925 = 8'h3 < length_1 ? _GEN_3765 : _GEN_3605; // @[executor.scala 308:60]
  wire [7:0] _GEN_3926 = 8'h3 < length_1 ? _GEN_3766 : _GEN_3606; // @[executor.scala 308:60]
  wire [7:0] _GEN_3927 = 8'h3 < length_1 ? _GEN_3767 : _GEN_3607; // @[executor.scala 308:60]
  wire [7:0] _GEN_3928 = 8'h3 < length_1 ? _GEN_3768 : _GEN_3608; // @[executor.scala 308:60]
  wire [7:0] _GEN_3929 = 8'h3 < length_1 ? _GEN_3769 : _GEN_3609; // @[executor.scala 308:60]
  wire [7:0] _GEN_3930 = 8'h3 < length_1 ? _GEN_3770 : _GEN_3610; // @[executor.scala 308:60]
  wire [7:0] _GEN_3931 = 8'h3 < length_1 ? _GEN_3771 : _GEN_3611; // @[executor.scala 308:60]
  wire [7:0] _GEN_3932 = 8'h3 < length_1 ? _GEN_3772 : _GEN_3612; // @[executor.scala 308:60]
  wire [7:0] _GEN_3933 = 8'h3 < length_1 ? _GEN_3773 : _GEN_3613; // @[executor.scala 308:60]
  wire [7:0] _GEN_3934 = 8'h3 < length_1 ? _GEN_3774 : _GEN_3614; // @[executor.scala 308:60]
  wire [7:0] _GEN_3935 = 8'h3 < length_1 ? _GEN_3775 : _GEN_3615; // @[executor.scala 308:60]
  wire [7:0] _GEN_3936 = 8'h3 < length_1 ? _GEN_3776 : _GEN_3616; // @[executor.scala 308:60]
  wire [7:0] _GEN_3937 = 8'h3 < length_1 ? _GEN_3777 : _GEN_3617; // @[executor.scala 308:60]
  wire [7:0] _GEN_3938 = 8'h3 < length_1 ? _GEN_3778 : _GEN_3618; // @[executor.scala 308:60]
  wire [7:0] _GEN_3939 = 8'h3 < length_1 ? _GEN_3779 : _GEN_3619; // @[executor.scala 308:60]
  wire [7:0] _GEN_3940 = 8'h3 < length_1 ? _GEN_3780 : _GEN_3620; // @[executor.scala 308:60]
  wire [7:0] _GEN_3941 = 8'h3 < length_1 ? _GEN_3781 : _GEN_3621; // @[executor.scala 308:60]
  wire [7:0] _GEN_3942 = 8'h3 < length_1 ? _GEN_3782 : _GEN_3622; // @[executor.scala 308:60]
  wire [7:0] _GEN_3943 = 8'h3 < length_1 ? _GEN_3783 : _GEN_3623; // @[executor.scala 308:60]
  wire [7:0] _GEN_3944 = 8'h3 < length_1 ? _GEN_3784 : _GEN_3624; // @[executor.scala 308:60]
  wire [7:0] _GEN_3945 = 8'h3 < length_1 ? _GEN_3785 : _GEN_3625; // @[executor.scala 308:60]
  wire [7:0] _GEN_3946 = 8'h3 < length_1 ? _GEN_3786 : _GEN_3626; // @[executor.scala 308:60]
  wire [7:0] _GEN_3947 = 8'h3 < length_1 ? _GEN_3787 : _GEN_3627; // @[executor.scala 308:60]
  wire [7:0] _GEN_3948 = 8'h3 < length_1 ? _GEN_3788 : _GEN_3628; // @[executor.scala 308:60]
  wire [7:0] _GEN_3949 = 8'h3 < length_1 ? _GEN_3789 : _GEN_3629; // @[executor.scala 308:60]
  wire [7:0] _GEN_3950 = 8'h3 < length_1 ? _GEN_3790 : _GEN_3630; // @[executor.scala 308:60]
  wire [7:0] _GEN_3951 = 8'h3 < length_1 ? _GEN_3791 : _GEN_3631; // @[executor.scala 308:60]
  wire [7:0] _GEN_3952 = 8'h3 < length_1 ? _GEN_3792 : _GEN_3632; // @[executor.scala 308:60]
  wire [7:0] _GEN_3953 = 8'h3 < length_1 ? _GEN_3793 : _GEN_3633; // @[executor.scala 308:60]
  wire [7:0] _GEN_3954 = 8'h3 < length_1 ? _GEN_3794 : _GEN_3634; // @[executor.scala 308:60]
  wire [7:0] _GEN_3955 = 8'h3 < length_1 ? _GEN_3795 : _GEN_3635; // @[executor.scala 308:60]
  wire [7:0] _GEN_3956 = 8'h3 < length_1 ? _GEN_3796 : _GEN_3636; // @[executor.scala 308:60]
  wire [7:0] _GEN_3957 = 8'h3 < length_1 ? _GEN_3797 : _GEN_3637; // @[executor.scala 308:60]
  wire [7:0] _GEN_3958 = 8'h3 < length_1 ? _GEN_3798 : _GEN_3638; // @[executor.scala 308:60]
  wire [7:0] _GEN_3959 = 8'h3 < length_1 ? _GEN_3799 : _GEN_3639; // @[executor.scala 308:60]
  wire [7:0] _GEN_3960 = 8'h3 < length_1 ? _GEN_3800 : _GEN_3640; // @[executor.scala 308:60]
  wire [7:0] _GEN_3961 = 8'h3 < length_1 ? _GEN_3801 : _GEN_3641; // @[executor.scala 308:60]
  wire [7:0] _GEN_3962 = 8'h3 < length_1 ? _GEN_3802 : _GEN_3642; // @[executor.scala 308:60]
  wire [7:0] _GEN_3963 = 8'h3 < length_1 ? _GEN_3803 : _GEN_3643; // @[executor.scala 308:60]
  wire [7:0] _GEN_3964 = 8'h3 < length_1 ? _GEN_3804 : _GEN_3644; // @[executor.scala 308:60]
  wire [7:0] _GEN_3965 = 8'h3 < length_1 ? _GEN_3805 : _GEN_3645; // @[executor.scala 308:60]
  wire [7:0] _GEN_3966 = 8'h3 < length_1 ? _GEN_3806 : _GEN_3646; // @[executor.scala 308:60]
  wire [7:0] _GEN_3967 = 8'h3 < length_1 ? _GEN_3807 : _GEN_3647; // @[executor.scala 308:60]
  wire [7:0] _GEN_3968 = 8'h3 < length_1 ? _GEN_3808 : _GEN_3648; // @[executor.scala 308:60]
  wire [7:0] _GEN_3969 = 8'h3 < length_1 ? _GEN_3809 : _GEN_3649; // @[executor.scala 308:60]
  wire [7:0] _GEN_3970 = 8'h3 < length_1 ? _GEN_3810 : _GEN_3650; // @[executor.scala 308:60]
  wire [7:0] _GEN_3971 = 8'h3 < length_1 ? _GEN_3811 : _GEN_3651; // @[executor.scala 308:60]
  wire [7:0] _GEN_3972 = 8'h3 < length_1 ? _GEN_3812 : _GEN_3652; // @[executor.scala 308:60]
  wire [7:0] _GEN_3973 = 8'h3 < length_1 ? _GEN_3813 : _GEN_3653; // @[executor.scala 308:60]
  wire [7:0] _GEN_3974 = 8'h3 < length_1 ? _GEN_3814 : _GEN_3654; // @[executor.scala 308:60]
  wire [7:0] _GEN_3975 = 8'h3 < length_1 ? _GEN_3815 : _GEN_3655; // @[executor.scala 308:60]
  wire [7:0] _GEN_3976 = 8'h3 < length_1 ? _GEN_3816 : _GEN_3656; // @[executor.scala 308:60]
  wire [7:0] _GEN_3977 = 8'h3 < length_1 ? _GEN_3817 : _GEN_3657; // @[executor.scala 308:60]
  wire [7:0] _GEN_3978 = 8'h3 < length_1 ? _GEN_3818 : _GEN_3658; // @[executor.scala 308:60]
  wire [7:0] _GEN_3979 = 8'h3 < length_1 ? _GEN_3819 : _GEN_3659; // @[executor.scala 308:60]
  wire [7:0] _GEN_3980 = 8'h3 < length_1 ? _GEN_3820 : _GEN_3660; // @[executor.scala 308:60]
  wire [7:0] _GEN_3981 = 8'h3 < length_1 ? _GEN_3821 : _GEN_3661; // @[executor.scala 308:60]
  wire [7:0] _GEN_3982 = 8'h3 < length_1 ? _GEN_3822 : _GEN_3662; // @[executor.scala 308:60]
  wire [7:0] _GEN_3983 = 8'h3 < length_1 ? _GEN_3823 : _GEN_3663; // @[executor.scala 308:60]
  wire [7:0] _GEN_3984 = 8'h3 < length_1 ? _GEN_3824 : _GEN_3664; // @[executor.scala 308:60]
  wire [7:0] _GEN_3985 = 8'h3 < length_1 ? _GEN_3825 : _GEN_3665; // @[executor.scala 308:60]
  wire [7:0] _GEN_3986 = 8'h3 < length_1 ? _GEN_3826 : _GEN_3666; // @[executor.scala 308:60]
  wire [7:0] _GEN_3987 = 8'h3 < length_1 ? _GEN_3827 : _GEN_3667; // @[executor.scala 308:60]
  wire [7:0] _GEN_3988 = 8'h3 < length_1 ? _GEN_3828 : _GEN_3668; // @[executor.scala 308:60]
  wire [7:0] _GEN_3989 = 8'h3 < length_1 ? _GEN_3829 : _GEN_3669; // @[executor.scala 308:60]
  wire [7:0] _GEN_3990 = 8'h3 < length_1 ? _GEN_3830 : _GEN_3670; // @[executor.scala 308:60]
  wire [7:0] _GEN_3991 = 8'h3 < length_1 ? _GEN_3831 : _GEN_3671; // @[executor.scala 308:60]
  wire [7:0] _GEN_3992 = 8'h3 < length_1 ? _GEN_3832 : _GEN_3672; // @[executor.scala 308:60]
  wire [7:0] _GEN_3993 = 8'h3 < length_1 ? _GEN_3833 : _GEN_3673; // @[executor.scala 308:60]
  wire [7:0] _GEN_3994 = 8'h3 < length_1 ? _GEN_3834 : _GEN_3674; // @[executor.scala 308:60]
  wire [7:0] _GEN_3995 = 8'h3 < length_1 ? _GEN_3835 : _GEN_3675; // @[executor.scala 308:60]
  wire [7:0] _GEN_3996 = 8'h3 < length_1 ? _GEN_3836 : _GEN_3676; // @[executor.scala 308:60]
  wire [7:0] _GEN_3997 = 8'h3 < length_1 ? _GEN_3837 : _GEN_3677; // @[executor.scala 308:60]
  wire [7:0] _GEN_3998 = 8'h3 < length_1 ? _GEN_3838 : _GEN_3678; // @[executor.scala 308:60]
  wire [7:0] _GEN_3999 = 8'h3 < length_1 ? _GEN_3839 : _GEN_3679; // @[executor.scala 308:60]
  wire [7:0] _GEN_4000 = 8'h3 < length_1 ? _GEN_3840 : _GEN_3680; // @[executor.scala 308:60]
  wire [7:0] _GEN_4001 = 8'h3 < length_1 ? _GEN_3841 : _GEN_3681; // @[executor.scala 308:60]
  wire [7:0] field_byte_12 = field_1[31:24]; // @[executor.scala 305:57]
  wire [7:0] total_offset_12 = offset_1 + 8'h4; // @[executor.scala 307:57]
  wire [7:0] _GEN_4002 = 8'h0 == total_offset_12 ? field_byte_12 : _GEN_3842; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4003 = 8'h1 == total_offset_12 ? field_byte_12 : _GEN_3843; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4004 = 8'h2 == total_offset_12 ? field_byte_12 : _GEN_3844; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4005 = 8'h3 == total_offset_12 ? field_byte_12 : _GEN_3845; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4006 = 8'h4 == total_offset_12 ? field_byte_12 : _GEN_3846; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4007 = 8'h5 == total_offset_12 ? field_byte_12 : _GEN_3847; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4008 = 8'h6 == total_offset_12 ? field_byte_12 : _GEN_3848; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4009 = 8'h7 == total_offset_12 ? field_byte_12 : _GEN_3849; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4010 = 8'h8 == total_offset_12 ? field_byte_12 : _GEN_3850; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4011 = 8'h9 == total_offset_12 ? field_byte_12 : _GEN_3851; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4012 = 8'ha == total_offset_12 ? field_byte_12 : _GEN_3852; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4013 = 8'hb == total_offset_12 ? field_byte_12 : _GEN_3853; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4014 = 8'hc == total_offset_12 ? field_byte_12 : _GEN_3854; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4015 = 8'hd == total_offset_12 ? field_byte_12 : _GEN_3855; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4016 = 8'he == total_offset_12 ? field_byte_12 : _GEN_3856; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4017 = 8'hf == total_offset_12 ? field_byte_12 : _GEN_3857; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4018 = 8'h10 == total_offset_12 ? field_byte_12 : _GEN_3858; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4019 = 8'h11 == total_offset_12 ? field_byte_12 : _GEN_3859; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4020 = 8'h12 == total_offset_12 ? field_byte_12 : _GEN_3860; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4021 = 8'h13 == total_offset_12 ? field_byte_12 : _GEN_3861; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4022 = 8'h14 == total_offset_12 ? field_byte_12 : _GEN_3862; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4023 = 8'h15 == total_offset_12 ? field_byte_12 : _GEN_3863; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4024 = 8'h16 == total_offset_12 ? field_byte_12 : _GEN_3864; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4025 = 8'h17 == total_offset_12 ? field_byte_12 : _GEN_3865; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4026 = 8'h18 == total_offset_12 ? field_byte_12 : _GEN_3866; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4027 = 8'h19 == total_offset_12 ? field_byte_12 : _GEN_3867; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4028 = 8'h1a == total_offset_12 ? field_byte_12 : _GEN_3868; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4029 = 8'h1b == total_offset_12 ? field_byte_12 : _GEN_3869; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4030 = 8'h1c == total_offset_12 ? field_byte_12 : _GEN_3870; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4031 = 8'h1d == total_offset_12 ? field_byte_12 : _GEN_3871; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4032 = 8'h1e == total_offset_12 ? field_byte_12 : _GEN_3872; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4033 = 8'h1f == total_offset_12 ? field_byte_12 : _GEN_3873; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4034 = 8'h20 == total_offset_12 ? field_byte_12 : _GEN_3874; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4035 = 8'h21 == total_offset_12 ? field_byte_12 : _GEN_3875; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4036 = 8'h22 == total_offset_12 ? field_byte_12 : _GEN_3876; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4037 = 8'h23 == total_offset_12 ? field_byte_12 : _GEN_3877; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4038 = 8'h24 == total_offset_12 ? field_byte_12 : _GEN_3878; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4039 = 8'h25 == total_offset_12 ? field_byte_12 : _GEN_3879; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4040 = 8'h26 == total_offset_12 ? field_byte_12 : _GEN_3880; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4041 = 8'h27 == total_offset_12 ? field_byte_12 : _GEN_3881; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4042 = 8'h28 == total_offset_12 ? field_byte_12 : _GEN_3882; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4043 = 8'h29 == total_offset_12 ? field_byte_12 : _GEN_3883; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4044 = 8'h2a == total_offset_12 ? field_byte_12 : _GEN_3884; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4045 = 8'h2b == total_offset_12 ? field_byte_12 : _GEN_3885; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4046 = 8'h2c == total_offset_12 ? field_byte_12 : _GEN_3886; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4047 = 8'h2d == total_offset_12 ? field_byte_12 : _GEN_3887; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4048 = 8'h2e == total_offset_12 ? field_byte_12 : _GEN_3888; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4049 = 8'h2f == total_offset_12 ? field_byte_12 : _GEN_3889; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4050 = 8'h30 == total_offset_12 ? field_byte_12 : _GEN_3890; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4051 = 8'h31 == total_offset_12 ? field_byte_12 : _GEN_3891; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4052 = 8'h32 == total_offset_12 ? field_byte_12 : _GEN_3892; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4053 = 8'h33 == total_offset_12 ? field_byte_12 : _GEN_3893; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4054 = 8'h34 == total_offset_12 ? field_byte_12 : _GEN_3894; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4055 = 8'h35 == total_offset_12 ? field_byte_12 : _GEN_3895; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4056 = 8'h36 == total_offset_12 ? field_byte_12 : _GEN_3896; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4057 = 8'h37 == total_offset_12 ? field_byte_12 : _GEN_3897; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4058 = 8'h38 == total_offset_12 ? field_byte_12 : _GEN_3898; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4059 = 8'h39 == total_offset_12 ? field_byte_12 : _GEN_3899; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4060 = 8'h3a == total_offset_12 ? field_byte_12 : _GEN_3900; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4061 = 8'h3b == total_offset_12 ? field_byte_12 : _GEN_3901; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4062 = 8'h3c == total_offset_12 ? field_byte_12 : _GEN_3902; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4063 = 8'h3d == total_offset_12 ? field_byte_12 : _GEN_3903; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4064 = 8'h3e == total_offset_12 ? field_byte_12 : _GEN_3904; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4065 = 8'h3f == total_offset_12 ? field_byte_12 : _GEN_3905; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4066 = 8'h40 == total_offset_12 ? field_byte_12 : _GEN_3906; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4067 = 8'h41 == total_offset_12 ? field_byte_12 : _GEN_3907; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4068 = 8'h42 == total_offset_12 ? field_byte_12 : _GEN_3908; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4069 = 8'h43 == total_offset_12 ? field_byte_12 : _GEN_3909; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4070 = 8'h44 == total_offset_12 ? field_byte_12 : _GEN_3910; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4071 = 8'h45 == total_offset_12 ? field_byte_12 : _GEN_3911; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4072 = 8'h46 == total_offset_12 ? field_byte_12 : _GEN_3912; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4073 = 8'h47 == total_offset_12 ? field_byte_12 : _GEN_3913; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4074 = 8'h48 == total_offset_12 ? field_byte_12 : _GEN_3914; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4075 = 8'h49 == total_offset_12 ? field_byte_12 : _GEN_3915; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4076 = 8'h4a == total_offset_12 ? field_byte_12 : _GEN_3916; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4077 = 8'h4b == total_offset_12 ? field_byte_12 : _GEN_3917; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4078 = 8'h4c == total_offset_12 ? field_byte_12 : _GEN_3918; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4079 = 8'h4d == total_offset_12 ? field_byte_12 : _GEN_3919; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4080 = 8'h4e == total_offset_12 ? field_byte_12 : _GEN_3920; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4081 = 8'h4f == total_offset_12 ? field_byte_12 : _GEN_3921; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4082 = 8'h50 == total_offset_12 ? field_byte_12 : _GEN_3922; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4083 = 8'h51 == total_offset_12 ? field_byte_12 : _GEN_3923; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4084 = 8'h52 == total_offset_12 ? field_byte_12 : _GEN_3924; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4085 = 8'h53 == total_offset_12 ? field_byte_12 : _GEN_3925; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4086 = 8'h54 == total_offset_12 ? field_byte_12 : _GEN_3926; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4087 = 8'h55 == total_offset_12 ? field_byte_12 : _GEN_3927; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4088 = 8'h56 == total_offset_12 ? field_byte_12 : _GEN_3928; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4089 = 8'h57 == total_offset_12 ? field_byte_12 : _GEN_3929; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4090 = 8'h58 == total_offset_12 ? field_byte_12 : _GEN_3930; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4091 = 8'h59 == total_offset_12 ? field_byte_12 : _GEN_3931; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4092 = 8'h5a == total_offset_12 ? field_byte_12 : _GEN_3932; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4093 = 8'h5b == total_offset_12 ? field_byte_12 : _GEN_3933; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4094 = 8'h5c == total_offset_12 ? field_byte_12 : _GEN_3934; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4095 = 8'h5d == total_offset_12 ? field_byte_12 : _GEN_3935; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4096 = 8'h5e == total_offset_12 ? field_byte_12 : _GEN_3936; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4097 = 8'h5f == total_offset_12 ? field_byte_12 : _GEN_3937; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4098 = 8'h60 == total_offset_12 ? field_byte_12 : _GEN_3938; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4099 = 8'h61 == total_offset_12 ? field_byte_12 : _GEN_3939; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4100 = 8'h62 == total_offset_12 ? field_byte_12 : _GEN_3940; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4101 = 8'h63 == total_offset_12 ? field_byte_12 : _GEN_3941; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4102 = 8'h64 == total_offset_12 ? field_byte_12 : _GEN_3942; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4103 = 8'h65 == total_offset_12 ? field_byte_12 : _GEN_3943; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4104 = 8'h66 == total_offset_12 ? field_byte_12 : _GEN_3944; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4105 = 8'h67 == total_offset_12 ? field_byte_12 : _GEN_3945; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4106 = 8'h68 == total_offset_12 ? field_byte_12 : _GEN_3946; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4107 = 8'h69 == total_offset_12 ? field_byte_12 : _GEN_3947; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4108 = 8'h6a == total_offset_12 ? field_byte_12 : _GEN_3948; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4109 = 8'h6b == total_offset_12 ? field_byte_12 : _GEN_3949; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4110 = 8'h6c == total_offset_12 ? field_byte_12 : _GEN_3950; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4111 = 8'h6d == total_offset_12 ? field_byte_12 : _GEN_3951; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4112 = 8'h6e == total_offset_12 ? field_byte_12 : _GEN_3952; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4113 = 8'h6f == total_offset_12 ? field_byte_12 : _GEN_3953; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4114 = 8'h70 == total_offset_12 ? field_byte_12 : _GEN_3954; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4115 = 8'h71 == total_offset_12 ? field_byte_12 : _GEN_3955; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4116 = 8'h72 == total_offset_12 ? field_byte_12 : _GEN_3956; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4117 = 8'h73 == total_offset_12 ? field_byte_12 : _GEN_3957; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4118 = 8'h74 == total_offset_12 ? field_byte_12 : _GEN_3958; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4119 = 8'h75 == total_offset_12 ? field_byte_12 : _GEN_3959; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4120 = 8'h76 == total_offset_12 ? field_byte_12 : _GEN_3960; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4121 = 8'h77 == total_offset_12 ? field_byte_12 : _GEN_3961; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4122 = 8'h78 == total_offset_12 ? field_byte_12 : _GEN_3962; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4123 = 8'h79 == total_offset_12 ? field_byte_12 : _GEN_3963; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4124 = 8'h7a == total_offset_12 ? field_byte_12 : _GEN_3964; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4125 = 8'h7b == total_offset_12 ? field_byte_12 : _GEN_3965; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4126 = 8'h7c == total_offset_12 ? field_byte_12 : _GEN_3966; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4127 = 8'h7d == total_offset_12 ? field_byte_12 : _GEN_3967; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4128 = 8'h7e == total_offset_12 ? field_byte_12 : _GEN_3968; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4129 = 8'h7f == total_offset_12 ? field_byte_12 : _GEN_3969; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4130 = 8'h80 == total_offset_12 ? field_byte_12 : _GEN_3970; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4131 = 8'h81 == total_offset_12 ? field_byte_12 : _GEN_3971; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4132 = 8'h82 == total_offset_12 ? field_byte_12 : _GEN_3972; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4133 = 8'h83 == total_offset_12 ? field_byte_12 : _GEN_3973; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4134 = 8'h84 == total_offset_12 ? field_byte_12 : _GEN_3974; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4135 = 8'h85 == total_offset_12 ? field_byte_12 : _GEN_3975; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4136 = 8'h86 == total_offset_12 ? field_byte_12 : _GEN_3976; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4137 = 8'h87 == total_offset_12 ? field_byte_12 : _GEN_3977; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4138 = 8'h88 == total_offset_12 ? field_byte_12 : _GEN_3978; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4139 = 8'h89 == total_offset_12 ? field_byte_12 : _GEN_3979; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4140 = 8'h8a == total_offset_12 ? field_byte_12 : _GEN_3980; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4141 = 8'h8b == total_offset_12 ? field_byte_12 : _GEN_3981; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4142 = 8'h8c == total_offset_12 ? field_byte_12 : _GEN_3982; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4143 = 8'h8d == total_offset_12 ? field_byte_12 : _GEN_3983; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4144 = 8'h8e == total_offset_12 ? field_byte_12 : _GEN_3984; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4145 = 8'h8f == total_offset_12 ? field_byte_12 : _GEN_3985; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4146 = 8'h90 == total_offset_12 ? field_byte_12 : _GEN_3986; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4147 = 8'h91 == total_offset_12 ? field_byte_12 : _GEN_3987; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4148 = 8'h92 == total_offset_12 ? field_byte_12 : _GEN_3988; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4149 = 8'h93 == total_offset_12 ? field_byte_12 : _GEN_3989; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4150 = 8'h94 == total_offset_12 ? field_byte_12 : _GEN_3990; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4151 = 8'h95 == total_offset_12 ? field_byte_12 : _GEN_3991; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4152 = 8'h96 == total_offset_12 ? field_byte_12 : _GEN_3992; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4153 = 8'h97 == total_offset_12 ? field_byte_12 : _GEN_3993; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4154 = 8'h98 == total_offset_12 ? field_byte_12 : _GEN_3994; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4155 = 8'h99 == total_offset_12 ? field_byte_12 : _GEN_3995; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4156 = 8'h9a == total_offset_12 ? field_byte_12 : _GEN_3996; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4157 = 8'h9b == total_offset_12 ? field_byte_12 : _GEN_3997; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4158 = 8'h9c == total_offset_12 ? field_byte_12 : _GEN_3998; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4159 = 8'h9d == total_offset_12 ? field_byte_12 : _GEN_3999; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4160 = 8'h9e == total_offset_12 ? field_byte_12 : _GEN_4000; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4161 = 8'h9f == total_offset_12 ? field_byte_12 : _GEN_4001; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4162 = 8'h4 < length_1 ? _GEN_4002 : _GEN_3842; // @[executor.scala 308:60]
  wire [7:0] _GEN_4163 = 8'h4 < length_1 ? _GEN_4003 : _GEN_3843; // @[executor.scala 308:60]
  wire [7:0] _GEN_4164 = 8'h4 < length_1 ? _GEN_4004 : _GEN_3844; // @[executor.scala 308:60]
  wire [7:0] _GEN_4165 = 8'h4 < length_1 ? _GEN_4005 : _GEN_3845; // @[executor.scala 308:60]
  wire [7:0] _GEN_4166 = 8'h4 < length_1 ? _GEN_4006 : _GEN_3846; // @[executor.scala 308:60]
  wire [7:0] _GEN_4167 = 8'h4 < length_1 ? _GEN_4007 : _GEN_3847; // @[executor.scala 308:60]
  wire [7:0] _GEN_4168 = 8'h4 < length_1 ? _GEN_4008 : _GEN_3848; // @[executor.scala 308:60]
  wire [7:0] _GEN_4169 = 8'h4 < length_1 ? _GEN_4009 : _GEN_3849; // @[executor.scala 308:60]
  wire [7:0] _GEN_4170 = 8'h4 < length_1 ? _GEN_4010 : _GEN_3850; // @[executor.scala 308:60]
  wire [7:0] _GEN_4171 = 8'h4 < length_1 ? _GEN_4011 : _GEN_3851; // @[executor.scala 308:60]
  wire [7:0] _GEN_4172 = 8'h4 < length_1 ? _GEN_4012 : _GEN_3852; // @[executor.scala 308:60]
  wire [7:0] _GEN_4173 = 8'h4 < length_1 ? _GEN_4013 : _GEN_3853; // @[executor.scala 308:60]
  wire [7:0] _GEN_4174 = 8'h4 < length_1 ? _GEN_4014 : _GEN_3854; // @[executor.scala 308:60]
  wire [7:0] _GEN_4175 = 8'h4 < length_1 ? _GEN_4015 : _GEN_3855; // @[executor.scala 308:60]
  wire [7:0] _GEN_4176 = 8'h4 < length_1 ? _GEN_4016 : _GEN_3856; // @[executor.scala 308:60]
  wire [7:0] _GEN_4177 = 8'h4 < length_1 ? _GEN_4017 : _GEN_3857; // @[executor.scala 308:60]
  wire [7:0] _GEN_4178 = 8'h4 < length_1 ? _GEN_4018 : _GEN_3858; // @[executor.scala 308:60]
  wire [7:0] _GEN_4179 = 8'h4 < length_1 ? _GEN_4019 : _GEN_3859; // @[executor.scala 308:60]
  wire [7:0] _GEN_4180 = 8'h4 < length_1 ? _GEN_4020 : _GEN_3860; // @[executor.scala 308:60]
  wire [7:0] _GEN_4181 = 8'h4 < length_1 ? _GEN_4021 : _GEN_3861; // @[executor.scala 308:60]
  wire [7:0] _GEN_4182 = 8'h4 < length_1 ? _GEN_4022 : _GEN_3862; // @[executor.scala 308:60]
  wire [7:0] _GEN_4183 = 8'h4 < length_1 ? _GEN_4023 : _GEN_3863; // @[executor.scala 308:60]
  wire [7:0] _GEN_4184 = 8'h4 < length_1 ? _GEN_4024 : _GEN_3864; // @[executor.scala 308:60]
  wire [7:0] _GEN_4185 = 8'h4 < length_1 ? _GEN_4025 : _GEN_3865; // @[executor.scala 308:60]
  wire [7:0] _GEN_4186 = 8'h4 < length_1 ? _GEN_4026 : _GEN_3866; // @[executor.scala 308:60]
  wire [7:0] _GEN_4187 = 8'h4 < length_1 ? _GEN_4027 : _GEN_3867; // @[executor.scala 308:60]
  wire [7:0] _GEN_4188 = 8'h4 < length_1 ? _GEN_4028 : _GEN_3868; // @[executor.scala 308:60]
  wire [7:0] _GEN_4189 = 8'h4 < length_1 ? _GEN_4029 : _GEN_3869; // @[executor.scala 308:60]
  wire [7:0] _GEN_4190 = 8'h4 < length_1 ? _GEN_4030 : _GEN_3870; // @[executor.scala 308:60]
  wire [7:0] _GEN_4191 = 8'h4 < length_1 ? _GEN_4031 : _GEN_3871; // @[executor.scala 308:60]
  wire [7:0] _GEN_4192 = 8'h4 < length_1 ? _GEN_4032 : _GEN_3872; // @[executor.scala 308:60]
  wire [7:0] _GEN_4193 = 8'h4 < length_1 ? _GEN_4033 : _GEN_3873; // @[executor.scala 308:60]
  wire [7:0] _GEN_4194 = 8'h4 < length_1 ? _GEN_4034 : _GEN_3874; // @[executor.scala 308:60]
  wire [7:0] _GEN_4195 = 8'h4 < length_1 ? _GEN_4035 : _GEN_3875; // @[executor.scala 308:60]
  wire [7:0] _GEN_4196 = 8'h4 < length_1 ? _GEN_4036 : _GEN_3876; // @[executor.scala 308:60]
  wire [7:0] _GEN_4197 = 8'h4 < length_1 ? _GEN_4037 : _GEN_3877; // @[executor.scala 308:60]
  wire [7:0] _GEN_4198 = 8'h4 < length_1 ? _GEN_4038 : _GEN_3878; // @[executor.scala 308:60]
  wire [7:0] _GEN_4199 = 8'h4 < length_1 ? _GEN_4039 : _GEN_3879; // @[executor.scala 308:60]
  wire [7:0] _GEN_4200 = 8'h4 < length_1 ? _GEN_4040 : _GEN_3880; // @[executor.scala 308:60]
  wire [7:0] _GEN_4201 = 8'h4 < length_1 ? _GEN_4041 : _GEN_3881; // @[executor.scala 308:60]
  wire [7:0] _GEN_4202 = 8'h4 < length_1 ? _GEN_4042 : _GEN_3882; // @[executor.scala 308:60]
  wire [7:0] _GEN_4203 = 8'h4 < length_1 ? _GEN_4043 : _GEN_3883; // @[executor.scala 308:60]
  wire [7:0] _GEN_4204 = 8'h4 < length_1 ? _GEN_4044 : _GEN_3884; // @[executor.scala 308:60]
  wire [7:0] _GEN_4205 = 8'h4 < length_1 ? _GEN_4045 : _GEN_3885; // @[executor.scala 308:60]
  wire [7:0] _GEN_4206 = 8'h4 < length_1 ? _GEN_4046 : _GEN_3886; // @[executor.scala 308:60]
  wire [7:0] _GEN_4207 = 8'h4 < length_1 ? _GEN_4047 : _GEN_3887; // @[executor.scala 308:60]
  wire [7:0] _GEN_4208 = 8'h4 < length_1 ? _GEN_4048 : _GEN_3888; // @[executor.scala 308:60]
  wire [7:0] _GEN_4209 = 8'h4 < length_1 ? _GEN_4049 : _GEN_3889; // @[executor.scala 308:60]
  wire [7:0] _GEN_4210 = 8'h4 < length_1 ? _GEN_4050 : _GEN_3890; // @[executor.scala 308:60]
  wire [7:0] _GEN_4211 = 8'h4 < length_1 ? _GEN_4051 : _GEN_3891; // @[executor.scala 308:60]
  wire [7:0] _GEN_4212 = 8'h4 < length_1 ? _GEN_4052 : _GEN_3892; // @[executor.scala 308:60]
  wire [7:0] _GEN_4213 = 8'h4 < length_1 ? _GEN_4053 : _GEN_3893; // @[executor.scala 308:60]
  wire [7:0] _GEN_4214 = 8'h4 < length_1 ? _GEN_4054 : _GEN_3894; // @[executor.scala 308:60]
  wire [7:0] _GEN_4215 = 8'h4 < length_1 ? _GEN_4055 : _GEN_3895; // @[executor.scala 308:60]
  wire [7:0] _GEN_4216 = 8'h4 < length_1 ? _GEN_4056 : _GEN_3896; // @[executor.scala 308:60]
  wire [7:0] _GEN_4217 = 8'h4 < length_1 ? _GEN_4057 : _GEN_3897; // @[executor.scala 308:60]
  wire [7:0] _GEN_4218 = 8'h4 < length_1 ? _GEN_4058 : _GEN_3898; // @[executor.scala 308:60]
  wire [7:0] _GEN_4219 = 8'h4 < length_1 ? _GEN_4059 : _GEN_3899; // @[executor.scala 308:60]
  wire [7:0] _GEN_4220 = 8'h4 < length_1 ? _GEN_4060 : _GEN_3900; // @[executor.scala 308:60]
  wire [7:0] _GEN_4221 = 8'h4 < length_1 ? _GEN_4061 : _GEN_3901; // @[executor.scala 308:60]
  wire [7:0] _GEN_4222 = 8'h4 < length_1 ? _GEN_4062 : _GEN_3902; // @[executor.scala 308:60]
  wire [7:0] _GEN_4223 = 8'h4 < length_1 ? _GEN_4063 : _GEN_3903; // @[executor.scala 308:60]
  wire [7:0] _GEN_4224 = 8'h4 < length_1 ? _GEN_4064 : _GEN_3904; // @[executor.scala 308:60]
  wire [7:0] _GEN_4225 = 8'h4 < length_1 ? _GEN_4065 : _GEN_3905; // @[executor.scala 308:60]
  wire [7:0] _GEN_4226 = 8'h4 < length_1 ? _GEN_4066 : _GEN_3906; // @[executor.scala 308:60]
  wire [7:0] _GEN_4227 = 8'h4 < length_1 ? _GEN_4067 : _GEN_3907; // @[executor.scala 308:60]
  wire [7:0] _GEN_4228 = 8'h4 < length_1 ? _GEN_4068 : _GEN_3908; // @[executor.scala 308:60]
  wire [7:0] _GEN_4229 = 8'h4 < length_1 ? _GEN_4069 : _GEN_3909; // @[executor.scala 308:60]
  wire [7:0] _GEN_4230 = 8'h4 < length_1 ? _GEN_4070 : _GEN_3910; // @[executor.scala 308:60]
  wire [7:0] _GEN_4231 = 8'h4 < length_1 ? _GEN_4071 : _GEN_3911; // @[executor.scala 308:60]
  wire [7:0] _GEN_4232 = 8'h4 < length_1 ? _GEN_4072 : _GEN_3912; // @[executor.scala 308:60]
  wire [7:0] _GEN_4233 = 8'h4 < length_1 ? _GEN_4073 : _GEN_3913; // @[executor.scala 308:60]
  wire [7:0] _GEN_4234 = 8'h4 < length_1 ? _GEN_4074 : _GEN_3914; // @[executor.scala 308:60]
  wire [7:0] _GEN_4235 = 8'h4 < length_1 ? _GEN_4075 : _GEN_3915; // @[executor.scala 308:60]
  wire [7:0] _GEN_4236 = 8'h4 < length_1 ? _GEN_4076 : _GEN_3916; // @[executor.scala 308:60]
  wire [7:0] _GEN_4237 = 8'h4 < length_1 ? _GEN_4077 : _GEN_3917; // @[executor.scala 308:60]
  wire [7:0] _GEN_4238 = 8'h4 < length_1 ? _GEN_4078 : _GEN_3918; // @[executor.scala 308:60]
  wire [7:0] _GEN_4239 = 8'h4 < length_1 ? _GEN_4079 : _GEN_3919; // @[executor.scala 308:60]
  wire [7:0] _GEN_4240 = 8'h4 < length_1 ? _GEN_4080 : _GEN_3920; // @[executor.scala 308:60]
  wire [7:0] _GEN_4241 = 8'h4 < length_1 ? _GEN_4081 : _GEN_3921; // @[executor.scala 308:60]
  wire [7:0] _GEN_4242 = 8'h4 < length_1 ? _GEN_4082 : _GEN_3922; // @[executor.scala 308:60]
  wire [7:0] _GEN_4243 = 8'h4 < length_1 ? _GEN_4083 : _GEN_3923; // @[executor.scala 308:60]
  wire [7:0] _GEN_4244 = 8'h4 < length_1 ? _GEN_4084 : _GEN_3924; // @[executor.scala 308:60]
  wire [7:0] _GEN_4245 = 8'h4 < length_1 ? _GEN_4085 : _GEN_3925; // @[executor.scala 308:60]
  wire [7:0] _GEN_4246 = 8'h4 < length_1 ? _GEN_4086 : _GEN_3926; // @[executor.scala 308:60]
  wire [7:0] _GEN_4247 = 8'h4 < length_1 ? _GEN_4087 : _GEN_3927; // @[executor.scala 308:60]
  wire [7:0] _GEN_4248 = 8'h4 < length_1 ? _GEN_4088 : _GEN_3928; // @[executor.scala 308:60]
  wire [7:0] _GEN_4249 = 8'h4 < length_1 ? _GEN_4089 : _GEN_3929; // @[executor.scala 308:60]
  wire [7:0] _GEN_4250 = 8'h4 < length_1 ? _GEN_4090 : _GEN_3930; // @[executor.scala 308:60]
  wire [7:0] _GEN_4251 = 8'h4 < length_1 ? _GEN_4091 : _GEN_3931; // @[executor.scala 308:60]
  wire [7:0] _GEN_4252 = 8'h4 < length_1 ? _GEN_4092 : _GEN_3932; // @[executor.scala 308:60]
  wire [7:0] _GEN_4253 = 8'h4 < length_1 ? _GEN_4093 : _GEN_3933; // @[executor.scala 308:60]
  wire [7:0] _GEN_4254 = 8'h4 < length_1 ? _GEN_4094 : _GEN_3934; // @[executor.scala 308:60]
  wire [7:0] _GEN_4255 = 8'h4 < length_1 ? _GEN_4095 : _GEN_3935; // @[executor.scala 308:60]
  wire [7:0] _GEN_4256 = 8'h4 < length_1 ? _GEN_4096 : _GEN_3936; // @[executor.scala 308:60]
  wire [7:0] _GEN_4257 = 8'h4 < length_1 ? _GEN_4097 : _GEN_3937; // @[executor.scala 308:60]
  wire [7:0] _GEN_4258 = 8'h4 < length_1 ? _GEN_4098 : _GEN_3938; // @[executor.scala 308:60]
  wire [7:0] _GEN_4259 = 8'h4 < length_1 ? _GEN_4099 : _GEN_3939; // @[executor.scala 308:60]
  wire [7:0] _GEN_4260 = 8'h4 < length_1 ? _GEN_4100 : _GEN_3940; // @[executor.scala 308:60]
  wire [7:0] _GEN_4261 = 8'h4 < length_1 ? _GEN_4101 : _GEN_3941; // @[executor.scala 308:60]
  wire [7:0] _GEN_4262 = 8'h4 < length_1 ? _GEN_4102 : _GEN_3942; // @[executor.scala 308:60]
  wire [7:0] _GEN_4263 = 8'h4 < length_1 ? _GEN_4103 : _GEN_3943; // @[executor.scala 308:60]
  wire [7:0] _GEN_4264 = 8'h4 < length_1 ? _GEN_4104 : _GEN_3944; // @[executor.scala 308:60]
  wire [7:0] _GEN_4265 = 8'h4 < length_1 ? _GEN_4105 : _GEN_3945; // @[executor.scala 308:60]
  wire [7:0] _GEN_4266 = 8'h4 < length_1 ? _GEN_4106 : _GEN_3946; // @[executor.scala 308:60]
  wire [7:0] _GEN_4267 = 8'h4 < length_1 ? _GEN_4107 : _GEN_3947; // @[executor.scala 308:60]
  wire [7:0] _GEN_4268 = 8'h4 < length_1 ? _GEN_4108 : _GEN_3948; // @[executor.scala 308:60]
  wire [7:0] _GEN_4269 = 8'h4 < length_1 ? _GEN_4109 : _GEN_3949; // @[executor.scala 308:60]
  wire [7:0] _GEN_4270 = 8'h4 < length_1 ? _GEN_4110 : _GEN_3950; // @[executor.scala 308:60]
  wire [7:0] _GEN_4271 = 8'h4 < length_1 ? _GEN_4111 : _GEN_3951; // @[executor.scala 308:60]
  wire [7:0] _GEN_4272 = 8'h4 < length_1 ? _GEN_4112 : _GEN_3952; // @[executor.scala 308:60]
  wire [7:0] _GEN_4273 = 8'h4 < length_1 ? _GEN_4113 : _GEN_3953; // @[executor.scala 308:60]
  wire [7:0] _GEN_4274 = 8'h4 < length_1 ? _GEN_4114 : _GEN_3954; // @[executor.scala 308:60]
  wire [7:0] _GEN_4275 = 8'h4 < length_1 ? _GEN_4115 : _GEN_3955; // @[executor.scala 308:60]
  wire [7:0] _GEN_4276 = 8'h4 < length_1 ? _GEN_4116 : _GEN_3956; // @[executor.scala 308:60]
  wire [7:0] _GEN_4277 = 8'h4 < length_1 ? _GEN_4117 : _GEN_3957; // @[executor.scala 308:60]
  wire [7:0] _GEN_4278 = 8'h4 < length_1 ? _GEN_4118 : _GEN_3958; // @[executor.scala 308:60]
  wire [7:0] _GEN_4279 = 8'h4 < length_1 ? _GEN_4119 : _GEN_3959; // @[executor.scala 308:60]
  wire [7:0] _GEN_4280 = 8'h4 < length_1 ? _GEN_4120 : _GEN_3960; // @[executor.scala 308:60]
  wire [7:0] _GEN_4281 = 8'h4 < length_1 ? _GEN_4121 : _GEN_3961; // @[executor.scala 308:60]
  wire [7:0] _GEN_4282 = 8'h4 < length_1 ? _GEN_4122 : _GEN_3962; // @[executor.scala 308:60]
  wire [7:0] _GEN_4283 = 8'h4 < length_1 ? _GEN_4123 : _GEN_3963; // @[executor.scala 308:60]
  wire [7:0] _GEN_4284 = 8'h4 < length_1 ? _GEN_4124 : _GEN_3964; // @[executor.scala 308:60]
  wire [7:0] _GEN_4285 = 8'h4 < length_1 ? _GEN_4125 : _GEN_3965; // @[executor.scala 308:60]
  wire [7:0] _GEN_4286 = 8'h4 < length_1 ? _GEN_4126 : _GEN_3966; // @[executor.scala 308:60]
  wire [7:0] _GEN_4287 = 8'h4 < length_1 ? _GEN_4127 : _GEN_3967; // @[executor.scala 308:60]
  wire [7:0] _GEN_4288 = 8'h4 < length_1 ? _GEN_4128 : _GEN_3968; // @[executor.scala 308:60]
  wire [7:0] _GEN_4289 = 8'h4 < length_1 ? _GEN_4129 : _GEN_3969; // @[executor.scala 308:60]
  wire [7:0] _GEN_4290 = 8'h4 < length_1 ? _GEN_4130 : _GEN_3970; // @[executor.scala 308:60]
  wire [7:0] _GEN_4291 = 8'h4 < length_1 ? _GEN_4131 : _GEN_3971; // @[executor.scala 308:60]
  wire [7:0] _GEN_4292 = 8'h4 < length_1 ? _GEN_4132 : _GEN_3972; // @[executor.scala 308:60]
  wire [7:0] _GEN_4293 = 8'h4 < length_1 ? _GEN_4133 : _GEN_3973; // @[executor.scala 308:60]
  wire [7:0] _GEN_4294 = 8'h4 < length_1 ? _GEN_4134 : _GEN_3974; // @[executor.scala 308:60]
  wire [7:0] _GEN_4295 = 8'h4 < length_1 ? _GEN_4135 : _GEN_3975; // @[executor.scala 308:60]
  wire [7:0] _GEN_4296 = 8'h4 < length_1 ? _GEN_4136 : _GEN_3976; // @[executor.scala 308:60]
  wire [7:0] _GEN_4297 = 8'h4 < length_1 ? _GEN_4137 : _GEN_3977; // @[executor.scala 308:60]
  wire [7:0] _GEN_4298 = 8'h4 < length_1 ? _GEN_4138 : _GEN_3978; // @[executor.scala 308:60]
  wire [7:0] _GEN_4299 = 8'h4 < length_1 ? _GEN_4139 : _GEN_3979; // @[executor.scala 308:60]
  wire [7:0] _GEN_4300 = 8'h4 < length_1 ? _GEN_4140 : _GEN_3980; // @[executor.scala 308:60]
  wire [7:0] _GEN_4301 = 8'h4 < length_1 ? _GEN_4141 : _GEN_3981; // @[executor.scala 308:60]
  wire [7:0] _GEN_4302 = 8'h4 < length_1 ? _GEN_4142 : _GEN_3982; // @[executor.scala 308:60]
  wire [7:0] _GEN_4303 = 8'h4 < length_1 ? _GEN_4143 : _GEN_3983; // @[executor.scala 308:60]
  wire [7:0] _GEN_4304 = 8'h4 < length_1 ? _GEN_4144 : _GEN_3984; // @[executor.scala 308:60]
  wire [7:0] _GEN_4305 = 8'h4 < length_1 ? _GEN_4145 : _GEN_3985; // @[executor.scala 308:60]
  wire [7:0] _GEN_4306 = 8'h4 < length_1 ? _GEN_4146 : _GEN_3986; // @[executor.scala 308:60]
  wire [7:0] _GEN_4307 = 8'h4 < length_1 ? _GEN_4147 : _GEN_3987; // @[executor.scala 308:60]
  wire [7:0] _GEN_4308 = 8'h4 < length_1 ? _GEN_4148 : _GEN_3988; // @[executor.scala 308:60]
  wire [7:0] _GEN_4309 = 8'h4 < length_1 ? _GEN_4149 : _GEN_3989; // @[executor.scala 308:60]
  wire [7:0] _GEN_4310 = 8'h4 < length_1 ? _GEN_4150 : _GEN_3990; // @[executor.scala 308:60]
  wire [7:0] _GEN_4311 = 8'h4 < length_1 ? _GEN_4151 : _GEN_3991; // @[executor.scala 308:60]
  wire [7:0] _GEN_4312 = 8'h4 < length_1 ? _GEN_4152 : _GEN_3992; // @[executor.scala 308:60]
  wire [7:0] _GEN_4313 = 8'h4 < length_1 ? _GEN_4153 : _GEN_3993; // @[executor.scala 308:60]
  wire [7:0] _GEN_4314 = 8'h4 < length_1 ? _GEN_4154 : _GEN_3994; // @[executor.scala 308:60]
  wire [7:0] _GEN_4315 = 8'h4 < length_1 ? _GEN_4155 : _GEN_3995; // @[executor.scala 308:60]
  wire [7:0] _GEN_4316 = 8'h4 < length_1 ? _GEN_4156 : _GEN_3996; // @[executor.scala 308:60]
  wire [7:0] _GEN_4317 = 8'h4 < length_1 ? _GEN_4157 : _GEN_3997; // @[executor.scala 308:60]
  wire [7:0] _GEN_4318 = 8'h4 < length_1 ? _GEN_4158 : _GEN_3998; // @[executor.scala 308:60]
  wire [7:0] _GEN_4319 = 8'h4 < length_1 ? _GEN_4159 : _GEN_3999; // @[executor.scala 308:60]
  wire [7:0] _GEN_4320 = 8'h4 < length_1 ? _GEN_4160 : _GEN_4000; // @[executor.scala 308:60]
  wire [7:0] _GEN_4321 = 8'h4 < length_1 ? _GEN_4161 : _GEN_4001; // @[executor.scala 308:60]
  wire [7:0] field_byte_13 = field_1[23:16]; // @[executor.scala 305:57]
  wire [7:0] total_offset_13 = offset_1 + 8'h5; // @[executor.scala 307:57]
  wire [7:0] _GEN_4322 = 8'h0 == total_offset_13 ? field_byte_13 : _GEN_4162; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4323 = 8'h1 == total_offset_13 ? field_byte_13 : _GEN_4163; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4324 = 8'h2 == total_offset_13 ? field_byte_13 : _GEN_4164; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4325 = 8'h3 == total_offset_13 ? field_byte_13 : _GEN_4165; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4326 = 8'h4 == total_offset_13 ? field_byte_13 : _GEN_4166; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4327 = 8'h5 == total_offset_13 ? field_byte_13 : _GEN_4167; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4328 = 8'h6 == total_offset_13 ? field_byte_13 : _GEN_4168; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4329 = 8'h7 == total_offset_13 ? field_byte_13 : _GEN_4169; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4330 = 8'h8 == total_offset_13 ? field_byte_13 : _GEN_4170; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4331 = 8'h9 == total_offset_13 ? field_byte_13 : _GEN_4171; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4332 = 8'ha == total_offset_13 ? field_byte_13 : _GEN_4172; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4333 = 8'hb == total_offset_13 ? field_byte_13 : _GEN_4173; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4334 = 8'hc == total_offset_13 ? field_byte_13 : _GEN_4174; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4335 = 8'hd == total_offset_13 ? field_byte_13 : _GEN_4175; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4336 = 8'he == total_offset_13 ? field_byte_13 : _GEN_4176; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4337 = 8'hf == total_offset_13 ? field_byte_13 : _GEN_4177; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4338 = 8'h10 == total_offset_13 ? field_byte_13 : _GEN_4178; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4339 = 8'h11 == total_offset_13 ? field_byte_13 : _GEN_4179; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4340 = 8'h12 == total_offset_13 ? field_byte_13 : _GEN_4180; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4341 = 8'h13 == total_offset_13 ? field_byte_13 : _GEN_4181; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4342 = 8'h14 == total_offset_13 ? field_byte_13 : _GEN_4182; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4343 = 8'h15 == total_offset_13 ? field_byte_13 : _GEN_4183; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4344 = 8'h16 == total_offset_13 ? field_byte_13 : _GEN_4184; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4345 = 8'h17 == total_offset_13 ? field_byte_13 : _GEN_4185; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4346 = 8'h18 == total_offset_13 ? field_byte_13 : _GEN_4186; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4347 = 8'h19 == total_offset_13 ? field_byte_13 : _GEN_4187; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4348 = 8'h1a == total_offset_13 ? field_byte_13 : _GEN_4188; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4349 = 8'h1b == total_offset_13 ? field_byte_13 : _GEN_4189; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4350 = 8'h1c == total_offset_13 ? field_byte_13 : _GEN_4190; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4351 = 8'h1d == total_offset_13 ? field_byte_13 : _GEN_4191; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4352 = 8'h1e == total_offset_13 ? field_byte_13 : _GEN_4192; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4353 = 8'h1f == total_offset_13 ? field_byte_13 : _GEN_4193; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4354 = 8'h20 == total_offset_13 ? field_byte_13 : _GEN_4194; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4355 = 8'h21 == total_offset_13 ? field_byte_13 : _GEN_4195; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4356 = 8'h22 == total_offset_13 ? field_byte_13 : _GEN_4196; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4357 = 8'h23 == total_offset_13 ? field_byte_13 : _GEN_4197; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4358 = 8'h24 == total_offset_13 ? field_byte_13 : _GEN_4198; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4359 = 8'h25 == total_offset_13 ? field_byte_13 : _GEN_4199; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4360 = 8'h26 == total_offset_13 ? field_byte_13 : _GEN_4200; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4361 = 8'h27 == total_offset_13 ? field_byte_13 : _GEN_4201; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4362 = 8'h28 == total_offset_13 ? field_byte_13 : _GEN_4202; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4363 = 8'h29 == total_offset_13 ? field_byte_13 : _GEN_4203; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4364 = 8'h2a == total_offset_13 ? field_byte_13 : _GEN_4204; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4365 = 8'h2b == total_offset_13 ? field_byte_13 : _GEN_4205; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4366 = 8'h2c == total_offset_13 ? field_byte_13 : _GEN_4206; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4367 = 8'h2d == total_offset_13 ? field_byte_13 : _GEN_4207; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4368 = 8'h2e == total_offset_13 ? field_byte_13 : _GEN_4208; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4369 = 8'h2f == total_offset_13 ? field_byte_13 : _GEN_4209; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4370 = 8'h30 == total_offset_13 ? field_byte_13 : _GEN_4210; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4371 = 8'h31 == total_offset_13 ? field_byte_13 : _GEN_4211; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4372 = 8'h32 == total_offset_13 ? field_byte_13 : _GEN_4212; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4373 = 8'h33 == total_offset_13 ? field_byte_13 : _GEN_4213; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4374 = 8'h34 == total_offset_13 ? field_byte_13 : _GEN_4214; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4375 = 8'h35 == total_offset_13 ? field_byte_13 : _GEN_4215; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4376 = 8'h36 == total_offset_13 ? field_byte_13 : _GEN_4216; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4377 = 8'h37 == total_offset_13 ? field_byte_13 : _GEN_4217; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4378 = 8'h38 == total_offset_13 ? field_byte_13 : _GEN_4218; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4379 = 8'h39 == total_offset_13 ? field_byte_13 : _GEN_4219; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4380 = 8'h3a == total_offset_13 ? field_byte_13 : _GEN_4220; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4381 = 8'h3b == total_offset_13 ? field_byte_13 : _GEN_4221; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4382 = 8'h3c == total_offset_13 ? field_byte_13 : _GEN_4222; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4383 = 8'h3d == total_offset_13 ? field_byte_13 : _GEN_4223; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4384 = 8'h3e == total_offset_13 ? field_byte_13 : _GEN_4224; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4385 = 8'h3f == total_offset_13 ? field_byte_13 : _GEN_4225; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4386 = 8'h40 == total_offset_13 ? field_byte_13 : _GEN_4226; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4387 = 8'h41 == total_offset_13 ? field_byte_13 : _GEN_4227; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4388 = 8'h42 == total_offset_13 ? field_byte_13 : _GEN_4228; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4389 = 8'h43 == total_offset_13 ? field_byte_13 : _GEN_4229; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4390 = 8'h44 == total_offset_13 ? field_byte_13 : _GEN_4230; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4391 = 8'h45 == total_offset_13 ? field_byte_13 : _GEN_4231; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4392 = 8'h46 == total_offset_13 ? field_byte_13 : _GEN_4232; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4393 = 8'h47 == total_offset_13 ? field_byte_13 : _GEN_4233; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4394 = 8'h48 == total_offset_13 ? field_byte_13 : _GEN_4234; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4395 = 8'h49 == total_offset_13 ? field_byte_13 : _GEN_4235; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4396 = 8'h4a == total_offset_13 ? field_byte_13 : _GEN_4236; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4397 = 8'h4b == total_offset_13 ? field_byte_13 : _GEN_4237; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4398 = 8'h4c == total_offset_13 ? field_byte_13 : _GEN_4238; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4399 = 8'h4d == total_offset_13 ? field_byte_13 : _GEN_4239; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4400 = 8'h4e == total_offset_13 ? field_byte_13 : _GEN_4240; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4401 = 8'h4f == total_offset_13 ? field_byte_13 : _GEN_4241; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4402 = 8'h50 == total_offset_13 ? field_byte_13 : _GEN_4242; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4403 = 8'h51 == total_offset_13 ? field_byte_13 : _GEN_4243; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4404 = 8'h52 == total_offset_13 ? field_byte_13 : _GEN_4244; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4405 = 8'h53 == total_offset_13 ? field_byte_13 : _GEN_4245; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4406 = 8'h54 == total_offset_13 ? field_byte_13 : _GEN_4246; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4407 = 8'h55 == total_offset_13 ? field_byte_13 : _GEN_4247; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4408 = 8'h56 == total_offset_13 ? field_byte_13 : _GEN_4248; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4409 = 8'h57 == total_offset_13 ? field_byte_13 : _GEN_4249; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4410 = 8'h58 == total_offset_13 ? field_byte_13 : _GEN_4250; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4411 = 8'h59 == total_offset_13 ? field_byte_13 : _GEN_4251; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4412 = 8'h5a == total_offset_13 ? field_byte_13 : _GEN_4252; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4413 = 8'h5b == total_offset_13 ? field_byte_13 : _GEN_4253; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4414 = 8'h5c == total_offset_13 ? field_byte_13 : _GEN_4254; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4415 = 8'h5d == total_offset_13 ? field_byte_13 : _GEN_4255; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4416 = 8'h5e == total_offset_13 ? field_byte_13 : _GEN_4256; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4417 = 8'h5f == total_offset_13 ? field_byte_13 : _GEN_4257; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4418 = 8'h60 == total_offset_13 ? field_byte_13 : _GEN_4258; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4419 = 8'h61 == total_offset_13 ? field_byte_13 : _GEN_4259; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4420 = 8'h62 == total_offset_13 ? field_byte_13 : _GEN_4260; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4421 = 8'h63 == total_offset_13 ? field_byte_13 : _GEN_4261; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4422 = 8'h64 == total_offset_13 ? field_byte_13 : _GEN_4262; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4423 = 8'h65 == total_offset_13 ? field_byte_13 : _GEN_4263; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4424 = 8'h66 == total_offset_13 ? field_byte_13 : _GEN_4264; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4425 = 8'h67 == total_offset_13 ? field_byte_13 : _GEN_4265; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4426 = 8'h68 == total_offset_13 ? field_byte_13 : _GEN_4266; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4427 = 8'h69 == total_offset_13 ? field_byte_13 : _GEN_4267; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4428 = 8'h6a == total_offset_13 ? field_byte_13 : _GEN_4268; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4429 = 8'h6b == total_offset_13 ? field_byte_13 : _GEN_4269; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4430 = 8'h6c == total_offset_13 ? field_byte_13 : _GEN_4270; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4431 = 8'h6d == total_offset_13 ? field_byte_13 : _GEN_4271; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4432 = 8'h6e == total_offset_13 ? field_byte_13 : _GEN_4272; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4433 = 8'h6f == total_offset_13 ? field_byte_13 : _GEN_4273; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4434 = 8'h70 == total_offset_13 ? field_byte_13 : _GEN_4274; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4435 = 8'h71 == total_offset_13 ? field_byte_13 : _GEN_4275; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4436 = 8'h72 == total_offset_13 ? field_byte_13 : _GEN_4276; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4437 = 8'h73 == total_offset_13 ? field_byte_13 : _GEN_4277; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4438 = 8'h74 == total_offset_13 ? field_byte_13 : _GEN_4278; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4439 = 8'h75 == total_offset_13 ? field_byte_13 : _GEN_4279; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4440 = 8'h76 == total_offset_13 ? field_byte_13 : _GEN_4280; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4441 = 8'h77 == total_offset_13 ? field_byte_13 : _GEN_4281; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4442 = 8'h78 == total_offset_13 ? field_byte_13 : _GEN_4282; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4443 = 8'h79 == total_offset_13 ? field_byte_13 : _GEN_4283; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4444 = 8'h7a == total_offset_13 ? field_byte_13 : _GEN_4284; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4445 = 8'h7b == total_offset_13 ? field_byte_13 : _GEN_4285; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4446 = 8'h7c == total_offset_13 ? field_byte_13 : _GEN_4286; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4447 = 8'h7d == total_offset_13 ? field_byte_13 : _GEN_4287; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4448 = 8'h7e == total_offset_13 ? field_byte_13 : _GEN_4288; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4449 = 8'h7f == total_offset_13 ? field_byte_13 : _GEN_4289; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4450 = 8'h80 == total_offset_13 ? field_byte_13 : _GEN_4290; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4451 = 8'h81 == total_offset_13 ? field_byte_13 : _GEN_4291; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4452 = 8'h82 == total_offset_13 ? field_byte_13 : _GEN_4292; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4453 = 8'h83 == total_offset_13 ? field_byte_13 : _GEN_4293; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4454 = 8'h84 == total_offset_13 ? field_byte_13 : _GEN_4294; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4455 = 8'h85 == total_offset_13 ? field_byte_13 : _GEN_4295; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4456 = 8'h86 == total_offset_13 ? field_byte_13 : _GEN_4296; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4457 = 8'h87 == total_offset_13 ? field_byte_13 : _GEN_4297; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4458 = 8'h88 == total_offset_13 ? field_byte_13 : _GEN_4298; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4459 = 8'h89 == total_offset_13 ? field_byte_13 : _GEN_4299; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4460 = 8'h8a == total_offset_13 ? field_byte_13 : _GEN_4300; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4461 = 8'h8b == total_offset_13 ? field_byte_13 : _GEN_4301; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4462 = 8'h8c == total_offset_13 ? field_byte_13 : _GEN_4302; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4463 = 8'h8d == total_offset_13 ? field_byte_13 : _GEN_4303; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4464 = 8'h8e == total_offset_13 ? field_byte_13 : _GEN_4304; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4465 = 8'h8f == total_offset_13 ? field_byte_13 : _GEN_4305; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4466 = 8'h90 == total_offset_13 ? field_byte_13 : _GEN_4306; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4467 = 8'h91 == total_offset_13 ? field_byte_13 : _GEN_4307; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4468 = 8'h92 == total_offset_13 ? field_byte_13 : _GEN_4308; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4469 = 8'h93 == total_offset_13 ? field_byte_13 : _GEN_4309; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4470 = 8'h94 == total_offset_13 ? field_byte_13 : _GEN_4310; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4471 = 8'h95 == total_offset_13 ? field_byte_13 : _GEN_4311; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4472 = 8'h96 == total_offset_13 ? field_byte_13 : _GEN_4312; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4473 = 8'h97 == total_offset_13 ? field_byte_13 : _GEN_4313; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4474 = 8'h98 == total_offset_13 ? field_byte_13 : _GEN_4314; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4475 = 8'h99 == total_offset_13 ? field_byte_13 : _GEN_4315; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4476 = 8'h9a == total_offset_13 ? field_byte_13 : _GEN_4316; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4477 = 8'h9b == total_offset_13 ? field_byte_13 : _GEN_4317; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4478 = 8'h9c == total_offset_13 ? field_byte_13 : _GEN_4318; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4479 = 8'h9d == total_offset_13 ? field_byte_13 : _GEN_4319; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4480 = 8'h9e == total_offset_13 ? field_byte_13 : _GEN_4320; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4481 = 8'h9f == total_offset_13 ? field_byte_13 : _GEN_4321; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4482 = 8'h5 < length_1 ? _GEN_4322 : _GEN_4162; // @[executor.scala 308:60]
  wire [7:0] _GEN_4483 = 8'h5 < length_1 ? _GEN_4323 : _GEN_4163; // @[executor.scala 308:60]
  wire [7:0] _GEN_4484 = 8'h5 < length_1 ? _GEN_4324 : _GEN_4164; // @[executor.scala 308:60]
  wire [7:0] _GEN_4485 = 8'h5 < length_1 ? _GEN_4325 : _GEN_4165; // @[executor.scala 308:60]
  wire [7:0] _GEN_4486 = 8'h5 < length_1 ? _GEN_4326 : _GEN_4166; // @[executor.scala 308:60]
  wire [7:0] _GEN_4487 = 8'h5 < length_1 ? _GEN_4327 : _GEN_4167; // @[executor.scala 308:60]
  wire [7:0] _GEN_4488 = 8'h5 < length_1 ? _GEN_4328 : _GEN_4168; // @[executor.scala 308:60]
  wire [7:0] _GEN_4489 = 8'h5 < length_1 ? _GEN_4329 : _GEN_4169; // @[executor.scala 308:60]
  wire [7:0] _GEN_4490 = 8'h5 < length_1 ? _GEN_4330 : _GEN_4170; // @[executor.scala 308:60]
  wire [7:0] _GEN_4491 = 8'h5 < length_1 ? _GEN_4331 : _GEN_4171; // @[executor.scala 308:60]
  wire [7:0] _GEN_4492 = 8'h5 < length_1 ? _GEN_4332 : _GEN_4172; // @[executor.scala 308:60]
  wire [7:0] _GEN_4493 = 8'h5 < length_1 ? _GEN_4333 : _GEN_4173; // @[executor.scala 308:60]
  wire [7:0] _GEN_4494 = 8'h5 < length_1 ? _GEN_4334 : _GEN_4174; // @[executor.scala 308:60]
  wire [7:0] _GEN_4495 = 8'h5 < length_1 ? _GEN_4335 : _GEN_4175; // @[executor.scala 308:60]
  wire [7:0] _GEN_4496 = 8'h5 < length_1 ? _GEN_4336 : _GEN_4176; // @[executor.scala 308:60]
  wire [7:0] _GEN_4497 = 8'h5 < length_1 ? _GEN_4337 : _GEN_4177; // @[executor.scala 308:60]
  wire [7:0] _GEN_4498 = 8'h5 < length_1 ? _GEN_4338 : _GEN_4178; // @[executor.scala 308:60]
  wire [7:0] _GEN_4499 = 8'h5 < length_1 ? _GEN_4339 : _GEN_4179; // @[executor.scala 308:60]
  wire [7:0] _GEN_4500 = 8'h5 < length_1 ? _GEN_4340 : _GEN_4180; // @[executor.scala 308:60]
  wire [7:0] _GEN_4501 = 8'h5 < length_1 ? _GEN_4341 : _GEN_4181; // @[executor.scala 308:60]
  wire [7:0] _GEN_4502 = 8'h5 < length_1 ? _GEN_4342 : _GEN_4182; // @[executor.scala 308:60]
  wire [7:0] _GEN_4503 = 8'h5 < length_1 ? _GEN_4343 : _GEN_4183; // @[executor.scala 308:60]
  wire [7:0] _GEN_4504 = 8'h5 < length_1 ? _GEN_4344 : _GEN_4184; // @[executor.scala 308:60]
  wire [7:0] _GEN_4505 = 8'h5 < length_1 ? _GEN_4345 : _GEN_4185; // @[executor.scala 308:60]
  wire [7:0] _GEN_4506 = 8'h5 < length_1 ? _GEN_4346 : _GEN_4186; // @[executor.scala 308:60]
  wire [7:0] _GEN_4507 = 8'h5 < length_1 ? _GEN_4347 : _GEN_4187; // @[executor.scala 308:60]
  wire [7:0] _GEN_4508 = 8'h5 < length_1 ? _GEN_4348 : _GEN_4188; // @[executor.scala 308:60]
  wire [7:0] _GEN_4509 = 8'h5 < length_1 ? _GEN_4349 : _GEN_4189; // @[executor.scala 308:60]
  wire [7:0] _GEN_4510 = 8'h5 < length_1 ? _GEN_4350 : _GEN_4190; // @[executor.scala 308:60]
  wire [7:0] _GEN_4511 = 8'h5 < length_1 ? _GEN_4351 : _GEN_4191; // @[executor.scala 308:60]
  wire [7:0] _GEN_4512 = 8'h5 < length_1 ? _GEN_4352 : _GEN_4192; // @[executor.scala 308:60]
  wire [7:0] _GEN_4513 = 8'h5 < length_1 ? _GEN_4353 : _GEN_4193; // @[executor.scala 308:60]
  wire [7:0] _GEN_4514 = 8'h5 < length_1 ? _GEN_4354 : _GEN_4194; // @[executor.scala 308:60]
  wire [7:0] _GEN_4515 = 8'h5 < length_1 ? _GEN_4355 : _GEN_4195; // @[executor.scala 308:60]
  wire [7:0] _GEN_4516 = 8'h5 < length_1 ? _GEN_4356 : _GEN_4196; // @[executor.scala 308:60]
  wire [7:0] _GEN_4517 = 8'h5 < length_1 ? _GEN_4357 : _GEN_4197; // @[executor.scala 308:60]
  wire [7:0] _GEN_4518 = 8'h5 < length_1 ? _GEN_4358 : _GEN_4198; // @[executor.scala 308:60]
  wire [7:0] _GEN_4519 = 8'h5 < length_1 ? _GEN_4359 : _GEN_4199; // @[executor.scala 308:60]
  wire [7:0] _GEN_4520 = 8'h5 < length_1 ? _GEN_4360 : _GEN_4200; // @[executor.scala 308:60]
  wire [7:0] _GEN_4521 = 8'h5 < length_1 ? _GEN_4361 : _GEN_4201; // @[executor.scala 308:60]
  wire [7:0] _GEN_4522 = 8'h5 < length_1 ? _GEN_4362 : _GEN_4202; // @[executor.scala 308:60]
  wire [7:0] _GEN_4523 = 8'h5 < length_1 ? _GEN_4363 : _GEN_4203; // @[executor.scala 308:60]
  wire [7:0] _GEN_4524 = 8'h5 < length_1 ? _GEN_4364 : _GEN_4204; // @[executor.scala 308:60]
  wire [7:0] _GEN_4525 = 8'h5 < length_1 ? _GEN_4365 : _GEN_4205; // @[executor.scala 308:60]
  wire [7:0] _GEN_4526 = 8'h5 < length_1 ? _GEN_4366 : _GEN_4206; // @[executor.scala 308:60]
  wire [7:0] _GEN_4527 = 8'h5 < length_1 ? _GEN_4367 : _GEN_4207; // @[executor.scala 308:60]
  wire [7:0] _GEN_4528 = 8'h5 < length_1 ? _GEN_4368 : _GEN_4208; // @[executor.scala 308:60]
  wire [7:0] _GEN_4529 = 8'h5 < length_1 ? _GEN_4369 : _GEN_4209; // @[executor.scala 308:60]
  wire [7:0] _GEN_4530 = 8'h5 < length_1 ? _GEN_4370 : _GEN_4210; // @[executor.scala 308:60]
  wire [7:0] _GEN_4531 = 8'h5 < length_1 ? _GEN_4371 : _GEN_4211; // @[executor.scala 308:60]
  wire [7:0] _GEN_4532 = 8'h5 < length_1 ? _GEN_4372 : _GEN_4212; // @[executor.scala 308:60]
  wire [7:0] _GEN_4533 = 8'h5 < length_1 ? _GEN_4373 : _GEN_4213; // @[executor.scala 308:60]
  wire [7:0] _GEN_4534 = 8'h5 < length_1 ? _GEN_4374 : _GEN_4214; // @[executor.scala 308:60]
  wire [7:0] _GEN_4535 = 8'h5 < length_1 ? _GEN_4375 : _GEN_4215; // @[executor.scala 308:60]
  wire [7:0] _GEN_4536 = 8'h5 < length_1 ? _GEN_4376 : _GEN_4216; // @[executor.scala 308:60]
  wire [7:0] _GEN_4537 = 8'h5 < length_1 ? _GEN_4377 : _GEN_4217; // @[executor.scala 308:60]
  wire [7:0] _GEN_4538 = 8'h5 < length_1 ? _GEN_4378 : _GEN_4218; // @[executor.scala 308:60]
  wire [7:0] _GEN_4539 = 8'h5 < length_1 ? _GEN_4379 : _GEN_4219; // @[executor.scala 308:60]
  wire [7:0] _GEN_4540 = 8'h5 < length_1 ? _GEN_4380 : _GEN_4220; // @[executor.scala 308:60]
  wire [7:0] _GEN_4541 = 8'h5 < length_1 ? _GEN_4381 : _GEN_4221; // @[executor.scala 308:60]
  wire [7:0] _GEN_4542 = 8'h5 < length_1 ? _GEN_4382 : _GEN_4222; // @[executor.scala 308:60]
  wire [7:0] _GEN_4543 = 8'h5 < length_1 ? _GEN_4383 : _GEN_4223; // @[executor.scala 308:60]
  wire [7:0] _GEN_4544 = 8'h5 < length_1 ? _GEN_4384 : _GEN_4224; // @[executor.scala 308:60]
  wire [7:0] _GEN_4545 = 8'h5 < length_1 ? _GEN_4385 : _GEN_4225; // @[executor.scala 308:60]
  wire [7:0] _GEN_4546 = 8'h5 < length_1 ? _GEN_4386 : _GEN_4226; // @[executor.scala 308:60]
  wire [7:0] _GEN_4547 = 8'h5 < length_1 ? _GEN_4387 : _GEN_4227; // @[executor.scala 308:60]
  wire [7:0] _GEN_4548 = 8'h5 < length_1 ? _GEN_4388 : _GEN_4228; // @[executor.scala 308:60]
  wire [7:0] _GEN_4549 = 8'h5 < length_1 ? _GEN_4389 : _GEN_4229; // @[executor.scala 308:60]
  wire [7:0] _GEN_4550 = 8'h5 < length_1 ? _GEN_4390 : _GEN_4230; // @[executor.scala 308:60]
  wire [7:0] _GEN_4551 = 8'h5 < length_1 ? _GEN_4391 : _GEN_4231; // @[executor.scala 308:60]
  wire [7:0] _GEN_4552 = 8'h5 < length_1 ? _GEN_4392 : _GEN_4232; // @[executor.scala 308:60]
  wire [7:0] _GEN_4553 = 8'h5 < length_1 ? _GEN_4393 : _GEN_4233; // @[executor.scala 308:60]
  wire [7:0] _GEN_4554 = 8'h5 < length_1 ? _GEN_4394 : _GEN_4234; // @[executor.scala 308:60]
  wire [7:0] _GEN_4555 = 8'h5 < length_1 ? _GEN_4395 : _GEN_4235; // @[executor.scala 308:60]
  wire [7:0] _GEN_4556 = 8'h5 < length_1 ? _GEN_4396 : _GEN_4236; // @[executor.scala 308:60]
  wire [7:0] _GEN_4557 = 8'h5 < length_1 ? _GEN_4397 : _GEN_4237; // @[executor.scala 308:60]
  wire [7:0] _GEN_4558 = 8'h5 < length_1 ? _GEN_4398 : _GEN_4238; // @[executor.scala 308:60]
  wire [7:0] _GEN_4559 = 8'h5 < length_1 ? _GEN_4399 : _GEN_4239; // @[executor.scala 308:60]
  wire [7:0] _GEN_4560 = 8'h5 < length_1 ? _GEN_4400 : _GEN_4240; // @[executor.scala 308:60]
  wire [7:0] _GEN_4561 = 8'h5 < length_1 ? _GEN_4401 : _GEN_4241; // @[executor.scala 308:60]
  wire [7:0] _GEN_4562 = 8'h5 < length_1 ? _GEN_4402 : _GEN_4242; // @[executor.scala 308:60]
  wire [7:0] _GEN_4563 = 8'h5 < length_1 ? _GEN_4403 : _GEN_4243; // @[executor.scala 308:60]
  wire [7:0] _GEN_4564 = 8'h5 < length_1 ? _GEN_4404 : _GEN_4244; // @[executor.scala 308:60]
  wire [7:0] _GEN_4565 = 8'h5 < length_1 ? _GEN_4405 : _GEN_4245; // @[executor.scala 308:60]
  wire [7:0] _GEN_4566 = 8'h5 < length_1 ? _GEN_4406 : _GEN_4246; // @[executor.scala 308:60]
  wire [7:0] _GEN_4567 = 8'h5 < length_1 ? _GEN_4407 : _GEN_4247; // @[executor.scala 308:60]
  wire [7:0] _GEN_4568 = 8'h5 < length_1 ? _GEN_4408 : _GEN_4248; // @[executor.scala 308:60]
  wire [7:0] _GEN_4569 = 8'h5 < length_1 ? _GEN_4409 : _GEN_4249; // @[executor.scala 308:60]
  wire [7:0] _GEN_4570 = 8'h5 < length_1 ? _GEN_4410 : _GEN_4250; // @[executor.scala 308:60]
  wire [7:0] _GEN_4571 = 8'h5 < length_1 ? _GEN_4411 : _GEN_4251; // @[executor.scala 308:60]
  wire [7:0] _GEN_4572 = 8'h5 < length_1 ? _GEN_4412 : _GEN_4252; // @[executor.scala 308:60]
  wire [7:0] _GEN_4573 = 8'h5 < length_1 ? _GEN_4413 : _GEN_4253; // @[executor.scala 308:60]
  wire [7:0] _GEN_4574 = 8'h5 < length_1 ? _GEN_4414 : _GEN_4254; // @[executor.scala 308:60]
  wire [7:0] _GEN_4575 = 8'h5 < length_1 ? _GEN_4415 : _GEN_4255; // @[executor.scala 308:60]
  wire [7:0] _GEN_4576 = 8'h5 < length_1 ? _GEN_4416 : _GEN_4256; // @[executor.scala 308:60]
  wire [7:0] _GEN_4577 = 8'h5 < length_1 ? _GEN_4417 : _GEN_4257; // @[executor.scala 308:60]
  wire [7:0] _GEN_4578 = 8'h5 < length_1 ? _GEN_4418 : _GEN_4258; // @[executor.scala 308:60]
  wire [7:0] _GEN_4579 = 8'h5 < length_1 ? _GEN_4419 : _GEN_4259; // @[executor.scala 308:60]
  wire [7:0] _GEN_4580 = 8'h5 < length_1 ? _GEN_4420 : _GEN_4260; // @[executor.scala 308:60]
  wire [7:0] _GEN_4581 = 8'h5 < length_1 ? _GEN_4421 : _GEN_4261; // @[executor.scala 308:60]
  wire [7:0] _GEN_4582 = 8'h5 < length_1 ? _GEN_4422 : _GEN_4262; // @[executor.scala 308:60]
  wire [7:0] _GEN_4583 = 8'h5 < length_1 ? _GEN_4423 : _GEN_4263; // @[executor.scala 308:60]
  wire [7:0] _GEN_4584 = 8'h5 < length_1 ? _GEN_4424 : _GEN_4264; // @[executor.scala 308:60]
  wire [7:0] _GEN_4585 = 8'h5 < length_1 ? _GEN_4425 : _GEN_4265; // @[executor.scala 308:60]
  wire [7:0] _GEN_4586 = 8'h5 < length_1 ? _GEN_4426 : _GEN_4266; // @[executor.scala 308:60]
  wire [7:0] _GEN_4587 = 8'h5 < length_1 ? _GEN_4427 : _GEN_4267; // @[executor.scala 308:60]
  wire [7:0] _GEN_4588 = 8'h5 < length_1 ? _GEN_4428 : _GEN_4268; // @[executor.scala 308:60]
  wire [7:0] _GEN_4589 = 8'h5 < length_1 ? _GEN_4429 : _GEN_4269; // @[executor.scala 308:60]
  wire [7:0] _GEN_4590 = 8'h5 < length_1 ? _GEN_4430 : _GEN_4270; // @[executor.scala 308:60]
  wire [7:0] _GEN_4591 = 8'h5 < length_1 ? _GEN_4431 : _GEN_4271; // @[executor.scala 308:60]
  wire [7:0] _GEN_4592 = 8'h5 < length_1 ? _GEN_4432 : _GEN_4272; // @[executor.scala 308:60]
  wire [7:0] _GEN_4593 = 8'h5 < length_1 ? _GEN_4433 : _GEN_4273; // @[executor.scala 308:60]
  wire [7:0] _GEN_4594 = 8'h5 < length_1 ? _GEN_4434 : _GEN_4274; // @[executor.scala 308:60]
  wire [7:0] _GEN_4595 = 8'h5 < length_1 ? _GEN_4435 : _GEN_4275; // @[executor.scala 308:60]
  wire [7:0] _GEN_4596 = 8'h5 < length_1 ? _GEN_4436 : _GEN_4276; // @[executor.scala 308:60]
  wire [7:0] _GEN_4597 = 8'h5 < length_1 ? _GEN_4437 : _GEN_4277; // @[executor.scala 308:60]
  wire [7:0] _GEN_4598 = 8'h5 < length_1 ? _GEN_4438 : _GEN_4278; // @[executor.scala 308:60]
  wire [7:0] _GEN_4599 = 8'h5 < length_1 ? _GEN_4439 : _GEN_4279; // @[executor.scala 308:60]
  wire [7:0] _GEN_4600 = 8'h5 < length_1 ? _GEN_4440 : _GEN_4280; // @[executor.scala 308:60]
  wire [7:0] _GEN_4601 = 8'h5 < length_1 ? _GEN_4441 : _GEN_4281; // @[executor.scala 308:60]
  wire [7:0] _GEN_4602 = 8'h5 < length_1 ? _GEN_4442 : _GEN_4282; // @[executor.scala 308:60]
  wire [7:0] _GEN_4603 = 8'h5 < length_1 ? _GEN_4443 : _GEN_4283; // @[executor.scala 308:60]
  wire [7:0] _GEN_4604 = 8'h5 < length_1 ? _GEN_4444 : _GEN_4284; // @[executor.scala 308:60]
  wire [7:0] _GEN_4605 = 8'h5 < length_1 ? _GEN_4445 : _GEN_4285; // @[executor.scala 308:60]
  wire [7:0] _GEN_4606 = 8'h5 < length_1 ? _GEN_4446 : _GEN_4286; // @[executor.scala 308:60]
  wire [7:0] _GEN_4607 = 8'h5 < length_1 ? _GEN_4447 : _GEN_4287; // @[executor.scala 308:60]
  wire [7:0] _GEN_4608 = 8'h5 < length_1 ? _GEN_4448 : _GEN_4288; // @[executor.scala 308:60]
  wire [7:0] _GEN_4609 = 8'h5 < length_1 ? _GEN_4449 : _GEN_4289; // @[executor.scala 308:60]
  wire [7:0] _GEN_4610 = 8'h5 < length_1 ? _GEN_4450 : _GEN_4290; // @[executor.scala 308:60]
  wire [7:0] _GEN_4611 = 8'h5 < length_1 ? _GEN_4451 : _GEN_4291; // @[executor.scala 308:60]
  wire [7:0] _GEN_4612 = 8'h5 < length_1 ? _GEN_4452 : _GEN_4292; // @[executor.scala 308:60]
  wire [7:0] _GEN_4613 = 8'h5 < length_1 ? _GEN_4453 : _GEN_4293; // @[executor.scala 308:60]
  wire [7:0] _GEN_4614 = 8'h5 < length_1 ? _GEN_4454 : _GEN_4294; // @[executor.scala 308:60]
  wire [7:0] _GEN_4615 = 8'h5 < length_1 ? _GEN_4455 : _GEN_4295; // @[executor.scala 308:60]
  wire [7:0] _GEN_4616 = 8'h5 < length_1 ? _GEN_4456 : _GEN_4296; // @[executor.scala 308:60]
  wire [7:0] _GEN_4617 = 8'h5 < length_1 ? _GEN_4457 : _GEN_4297; // @[executor.scala 308:60]
  wire [7:0] _GEN_4618 = 8'h5 < length_1 ? _GEN_4458 : _GEN_4298; // @[executor.scala 308:60]
  wire [7:0] _GEN_4619 = 8'h5 < length_1 ? _GEN_4459 : _GEN_4299; // @[executor.scala 308:60]
  wire [7:0] _GEN_4620 = 8'h5 < length_1 ? _GEN_4460 : _GEN_4300; // @[executor.scala 308:60]
  wire [7:0] _GEN_4621 = 8'h5 < length_1 ? _GEN_4461 : _GEN_4301; // @[executor.scala 308:60]
  wire [7:0] _GEN_4622 = 8'h5 < length_1 ? _GEN_4462 : _GEN_4302; // @[executor.scala 308:60]
  wire [7:0] _GEN_4623 = 8'h5 < length_1 ? _GEN_4463 : _GEN_4303; // @[executor.scala 308:60]
  wire [7:0] _GEN_4624 = 8'h5 < length_1 ? _GEN_4464 : _GEN_4304; // @[executor.scala 308:60]
  wire [7:0] _GEN_4625 = 8'h5 < length_1 ? _GEN_4465 : _GEN_4305; // @[executor.scala 308:60]
  wire [7:0] _GEN_4626 = 8'h5 < length_1 ? _GEN_4466 : _GEN_4306; // @[executor.scala 308:60]
  wire [7:0] _GEN_4627 = 8'h5 < length_1 ? _GEN_4467 : _GEN_4307; // @[executor.scala 308:60]
  wire [7:0] _GEN_4628 = 8'h5 < length_1 ? _GEN_4468 : _GEN_4308; // @[executor.scala 308:60]
  wire [7:0] _GEN_4629 = 8'h5 < length_1 ? _GEN_4469 : _GEN_4309; // @[executor.scala 308:60]
  wire [7:0] _GEN_4630 = 8'h5 < length_1 ? _GEN_4470 : _GEN_4310; // @[executor.scala 308:60]
  wire [7:0] _GEN_4631 = 8'h5 < length_1 ? _GEN_4471 : _GEN_4311; // @[executor.scala 308:60]
  wire [7:0] _GEN_4632 = 8'h5 < length_1 ? _GEN_4472 : _GEN_4312; // @[executor.scala 308:60]
  wire [7:0] _GEN_4633 = 8'h5 < length_1 ? _GEN_4473 : _GEN_4313; // @[executor.scala 308:60]
  wire [7:0] _GEN_4634 = 8'h5 < length_1 ? _GEN_4474 : _GEN_4314; // @[executor.scala 308:60]
  wire [7:0] _GEN_4635 = 8'h5 < length_1 ? _GEN_4475 : _GEN_4315; // @[executor.scala 308:60]
  wire [7:0] _GEN_4636 = 8'h5 < length_1 ? _GEN_4476 : _GEN_4316; // @[executor.scala 308:60]
  wire [7:0] _GEN_4637 = 8'h5 < length_1 ? _GEN_4477 : _GEN_4317; // @[executor.scala 308:60]
  wire [7:0] _GEN_4638 = 8'h5 < length_1 ? _GEN_4478 : _GEN_4318; // @[executor.scala 308:60]
  wire [7:0] _GEN_4639 = 8'h5 < length_1 ? _GEN_4479 : _GEN_4319; // @[executor.scala 308:60]
  wire [7:0] _GEN_4640 = 8'h5 < length_1 ? _GEN_4480 : _GEN_4320; // @[executor.scala 308:60]
  wire [7:0] _GEN_4641 = 8'h5 < length_1 ? _GEN_4481 : _GEN_4321; // @[executor.scala 308:60]
  wire [7:0] field_byte_14 = field_1[15:8]; // @[executor.scala 305:57]
  wire [7:0] total_offset_14 = offset_1 + 8'h6; // @[executor.scala 307:57]
  wire [7:0] _GEN_4642 = 8'h0 == total_offset_14 ? field_byte_14 : _GEN_4482; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4643 = 8'h1 == total_offset_14 ? field_byte_14 : _GEN_4483; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4644 = 8'h2 == total_offset_14 ? field_byte_14 : _GEN_4484; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4645 = 8'h3 == total_offset_14 ? field_byte_14 : _GEN_4485; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4646 = 8'h4 == total_offset_14 ? field_byte_14 : _GEN_4486; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4647 = 8'h5 == total_offset_14 ? field_byte_14 : _GEN_4487; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4648 = 8'h6 == total_offset_14 ? field_byte_14 : _GEN_4488; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4649 = 8'h7 == total_offset_14 ? field_byte_14 : _GEN_4489; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4650 = 8'h8 == total_offset_14 ? field_byte_14 : _GEN_4490; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4651 = 8'h9 == total_offset_14 ? field_byte_14 : _GEN_4491; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4652 = 8'ha == total_offset_14 ? field_byte_14 : _GEN_4492; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4653 = 8'hb == total_offset_14 ? field_byte_14 : _GEN_4493; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4654 = 8'hc == total_offset_14 ? field_byte_14 : _GEN_4494; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4655 = 8'hd == total_offset_14 ? field_byte_14 : _GEN_4495; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4656 = 8'he == total_offset_14 ? field_byte_14 : _GEN_4496; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4657 = 8'hf == total_offset_14 ? field_byte_14 : _GEN_4497; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4658 = 8'h10 == total_offset_14 ? field_byte_14 : _GEN_4498; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4659 = 8'h11 == total_offset_14 ? field_byte_14 : _GEN_4499; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4660 = 8'h12 == total_offset_14 ? field_byte_14 : _GEN_4500; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4661 = 8'h13 == total_offset_14 ? field_byte_14 : _GEN_4501; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4662 = 8'h14 == total_offset_14 ? field_byte_14 : _GEN_4502; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4663 = 8'h15 == total_offset_14 ? field_byte_14 : _GEN_4503; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4664 = 8'h16 == total_offset_14 ? field_byte_14 : _GEN_4504; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4665 = 8'h17 == total_offset_14 ? field_byte_14 : _GEN_4505; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4666 = 8'h18 == total_offset_14 ? field_byte_14 : _GEN_4506; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4667 = 8'h19 == total_offset_14 ? field_byte_14 : _GEN_4507; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4668 = 8'h1a == total_offset_14 ? field_byte_14 : _GEN_4508; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4669 = 8'h1b == total_offset_14 ? field_byte_14 : _GEN_4509; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4670 = 8'h1c == total_offset_14 ? field_byte_14 : _GEN_4510; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4671 = 8'h1d == total_offset_14 ? field_byte_14 : _GEN_4511; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4672 = 8'h1e == total_offset_14 ? field_byte_14 : _GEN_4512; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4673 = 8'h1f == total_offset_14 ? field_byte_14 : _GEN_4513; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4674 = 8'h20 == total_offset_14 ? field_byte_14 : _GEN_4514; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4675 = 8'h21 == total_offset_14 ? field_byte_14 : _GEN_4515; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4676 = 8'h22 == total_offset_14 ? field_byte_14 : _GEN_4516; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4677 = 8'h23 == total_offset_14 ? field_byte_14 : _GEN_4517; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4678 = 8'h24 == total_offset_14 ? field_byte_14 : _GEN_4518; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4679 = 8'h25 == total_offset_14 ? field_byte_14 : _GEN_4519; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4680 = 8'h26 == total_offset_14 ? field_byte_14 : _GEN_4520; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4681 = 8'h27 == total_offset_14 ? field_byte_14 : _GEN_4521; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4682 = 8'h28 == total_offset_14 ? field_byte_14 : _GEN_4522; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4683 = 8'h29 == total_offset_14 ? field_byte_14 : _GEN_4523; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4684 = 8'h2a == total_offset_14 ? field_byte_14 : _GEN_4524; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4685 = 8'h2b == total_offset_14 ? field_byte_14 : _GEN_4525; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4686 = 8'h2c == total_offset_14 ? field_byte_14 : _GEN_4526; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4687 = 8'h2d == total_offset_14 ? field_byte_14 : _GEN_4527; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4688 = 8'h2e == total_offset_14 ? field_byte_14 : _GEN_4528; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4689 = 8'h2f == total_offset_14 ? field_byte_14 : _GEN_4529; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4690 = 8'h30 == total_offset_14 ? field_byte_14 : _GEN_4530; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4691 = 8'h31 == total_offset_14 ? field_byte_14 : _GEN_4531; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4692 = 8'h32 == total_offset_14 ? field_byte_14 : _GEN_4532; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4693 = 8'h33 == total_offset_14 ? field_byte_14 : _GEN_4533; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4694 = 8'h34 == total_offset_14 ? field_byte_14 : _GEN_4534; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4695 = 8'h35 == total_offset_14 ? field_byte_14 : _GEN_4535; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4696 = 8'h36 == total_offset_14 ? field_byte_14 : _GEN_4536; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4697 = 8'h37 == total_offset_14 ? field_byte_14 : _GEN_4537; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4698 = 8'h38 == total_offset_14 ? field_byte_14 : _GEN_4538; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4699 = 8'h39 == total_offset_14 ? field_byte_14 : _GEN_4539; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4700 = 8'h3a == total_offset_14 ? field_byte_14 : _GEN_4540; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4701 = 8'h3b == total_offset_14 ? field_byte_14 : _GEN_4541; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4702 = 8'h3c == total_offset_14 ? field_byte_14 : _GEN_4542; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4703 = 8'h3d == total_offset_14 ? field_byte_14 : _GEN_4543; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4704 = 8'h3e == total_offset_14 ? field_byte_14 : _GEN_4544; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4705 = 8'h3f == total_offset_14 ? field_byte_14 : _GEN_4545; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4706 = 8'h40 == total_offset_14 ? field_byte_14 : _GEN_4546; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4707 = 8'h41 == total_offset_14 ? field_byte_14 : _GEN_4547; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4708 = 8'h42 == total_offset_14 ? field_byte_14 : _GEN_4548; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4709 = 8'h43 == total_offset_14 ? field_byte_14 : _GEN_4549; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4710 = 8'h44 == total_offset_14 ? field_byte_14 : _GEN_4550; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4711 = 8'h45 == total_offset_14 ? field_byte_14 : _GEN_4551; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4712 = 8'h46 == total_offset_14 ? field_byte_14 : _GEN_4552; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4713 = 8'h47 == total_offset_14 ? field_byte_14 : _GEN_4553; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4714 = 8'h48 == total_offset_14 ? field_byte_14 : _GEN_4554; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4715 = 8'h49 == total_offset_14 ? field_byte_14 : _GEN_4555; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4716 = 8'h4a == total_offset_14 ? field_byte_14 : _GEN_4556; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4717 = 8'h4b == total_offset_14 ? field_byte_14 : _GEN_4557; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4718 = 8'h4c == total_offset_14 ? field_byte_14 : _GEN_4558; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4719 = 8'h4d == total_offset_14 ? field_byte_14 : _GEN_4559; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4720 = 8'h4e == total_offset_14 ? field_byte_14 : _GEN_4560; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4721 = 8'h4f == total_offset_14 ? field_byte_14 : _GEN_4561; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4722 = 8'h50 == total_offset_14 ? field_byte_14 : _GEN_4562; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4723 = 8'h51 == total_offset_14 ? field_byte_14 : _GEN_4563; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4724 = 8'h52 == total_offset_14 ? field_byte_14 : _GEN_4564; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4725 = 8'h53 == total_offset_14 ? field_byte_14 : _GEN_4565; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4726 = 8'h54 == total_offset_14 ? field_byte_14 : _GEN_4566; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4727 = 8'h55 == total_offset_14 ? field_byte_14 : _GEN_4567; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4728 = 8'h56 == total_offset_14 ? field_byte_14 : _GEN_4568; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4729 = 8'h57 == total_offset_14 ? field_byte_14 : _GEN_4569; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4730 = 8'h58 == total_offset_14 ? field_byte_14 : _GEN_4570; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4731 = 8'h59 == total_offset_14 ? field_byte_14 : _GEN_4571; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4732 = 8'h5a == total_offset_14 ? field_byte_14 : _GEN_4572; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4733 = 8'h5b == total_offset_14 ? field_byte_14 : _GEN_4573; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4734 = 8'h5c == total_offset_14 ? field_byte_14 : _GEN_4574; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4735 = 8'h5d == total_offset_14 ? field_byte_14 : _GEN_4575; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4736 = 8'h5e == total_offset_14 ? field_byte_14 : _GEN_4576; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4737 = 8'h5f == total_offset_14 ? field_byte_14 : _GEN_4577; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4738 = 8'h60 == total_offset_14 ? field_byte_14 : _GEN_4578; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4739 = 8'h61 == total_offset_14 ? field_byte_14 : _GEN_4579; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4740 = 8'h62 == total_offset_14 ? field_byte_14 : _GEN_4580; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4741 = 8'h63 == total_offset_14 ? field_byte_14 : _GEN_4581; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4742 = 8'h64 == total_offset_14 ? field_byte_14 : _GEN_4582; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4743 = 8'h65 == total_offset_14 ? field_byte_14 : _GEN_4583; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4744 = 8'h66 == total_offset_14 ? field_byte_14 : _GEN_4584; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4745 = 8'h67 == total_offset_14 ? field_byte_14 : _GEN_4585; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4746 = 8'h68 == total_offset_14 ? field_byte_14 : _GEN_4586; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4747 = 8'h69 == total_offset_14 ? field_byte_14 : _GEN_4587; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4748 = 8'h6a == total_offset_14 ? field_byte_14 : _GEN_4588; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4749 = 8'h6b == total_offset_14 ? field_byte_14 : _GEN_4589; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4750 = 8'h6c == total_offset_14 ? field_byte_14 : _GEN_4590; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4751 = 8'h6d == total_offset_14 ? field_byte_14 : _GEN_4591; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4752 = 8'h6e == total_offset_14 ? field_byte_14 : _GEN_4592; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4753 = 8'h6f == total_offset_14 ? field_byte_14 : _GEN_4593; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4754 = 8'h70 == total_offset_14 ? field_byte_14 : _GEN_4594; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4755 = 8'h71 == total_offset_14 ? field_byte_14 : _GEN_4595; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4756 = 8'h72 == total_offset_14 ? field_byte_14 : _GEN_4596; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4757 = 8'h73 == total_offset_14 ? field_byte_14 : _GEN_4597; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4758 = 8'h74 == total_offset_14 ? field_byte_14 : _GEN_4598; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4759 = 8'h75 == total_offset_14 ? field_byte_14 : _GEN_4599; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4760 = 8'h76 == total_offset_14 ? field_byte_14 : _GEN_4600; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4761 = 8'h77 == total_offset_14 ? field_byte_14 : _GEN_4601; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4762 = 8'h78 == total_offset_14 ? field_byte_14 : _GEN_4602; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4763 = 8'h79 == total_offset_14 ? field_byte_14 : _GEN_4603; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4764 = 8'h7a == total_offset_14 ? field_byte_14 : _GEN_4604; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4765 = 8'h7b == total_offset_14 ? field_byte_14 : _GEN_4605; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4766 = 8'h7c == total_offset_14 ? field_byte_14 : _GEN_4606; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4767 = 8'h7d == total_offset_14 ? field_byte_14 : _GEN_4607; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4768 = 8'h7e == total_offset_14 ? field_byte_14 : _GEN_4608; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4769 = 8'h7f == total_offset_14 ? field_byte_14 : _GEN_4609; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4770 = 8'h80 == total_offset_14 ? field_byte_14 : _GEN_4610; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4771 = 8'h81 == total_offset_14 ? field_byte_14 : _GEN_4611; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4772 = 8'h82 == total_offset_14 ? field_byte_14 : _GEN_4612; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4773 = 8'h83 == total_offset_14 ? field_byte_14 : _GEN_4613; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4774 = 8'h84 == total_offset_14 ? field_byte_14 : _GEN_4614; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4775 = 8'h85 == total_offset_14 ? field_byte_14 : _GEN_4615; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4776 = 8'h86 == total_offset_14 ? field_byte_14 : _GEN_4616; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4777 = 8'h87 == total_offset_14 ? field_byte_14 : _GEN_4617; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4778 = 8'h88 == total_offset_14 ? field_byte_14 : _GEN_4618; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4779 = 8'h89 == total_offset_14 ? field_byte_14 : _GEN_4619; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4780 = 8'h8a == total_offset_14 ? field_byte_14 : _GEN_4620; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4781 = 8'h8b == total_offset_14 ? field_byte_14 : _GEN_4621; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4782 = 8'h8c == total_offset_14 ? field_byte_14 : _GEN_4622; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4783 = 8'h8d == total_offset_14 ? field_byte_14 : _GEN_4623; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4784 = 8'h8e == total_offset_14 ? field_byte_14 : _GEN_4624; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4785 = 8'h8f == total_offset_14 ? field_byte_14 : _GEN_4625; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4786 = 8'h90 == total_offset_14 ? field_byte_14 : _GEN_4626; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4787 = 8'h91 == total_offset_14 ? field_byte_14 : _GEN_4627; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4788 = 8'h92 == total_offset_14 ? field_byte_14 : _GEN_4628; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4789 = 8'h93 == total_offset_14 ? field_byte_14 : _GEN_4629; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4790 = 8'h94 == total_offset_14 ? field_byte_14 : _GEN_4630; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4791 = 8'h95 == total_offset_14 ? field_byte_14 : _GEN_4631; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4792 = 8'h96 == total_offset_14 ? field_byte_14 : _GEN_4632; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4793 = 8'h97 == total_offset_14 ? field_byte_14 : _GEN_4633; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4794 = 8'h98 == total_offset_14 ? field_byte_14 : _GEN_4634; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4795 = 8'h99 == total_offset_14 ? field_byte_14 : _GEN_4635; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4796 = 8'h9a == total_offset_14 ? field_byte_14 : _GEN_4636; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4797 = 8'h9b == total_offset_14 ? field_byte_14 : _GEN_4637; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4798 = 8'h9c == total_offset_14 ? field_byte_14 : _GEN_4638; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4799 = 8'h9d == total_offset_14 ? field_byte_14 : _GEN_4639; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4800 = 8'h9e == total_offset_14 ? field_byte_14 : _GEN_4640; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4801 = 8'h9f == total_offset_14 ? field_byte_14 : _GEN_4641; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4802 = 8'h6 < length_1 ? _GEN_4642 : _GEN_4482; // @[executor.scala 308:60]
  wire [7:0] _GEN_4803 = 8'h6 < length_1 ? _GEN_4643 : _GEN_4483; // @[executor.scala 308:60]
  wire [7:0] _GEN_4804 = 8'h6 < length_1 ? _GEN_4644 : _GEN_4484; // @[executor.scala 308:60]
  wire [7:0] _GEN_4805 = 8'h6 < length_1 ? _GEN_4645 : _GEN_4485; // @[executor.scala 308:60]
  wire [7:0] _GEN_4806 = 8'h6 < length_1 ? _GEN_4646 : _GEN_4486; // @[executor.scala 308:60]
  wire [7:0] _GEN_4807 = 8'h6 < length_1 ? _GEN_4647 : _GEN_4487; // @[executor.scala 308:60]
  wire [7:0] _GEN_4808 = 8'h6 < length_1 ? _GEN_4648 : _GEN_4488; // @[executor.scala 308:60]
  wire [7:0] _GEN_4809 = 8'h6 < length_1 ? _GEN_4649 : _GEN_4489; // @[executor.scala 308:60]
  wire [7:0] _GEN_4810 = 8'h6 < length_1 ? _GEN_4650 : _GEN_4490; // @[executor.scala 308:60]
  wire [7:0] _GEN_4811 = 8'h6 < length_1 ? _GEN_4651 : _GEN_4491; // @[executor.scala 308:60]
  wire [7:0] _GEN_4812 = 8'h6 < length_1 ? _GEN_4652 : _GEN_4492; // @[executor.scala 308:60]
  wire [7:0] _GEN_4813 = 8'h6 < length_1 ? _GEN_4653 : _GEN_4493; // @[executor.scala 308:60]
  wire [7:0] _GEN_4814 = 8'h6 < length_1 ? _GEN_4654 : _GEN_4494; // @[executor.scala 308:60]
  wire [7:0] _GEN_4815 = 8'h6 < length_1 ? _GEN_4655 : _GEN_4495; // @[executor.scala 308:60]
  wire [7:0] _GEN_4816 = 8'h6 < length_1 ? _GEN_4656 : _GEN_4496; // @[executor.scala 308:60]
  wire [7:0] _GEN_4817 = 8'h6 < length_1 ? _GEN_4657 : _GEN_4497; // @[executor.scala 308:60]
  wire [7:0] _GEN_4818 = 8'h6 < length_1 ? _GEN_4658 : _GEN_4498; // @[executor.scala 308:60]
  wire [7:0] _GEN_4819 = 8'h6 < length_1 ? _GEN_4659 : _GEN_4499; // @[executor.scala 308:60]
  wire [7:0] _GEN_4820 = 8'h6 < length_1 ? _GEN_4660 : _GEN_4500; // @[executor.scala 308:60]
  wire [7:0] _GEN_4821 = 8'h6 < length_1 ? _GEN_4661 : _GEN_4501; // @[executor.scala 308:60]
  wire [7:0] _GEN_4822 = 8'h6 < length_1 ? _GEN_4662 : _GEN_4502; // @[executor.scala 308:60]
  wire [7:0] _GEN_4823 = 8'h6 < length_1 ? _GEN_4663 : _GEN_4503; // @[executor.scala 308:60]
  wire [7:0] _GEN_4824 = 8'h6 < length_1 ? _GEN_4664 : _GEN_4504; // @[executor.scala 308:60]
  wire [7:0] _GEN_4825 = 8'h6 < length_1 ? _GEN_4665 : _GEN_4505; // @[executor.scala 308:60]
  wire [7:0] _GEN_4826 = 8'h6 < length_1 ? _GEN_4666 : _GEN_4506; // @[executor.scala 308:60]
  wire [7:0] _GEN_4827 = 8'h6 < length_1 ? _GEN_4667 : _GEN_4507; // @[executor.scala 308:60]
  wire [7:0] _GEN_4828 = 8'h6 < length_1 ? _GEN_4668 : _GEN_4508; // @[executor.scala 308:60]
  wire [7:0] _GEN_4829 = 8'h6 < length_1 ? _GEN_4669 : _GEN_4509; // @[executor.scala 308:60]
  wire [7:0] _GEN_4830 = 8'h6 < length_1 ? _GEN_4670 : _GEN_4510; // @[executor.scala 308:60]
  wire [7:0] _GEN_4831 = 8'h6 < length_1 ? _GEN_4671 : _GEN_4511; // @[executor.scala 308:60]
  wire [7:0] _GEN_4832 = 8'h6 < length_1 ? _GEN_4672 : _GEN_4512; // @[executor.scala 308:60]
  wire [7:0] _GEN_4833 = 8'h6 < length_1 ? _GEN_4673 : _GEN_4513; // @[executor.scala 308:60]
  wire [7:0] _GEN_4834 = 8'h6 < length_1 ? _GEN_4674 : _GEN_4514; // @[executor.scala 308:60]
  wire [7:0] _GEN_4835 = 8'h6 < length_1 ? _GEN_4675 : _GEN_4515; // @[executor.scala 308:60]
  wire [7:0] _GEN_4836 = 8'h6 < length_1 ? _GEN_4676 : _GEN_4516; // @[executor.scala 308:60]
  wire [7:0] _GEN_4837 = 8'h6 < length_1 ? _GEN_4677 : _GEN_4517; // @[executor.scala 308:60]
  wire [7:0] _GEN_4838 = 8'h6 < length_1 ? _GEN_4678 : _GEN_4518; // @[executor.scala 308:60]
  wire [7:0] _GEN_4839 = 8'h6 < length_1 ? _GEN_4679 : _GEN_4519; // @[executor.scala 308:60]
  wire [7:0] _GEN_4840 = 8'h6 < length_1 ? _GEN_4680 : _GEN_4520; // @[executor.scala 308:60]
  wire [7:0] _GEN_4841 = 8'h6 < length_1 ? _GEN_4681 : _GEN_4521; // @[executor.scala 308:60]
  wire [7:0] _GEN_4842 = 8'h6 < length_1 ? _GEN_4682 : _GEN_4522; // @[executor.scala 308:60]
  wire [7:0] _GEN_4843 = 8'h6 < length_1 ? _GEN_4683 : _GEN_4523; // @[executor.scala 308:60]
  wire [7:0] _GEN_4844 = 8'h6 < length_1 ? _GEN_4684 : _GEN_4524; // @[executor.scala 308:60]
  wire [7:0] _GEN_4845 = 8'h6 < length_1 ? _GEN_4685 : _GEN_4525; // @[executor.scala 308:60]
  wire [7:0] _GEN_4846 = 8'h6 < length_1 ? _GEN_4686 : _GEN_4526; // @[executor.scala 308:60]
  wire [7:0] _GEN_4847 = 8'h6 < length_1 ? _GEN_4687 : _GEN_4527; // @[executor.scala 308:60]
  wire [7:0] _GEN_4848 = 8'h6 < length_1 ? _GEN_4688 : _GEN_4528; // @[executor.scala 308:60]
  wire [7:0] _GEN_4849 = 8'h6 < length_1 ? _GEN_4689 : _GEN_4529; // @[executor.scala 308:60]
  wire [7:0] _GEN_4850 = 8'h6 < length_1 ? _GEN_4690 : _GEN_4530; // @[executor.scala 308:60]
  wire [7:0] _GEN_4851 = 8'h6 < length_1 ? _GEN_4691 : _GEN_4531; // @[executor.scala 308:60]
  wire [7:0] _GEN_4852 = 8'h6 < length_1 ? _GEN_4692 : _GEN_4532; // @[executor.scala 308:60]
  wire [7:0] _GEN_4853 = 8'h6 < length_1 ? _GEN_4693 : _GEN_4533; // @[executor.scala 308:60]
  wire [7:0] _GEN_4854 = 8'h6 < length_1 ? _GEN_4694 : _GEN_4534; // @[executor.scala 308:60]
  wire [7:0] _GEN_4855 = 8'h6 < length_1 ? _GEN_4695 : _GEN_4535; // @[executor.scala 308:60]
  wire [7:0] _GEN_4856 = 8'h6 < length_1 ? _GEN_4696 : _GEN_4536; // @[executor.scala 308:60]
  wire [7:0] _GEN_4857 = 8'h6 < length_1 ? _GEN_4697 : _GEN_4537; // @[executor.scala 308:60]
  wire [7:0] _GEN_4858 = 8'h6 < length_1 ? _GEN_4698 : _GEN_4538; // @[executor.scala 308:60]
  wire [7:0] _GEN_4859 = 8'h6 < length_1 ? _GEN_4699 : _GEN_4539; // @[executor.scala 308:60]
  wire [7:0] _GEN_4860 = 8'h6 < length_1 ? _GEN_4700 : _GEN_4540; // @[executor.scala 308:60]
  wire [7:0] _GEN_4861 = 8'h6 < length_1 ? _GEN_4701 : _GEN_4541; // @[executor.scala 308:60]
  wire [7:0] _GEN_4862 = 8'h6 < length_1 ? _GEN_4702 : _GEN_4542; // @[executor.scala 308:60]
  wire [7:0] _GEN_4863 = 8'h6 < length_1 ? _GEN_4703 : _GEN_4543; // @[executor.scala 308:60]
  wire [7:0] _GEN_4864 = 8'h6 < length_1 ? _GEN_4704 : _GEN_4544; // @[executor.scala 308:60]
  wire [7:0] _GEN_4865 = 8'h6 < length_1 ? _GEN_4705 : _GEN_4545; // @[executor.scala 308:60]
  wire [7:0] _GEN_4866 = 8'h6 < length_1 ? _GEN_4706 : _GEN_4546; // @[executor.scala 308:60]
  wire [7:0] _GEN_4867 = 8'h6 < length_1 ? _GEN_4707 : _GEN_4547; // @[executor.scala 308:60]
  wire [7:0] _GEN_4868 = 8'h6 < length_1 ? _GEN_4708 : _GEN_4548; // @[executor.scala 308:60]
  wire [7:0] _GEN_4869 = 8'h6 < length_1 ? _GEN_4709 : _GEN_4549; // @[executor.scala 308:60]
  wire [7:0] _GEN_4870 = 8'h6 < length_1 ? _GEN_4710 : _GEN_4550; // @[executor.scala 308:60]
  wire [7:0] _GEN_4871 = 8'h6 < length_1 ? _GEN_4711 : _GEN_4551; // @[executor.scala 308:60]
  wire [7:0] _GEN_4872 = 8'h6 < length_1 ? _GEN_4712 : _GEN_4552; // @[executor.scala 308:60]
  wire [7:0] _GEN_4873 = 8'h6 < length_1 ? _GEN_4713 : _GEN_4553; // @[executor.scala 308:60]
  wire [7:0] _GEN_4874 = 8'h6 < length_1 ? _GEN_4714 : _GEN_4554; // @[executor.scala 308:60]
  wire [7:0] _GEN_4875 = 8'h6 < length_1 ? _GEN_4715 : _GEN_4555; // @[executor.scala 308:60]
  wire [7:0] _GEN_4876 = 8'h6 < length_1 ? _GEN_4716 : _GEN_4556; // @[executor.scala 308:60]
  wire [7:0] _GEN_4877 = 8'h6 < length_1 ? _GEN_4717 : _GEN_4557; // @[executor.scala 308:60]
  wire [7:0] _GEN_4878 = 8'h6 < length_1 ? _GEN_4718 : _GEN_4558; // @[executor.scala 308:60]
  wire [7:0] _GEN_4879 = 8'h6 < length_1 ? _GEN_4719 : _GEN_4559; // @[executor.scala 308:60]
  wire [7:0] _GEN_4880 = 8'h6 < length_1 ? _GEN_4720 : _GEN_4560; // @[executor.scala 308:60]
  wire [7:0] _GEN_4881 = 8'h6 < length_1 ? _GEN_4721 : _GEN_4561; // @[executor.scala 308:60]
  wire [7:0] _GEN_4882 = 8'h6 < length_1 ? _GEN_4722 : _GEN_4562; // @[executor.scala 308:60]
  wire [7:0] _GEN_4883 = 8'h6 < length_1 ? _GEN_4723 : _GEN_4563; // @[executor.scala 308:60]
  wire [7:0] _GEN_4884 = 8'h6 < length_1 ? _GEN_4724 : _GEN_4564; // @[executor.scala 308:60]
  wire [7:0] _GEN_4885 = 8'h6 < length_1 ? _GEN_4725 : _GEN_4565; // @[executor.scala 308:60]
  wire [7:0] _GEN_4886 = 8'h6 < length_1 ? _GEN_4726 : _GEN_4566; // @[executor.scala 308:60]
  wire [7:0] _GEN_4887 = 8'h6 < length_1 ? _GEN_4727 : _GEN_4567; // @[executor.scala 308:60]
  wire [7:0] _GEN_4888 = 8'h6 < length_1 ? _GEN_4728 : _GEN_4568; // @[executor.scala 308:60]
  wire [7:0] _GEN_4889 = 8'h6 < length_1 ? _GEN_4729 : _GEN_4569; // @[executor.scala 308:60]
  wire [7:0] _GEN_4890 = 8'h6 < length_1 ? _GEN_4730 : _GEN_4570; // @[executor.scala 308:60]
  wire [7:0] _GEN_4891 = 8'h6 < length_1 ? _GEN_4731 : _GEN_4571; // @[executor.scala 308:60]
  wire [7:0] _GEN_4892 = 8'h6 < length_1 ? _GEN_4732 : _GEN_4572; // @[executor.scala 308:60]
  wire [7:0] _GEN_4893 = 8'h6 < length_1 ? _GEN_4733 : _GEN_4573; // @[executor.scala 308:60]
  wire [7:0] _GEN_4894 = 8'h6 < length_1 ? _GEN_4734 : _GEN_4574; // @[executor.scala 308:60]
  wire [7:0] _GEN_4895 = 8'h6 < length_1 ? _GEN_4735 : _GEN_4575; // @[executor.scala 308:60]
  wire [7:0] _GEN_4896 = 8'h6 < length_1 ? _GEN_4736 : _GEN_4576; // @[executor.scala 308:60]
  wire [7:0] _GEN_4897 = 8'h6 < length_1 ? _GEN_4737 : _GEN_4577; // @[executor.scala 308:60]
  wire [7:0] _GEN_4898 = 8'h6 < length_1 ? _GEN_4738 : _GEN_4578; // @[executor.scala 308:60]
  wire [7:0] _GEN_4899 = 8'h6 < length_1 ? _GEN_4739 : _GEN_4579; // @[executor.scala 308:60]
  wire [7:0] _GEN_4900 = 8'h6 < length_1 ? _GEN_4740 : _GEN_4580; // @[executor.scala 308:60]
  wire [7:0] _GEN_4901 = 8'h6 < length_1 ? _GEN_4741 : _GEN_4581; // @[executor.scala 308:60]
  wire [7:0] _GEN_4902 = 8'h6 < length_1 ? _GEN_4742 : _GEN_4582; // @[executor.scala 308:60]
  wire [7:0] _GEN_4903 = 8'h6 < length_1 ? _GEN_4743 : _GEN_4583; // @[executor.scala 308:60]
  wire [7:0] _GEN_4904 = 8'h6 < length_1 ? _GEN_4744 : _GEN_4584; // @[executor.scala 308:60]
  wire [7:0] _GEN_4905 = 8'h6 < length_1 ? _GEN_4745 : _GEN_4585; // @[executor.scala 308:60]
  wire [7:0] _GEN_4906 = 8'h6 < length_1 ? _GEN_4746 : _GEN_4586; // @[executor.scala 308:60]
  wire [7:0] _GEN_4907 = 8'h6 < length_1 ? _GEN_4747 : _GEN_4587; // @[executor.scala 308:60]
  wire [7:0] _GEN_4908 = 8'h6 < length_1 ? _GEN_4748 : _GEN_4588; // @[executor.scala 308:60]
  wire [7:0] _GEN_4909 = 8'h6 < length_1 ? _GEN_4749 : _GEN_4589; // @[executor.scala 308:60]
  wire [7:0] _GEN_4910 = 8'h6 < length_1 ? _GEN_4750 : _GEN_4590; // @[executor.scala 308:60]
  wire [7:0] _GEN_4911 = 8'h6 < length_1 ? _GEN_4751 : _GEN_4591; // @[executor.scala 308:60]
  wire [7:0] _GEN_4912 = 8'h6 < length_1 ? _GEN_4752 : _GEN_4592; // @[executor.scala 308:60]
  wire [7:0] _GEN_4913 = 8'h6 < length_1 ? _GEN_4753 : _GEN_4593; // @[executor.scala 308:60]
  wire [7:0] _GEN_4914 = 8'h6 < length_1 ? _GEN_4754 : _GEN_4594; // @[executor.scala 308:60]
  wire [7:0] _GEN_4915 = 8'h6 < length_1 ? _GEN_4755 : _GEN_4595; // @[executor.scala 308:60]
  wire [7:0] _GEN_4916 = 8'h6 < length_1 ? _GEN_4756 : _GEN_4596; // @[executor.scala 308:60]
  wire [7:0] _GEN_4917 = 8'h6 < length_1 ? _GEN_4757 : _GEN_4597; // @[executor.scala 308:60]
  wire [7:0] _GEN_4918 = 8'h6 < length_1 ? _GEN_4758 : _GEN_4598; // @[executor.scala 308:60]
  wire [7:0] _GEN_4919 = 8'h6 < length_1 ? _GEN_4759 : _GEN_4599; // @[executor.scala 308:60]
  wire [7:0] _GEN_4920 = 8'h6 < length_1 ? _GEN_4760 : _GEN_4600; // @[executor.scala 308:60]
  wire [7:0] _GEN_4921 = 8'h6 < length_1 ? _GEN_4761 : _GEN_4601; // @[executor.scala 308:60]
  wire [7:0] _GEN_4922 = 8'h6 < length_1 ? _GEN_4762 : _GEN_4602; // @[executor.scala 308:60]
  wire [7:0] _GEN_4923 = 8'h6 < length_1 ? _GEN_4763 : _GEN_4603; // @[executor.scala 308:60]
  wire [7:0] _GEN_4924 = 8'h6 < length_1 ? _GEN_4764 : _GEN_4604; // @[executor.scala 308:60]
  wire [7:0] _GEN_4925 = 8'h6 < length_1 ? _GEN_4765 : _GEN_4605; // @[executor.scala 308:60]
  wire [7:0] _GEN_4926 = 8'h6 < length_1 ? _GEN_4766 : _GEN_4606; // @[executor.scala 308:60]
  wire [7:0] _GEN_4927 = 8'h6 < length_1 ? _GEN_4767 : _GEN_4607; // @[executor.scala 308:60]
  wire [7:0] _GEN_4928 = 8'h6 < length_1 ? _GEN_4768 : _GEN_4608; // @[executor.scala 308:60]
  wire [7:0] _GEN_4929 = 8'h6 < length_1 ? _GEN_4769 : _GEN_4609; // @[executor.scala 308:60]
  wire [7:0] _GEN_4930 = 8'h6 < length_1 ? _GEN_4770 : _GEN_4610; // @[executor.scala 308:60]
  wire [7:0] _GEN_4931 = 8'h6 < length_1 ? _GEN_4771 : _GEN_4611; // @[executor.scala 308:60]
  wire [7:0] _GEN_4932 = 8'h6 < length_1 ? _GEN_4772 : _GEN_4612; // @[executor.scala 308:60]
  wire [7:0] _GEN_4933 = 8'h6 < length_1 ? _GEN_4773 : _GEN_4613; // @[executor.scala 308:60]
  wire [7:0] _GEN_4934 = 8'h6 < length_1 ? _GEN_4774 : _GEN_4614; // @[executor.scala 308:60]
  wire [7:0] _GEN_4935 = 8'h6 < length_1 ? _GEN_4775 : _GEN_4615; // @[executor.scala 308:60]
  wire [7:0] _GEN_4936 = 8'h6 < length_1 ? _GEN_4776 : _GEN_4616; // @[executor.scala 308:60]
  wire [7:0] _GEN_4937 = 8'h6 < length_1 ? _GEN_4777 : _GEN_4617; // @[executor.scala 308:60]
  wire [7:0] _GEN_4938 = 8'h6 < length_1 ? _GEN_4778 : _GEN_4618; // @[executor.scala 308:60]
  wire [7:0] _GEN_4939 = 8'h6 < length_1 ? _GEN_4779 : _GEN_4619; // @[executor.scala 308:60]
  wire [7:0] _GEN_4940 = 8'h6 < length_1 ? _GEN_4780 : _GEN_4620; // @[executor.scala 308:60]
  wire [7:0] _GEN_4941 = 8'h6 < length_1 ? _GEN_4781 : _GEN_4621; // @[executor.scala 308:60]
  wire [7:0] _GEN_4942 = 8'h6 < length_1 ? _GEN_4782 : _GEN_4622; // @[executor.scala 308:60]
  wire [7:0] _GEN_4943 = 8'h6 < length_1 ? _GEN_4783 : _GEN_4623; // @[executor.scala 308:60]
  wire [7:0] _GEN_4944 = 8'h6 < length_1 ? _GEN_4784 : _GEN_4624; // @[executor.scala 308:60]
  wire [7:0] _GEN_4945 = 8'h6 < length_1 ? _GEN_4785 : _GEN_4625; // @[executor.scala 308:60]
  wire [7:0] _GEN_4946 = 8'h6 < length_1 ? _GEN_4786 : _GEN_4626; // @[executor.scala 308:60]
  wire [7:0] _GEN_4947 = 8'h6 < length_1 ? _GEN_4787 : _GEN_4627; // @[executor.scala 308:60]
  wire [7:0] _GEN_4948 = 8'h6 < length_1 ? _GEN_4788 : _GEN_4628; // @[executor.scala 308:60]
  wire [7:0] _GEN_4949 = 8'h6 < length_1 ? _GEN_4789 : _GEN_4629; // @[executor.scala 308:60]
  wire [7:0] _GEN_4950 = 8'h6 < length_1 ? _GEN_4790 : _GEN_4630; // @[executor.scala 308:60]
  wire [7:0] _GEN_4951 = 8'h6 < length_1 ? _GEN_4791 : _GEN_4631; // @[executor.scala 308:60]
  wire [7:0] _GEN_4952 = 8'h6 < length_1 ? _GEN_4792 : _GEN_4632; // @[executor.scala 308:60]
  wire [7:0] _GEN_4953 = 8'h6 < length_1 ? _GEN_4793 : _GEN_4633; // @[executor.scala 308:60]
  wire [7:0] _GEN_4954 = 8'h6 < length_1 ? _GEN_4794 : _GEN_4634; // @[executor.scala 308:60]
  wire [7:0] _GEN_4955 = 8'h6 < length_1 ? _GEN_4795 : _GEN_4635; // @[executor.scala 308:60]
  wire [7:0] _GEN_4956 = 8'h6 < length_1 ? _GEN_4796 : _GEN_4636; // @[executor.scala 308:60]
  wire [7:0] _GEN_4957 = 8'h6 < length_1 ? _GEN_4797 : _GEN_4637; // @[executor.scala 308:60]
  wire [7:0] _GEN_4958 = 8'h6 < length_1 ? _GEN_4798 : _GEN_4638; // @[executor.scala 308:60]
  wire [7:0] _GEN_4959 = 8'h6 < length_1 ? _GEN_4799 : _GEN_4639; // @[executor.scala 308:60]
  wire [7:0] _GEN_4960 = 8'h6 < length_1 ? _GEN_4800 : _GEN_4640; // @[executor.scala 308:60]
  wire [7:0] _GEN_4961 = 8'h6 < length_1 ? _GEN_4801 : _GEN_4641; // @[executor.scala 308:60]
  wire [7:0] field_byte_15 = field_1[7:0]; // @[executor.scala 305:57]
  wire [7:0] total_offset_15 = offset_1 + 8'h7; // @[executor.scala 307:57]
  wire [7:0] _GEN_4962 = 8'h0 == total_offset_15 ? field_byte_15 : _GEN_4802; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4963 = 8'h1 == total_offset_15 ? field_byte_15 : _GEN_4803; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4964 = 8'h2 == total_offset_15 ? field_byte_15 : _GEN_4804; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4965 = 8'h3 == total_offset_15 ? field_byte_15 : _GEN_4805; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4966 = 8'h4 == total_offset_15 ? field_byte_15 : _GEN_4806; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4967 = 8'h5 == total_offset_15 ? field_byte_15 : _GEN_4807; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4968 = 8'h6 == total_offset_15 ? field_byte_15 : _GEN_4808; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4969 = 8'h7 == total_offset_15 ? field_byte_15 : _GEN_4809; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4970 = 8'h8 == total_offset_15 ? field_byte_15 : _GEN_4810; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4971 = 8'h9 == total_offset_15 ? field_byte_15 : _GEN_4811; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4972 = 8'ha == total_offset_15 ? field_byte_15 : _GEN_4812; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4973 = 8'hb == total_offset_15 ? field_byte_15 : _GEN_4813; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4974 = 8'hc == total_offset_15 ? field_byte_15 : _GEN_4814; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4975 = 8'hd == total_offset_15 ? field_byte_15 : _GEN_4815; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4976 = 8'he == total_offset_15 ? field_byte_15 : _GEN_4816; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4977 = 8'hf == total_offset_15 ? field_byte_15 : _GEN_4817; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4978 = 8'h10 == total_offset_15 ? field_byte_15 : _GEN_4818; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4979 = 8'h11 == total_offset_15 ? field_byte_15 : _GEN_4819; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4980 = 8'h12 == total_offset_15 ? field_byte_15 : _GEN_4820; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4981 = 8'h13 == total_offset_15 ? field_byte_15 : _GEN_4821; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4982 = 8'h14 == total_offset_15 ? field_byte_15 : _GEN_4822; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4983 = 8'h15 == total_offset_15 ? field_byte_15 : _GEN_4823; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4984 = 8'h16 == total_offset_15 ? field_byte_15 : _GEN_4824; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4985 = 8'h17 == total_offset_15 ? field_byte_15 : _GEN_4825; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4986 = 8'h18 == total_offset_15 ? field_byte_15 : _GEN_4826; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4987 = 8'h19 == total_offset_15 ? field_byte_15 : _GEN_4827; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4988 = 8'h1a == total_offset_15 ? field_byte_15 : _GEN_4828; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4989 = 8'h1b == total_offset_15 ? field_byte_15 : _GEN_4829; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4990 = 8'h1c == total_offset_15 ? field_byte_15 : _GEN_4830; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4991 = 8'h1d == total_offset_15 ? field_byte_15 : _GEN_4831; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4992 = 8'h1e == total_offset_15 ? field_byte_15 : _GEN_4832; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4993 = 8'h1f == total_offset_15 ? field_byte_15 : _GEN_4833; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4994 = 8'h20 == total_offset_15 ? field_byte_15 : _GEN_4834; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4995 = 8'h21 == total_offset_15 ? field_byte_15 : _GEN_4835; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4996 = 8'h22 == total_offset_15 ? field_byte_15 : _GEN_4836; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4997 = 8'h23 == total_offset_15 ? field_byte_15 : _GEN_4837; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4998 = 8'h24 == total_offset_15 ? field_byte_15 : _GEN_4838; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_4999 = 8'h25 == total_offset_15 ? field_byte_15 : _GEN_4839; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5000 = 8'h26 == total_offset_15 ? field_byte_15 : _GEN_4840; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5001 = 8'h27 == total_offset_15 ? field_byte_15 : _GEN_4841; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5002 = 8'h28 == total_offset_15 ? field_byte_15 : _GEN_4842; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5003 = 8'h29 == total_offset_15 ? field_byte_15 : _GEN_4843; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5004 = 8'h2a == total_offset_15 ? field_byte_15 : _GEN_4844; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5005 = 8'h2b == total_offset_15 ? field_byte_15 : _GEN_4845; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5006 = 8'h2c == total_offset_15 ? field_byte_15 : _GEN_4846; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5007 = 8'h2d == total_offset_15 ? field_byte_15 : _GEN_4847; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5008 = 8'h2e == total_offset_15 ? field_byte_15 : _GEN_4848; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5009 = 8'h2f == total_offset_15 ? field_byte_15 : _GEN_4849; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5010 = 8'h30 == total_offset_15 ? field_byte_15 : _GEN_4850; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5011 = 8'h31 == total_offset_15 ? field_byte_15 : _GEN_4851; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5012 = 8'h32 == total_offset_15 ? field_byte_15 : _GEN_4852; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5013 = 8'h33 == total_offset_15 ? field_byte_15 : _GEN_4853; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5014 = 8'h34 == total_offset_15 ? field_byte_15 : _GEN_4854; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5015 = 8'h35 == total_offset_15 ? field_byte_15 : _GEN_4855; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5016 = 8'h36 == total_offset_15 ? field_byte_15 : _GEN_4856; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5017 = 8'h37 == total_offset_15 ? field_byte_15 : _GEN_4857; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5018 = 8'h38 == total_offset_15 ? field_byte_15 : _GEN_4858; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5019 = 8'h39 == total_offset_15 ? field_byte_15 : _GEN_4859; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5020 = 8'h3a == total_offset_15 ? field_byte_15 : _GEN_4860; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5021 = 8'h3b == total_offset_15 ? field_byte_15 : _GEN_4861; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5022 = 8'h3c == total_offset_15 ? field_byte_15 : _GEN_4862; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5023 = 8'h3d == total_offset_15 ? field_byte_15 : _GEN_4863; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5024 = 8'h3e == total_offset_15 ? field_byte_15 : _GEN_4864; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5025 = 8'h3f == total_offset_15 ? field_byte_15 : _GEN_4865; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5026 = 8'h40 == total_offset_15 ? field_byte_15 : _GEN_4866; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5027 = 8'h41 == total_offset_15 ? field_byte_15 : _GEN_4867; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5028 = 8'h42 == total_offset_15 ? field_byte_15 : _GEN_4868; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5029 = 8'h43 == total_offset_15 ? field_byte_15 : _GEN_4869; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5030 = 8'h44 == total_offset_15 ? field_byte_15 : _GEN_4870; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5031 = 8'h45 == total_offset_15 ? field_byte_15 : _GEN_4871; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5032 = 8'h46 == total_offset_15 ? field_byte_15 : _GEN_4872; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5033 = 8'h47 == total_offset_15 ? field_byte_15 : _GEN_4873; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5034 = 8'h48 == total_offset_15 ? field_byte_15 : _GEN_4874; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5035 = 8'h49 == total_offset_15 ? field_byte_15 : _GEN_4875; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5036 = 8'h4a == total_offset_15 ? field_byte_15 : _GEN_4876; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5037 = 8'h4b == total_offset_15 ? field_byte_15 : _GEN_4877; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5038 = 8'h4c == total_offset_15 ? field_byte_15 : _GEN_4878; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5039 = 8'h4d == total_offset_15 ? field_byte_15 : _GEN_4879; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5040 = 8'h4e == total_offset_15 ? field_byte_15 : _GEN_4880; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5041 = 8'h4f == total_offset_15 ? field_byte_15 : _GEN_4881; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5042 = 8'h50 == total_offset_15 ? field_byte_15 : _GEN_4882; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5043 = 8'h51 == total_offset_15 ? field_byte_15 : _GEN_4883; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5044 = 8'h52 == total_offset_15 ? field_byte_15 : _GEN_4884; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5045 = 8'h53 == total_offset_15 ? field_byte_15 : _GEN_4885; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5046 = 8'h54 == total_offset_15 ? field_byte_15 : _GEN_4886; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5047 = 8'h55 == total_offset_15 ? field_byte_15 : _GEN_4887; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5048 = 8'h56 == total_offset_15 ? field_byte_15 : _GEN_4888; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5049 = 8'h57 == total_offset_15 ? field_byte_15 : _GEN_4889; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5050 = 8'h58 == total_offset_15 ? field_byte_15 : _GEN_4890; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5051 = 8'h59 == total_offset_15 ? field_byte_15 : _GEN_4891; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5052 = 8'h5a == total_offset_15 ? field_byte_15 : _GEN_4892; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5053 = 8'h5b == total_offset_15 ? field_byte_15 : _GEN_4893; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5054 = 8'h5c == total_offset_15 ? field_byte_15 : _GEN_4894; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5055 = 8'h5d == total_offset_15 ? field_byte_15 : _GEN_4895; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5056 = 8'h5e == total_offset_15 ? field_byte_15 : _GEN_4896; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5057 = 8'h5f == total_offset_15 ? field_byte_15 : _GEN_4897; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5058 = 8'h60 == total_offset_15 ? field_byte_15 : _GEN_4898; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5059 = 8'h61 == total_offset_15 ? field_byte_15 : _GEN_4899; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5060 = 8'h62 == total_offset_15 ? field_byte_15 : _GEN_4900; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5061 = 8'h63 == total_offset_15 ? field_byte_15 : _GEN_4901; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5062 = 8'h64 == total_offset_15 ? field_byte_15 : _GEN_4902; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5063 = 8'h65 == total_offset_15 ? field_byte_15 : _GEN_4903; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5064 = 8'h66 == total_offset_15 ? field_byte_15 : _GEN_4904; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5065 = 8'h67 == total_offset_15 ? field_byte_15 : _GEN_4905; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5066 = 8'h68 == total_offset_15 ? field_byte_15 : _GEN_4906; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5067 = 8'h69 == total_offset_15 ? field_byte_15 : _GEN_4907; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5068 = 8'h6a == total_offset_15 ? field_byte_15 : _GEN_4908; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5069 = 8'h6b == total_offset_15 ? field_byte_15 : _GEN_4909; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5070 = 8'h6c == total_offset_15 ? field_byte_15 : _GEN_4910; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5071 = 8'h6d == total_offset_15 ? field_byte_15 : _GEN_4911; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5072 = 8'h6e == total_offset_15 ? field_byte_15 : _GEN_4912; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5073 = 8'h6f == total_offset_15 ? field_byte_15 : _GEN_4913; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5074 = 8'h70 == total_offset_15 ? field_byte_15 : _GEN_4914; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5075 = 8'h71 == total_offset_15 ? field_byte_15 : _GEN_4915; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5076 = 8'h72 == total_offset_15 ? field_byte_15 : _GEN_4916; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5077 = 8'h73 == total_offset_15 ? field_byte_15 : _GEN_4917; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5078 = 8'h74 == total_offset_15 ? field_byte_15 : _GEN_4918; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5079 = 8'h75 == total_offset_15 ? field_byte_15 : _GEN_4919; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5080 = 8'h76 == total_offset_15 ? field_byte_15 : _GEN_4920; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5081 = 8'h77 == total_offset_15 ? field_byte_15 : _GEN_4921; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5082 = 8'h78 == total_offset_15 ? field_byte_15 : _GEN_4922; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5083 = 8'h79 == total_offset_15 ? field_byte_15 : _GEN_4923; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5084 = 8'h7a == total_offset_15 ? field_byte_15 : _GEN_4924; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5085 = 8'h7b == total_offset_15 ? field_byte_15 : _GEN_4925; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5086 = 8'h7c == total_offset_15 ? field_byte_15 : _GEN_4926; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5087 = 8'h7d == total_offset_15 ? field_byte_15 : _GEN_4927; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5088 = 8'h7e == total_offset_15 ? field_byte_15 : _GEN_4928; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5089 = 8'h7f == total_offset_15 ? field_byte_15 : _GEN_4929; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5090 = 8'h80 == total_offset_15 ? field_byte_15 : _GEN_4930; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5091 = 8'h81 == total_offset_15 ? field_byte_15 : _GEN_4931; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5092 = 8'h82 == total_offset_15 ? field_byte_15 : _GEN_4932; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5093 = 8'h83 == total_offset_15 ? field_byte_15 : _GEN_4933; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5094 = 8'h84 == total_offset_15 ? field_byte_15 : _GEN_4934; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5095 = 8'h85 == total_offset_15 ? field_byte_15 : _GEN_4935; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5096 = 8'h86 == total_offset_15 ? field_byte_15 : _GEN_4936; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5097 = 8'h87 == total_offset_15 ? field_byte_15 : _GEN_4937; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5098 = 8'h88 == total_offset_15 ? field_byte_15 : _GEN_4938; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5099 = 8'h89 == total_offset_15 ? field_byte_15 : _GEN_4939; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5100 = 8'h8a == total_offset_15 ? field_byte_15 : _GEN_4940; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5101 = 8'h8b == total_offset_15 ? field_byte_15 : _GEN_4941; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5102 = 8'h8c == total_offset_15 ? field_byte_15 : _GEN_4942; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5103 = 8'h8d == total_offset_15 ? field_byte_15 : _GEN_4943; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5104 = 8'h8e == total_offset_15 ? field_byte_15 : _GEN_4944; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5105 = 8'h8f == total_offset_15 ? field_byte_15 : _GEN_4945; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5106 = 8'h90 == total_offset_15 ? field_byte_15 : _GEN_4946; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5107 = 8'h91 == total_offset_15 ? field_byte_15 : _GEN_4947; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5108 = 8'h92 == total_offset_15 ? field_byte_15 : _GEN_4948; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5109 = 8'h93 == total_offset_15 ? field_byte_15 : _GEN_4949; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5110 = 8'h94 == total_offset_15 ? field_byte_15 : _GEN_4950; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5111 = 8'h95 == total_offset_15 ? field_byte_15 : _GEN_4951; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5112 = 8'h96 == total_offset_15 ? field_byte_15 : _GEN_4952; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5113 = 8'h97 == total_offset_15 ? field_byte_15 : _GEN_4953; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5114 = 8'h98 == total_offset_15 ? field_byte_15 : _GEN_4954; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5115 = 8'h99 == total_offset_15 ? field_byte_15 : _GEN_4955; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5116 = 8'h9a == total_offset_15 ? field_byte_15 : _GEN_4956; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5117 = 8'h9b == total_offset_15 ? field_byte_15 : _GEN_4957; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5118 = 8'h9c == total_offset_15 ? field_byte_15 : _GEN_4958; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5119 = 8'h9d == total_offset_15 ? field_byte_15 : _GEN_4959; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5120 = 8'h9e == total_offset_15 ? field_byte_15 : _GEN_4960; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5121 = 8'h9f == total_offset_15 ? field_byte_15 : _GEN_4961; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5122 = 8'h7 < length_1 ? _GEN_4962 : _GEN_4802; // @[executor.scala 308:60]
  wire [7:0] _GEN_5123 = 8'h7 < length_1 ? _GEN_4963 : _GEN_4803; // @[executor.scala 308:60]
  wire [7:0] _GEN_5124 = 8'h7 < length_1 ? _GEN_4964 : _GEN_4804; // @[executor.scala 308:60]
  wire [7:0] _GEN_5125 = 8'h7 < length_1 ? _GEN_4965 : _GEN_4805; // @[executor.scala 308:60]
  wire [7:0] _GEN_5126 = 8'h7 < length_1 ? _GEN_4966 : _GEN_4806; // @[executor.scala 308:60]
  wire [7:0] _GEN_5127 = 8'h7 < length_1 ? _GEN_4967 : _GEN_4807; // @[executor.scala 308:60]
  wire [7:0] _GEN_5128 = 8'h7 < length_1 ? _GEN_4968 : _GEN_4808; // @[executor.scala 308:60]
  wire [7:0] _GEN_5129 = 8'h7 < length_1 ? _GEN_4969 : _GEN_4809; // @[executor.scala 308:60]
  wire [7:0] _GEN_5130 = 8'h7 < length_1 ? _GEN_4970 : _GEN_4810; // @[executor.scala 308:60]
  wire [7:0] _GEN_5131 = 8'h7 < length_1 ? _GEN_4971 : _GEN_4811; // @[executor.scala 308:60]
  wire [7:0] _GEN_5132 = 8'h7 < length_1 ? _GEN_4972 : _GEN_4812; // @[executor.scala 308:60]
  wire [7:0] _GEN_5133 = 8'h7 < length_1 ? _GEN_4973 : _GEN_4813; // @[executor.scala 308:60]
  wire [7:0] _GEN_5134 = 8'h7 < length_1 ? _GEN_4974 : _GEN_4814; // @[executor.scala 308:60]
  wire [7:0] _GEN_5135 = 8'h7 < length_1 ? _GEN_4975 : _GEN_4815; // @[executor.scala 308:60]
  wire [7:0] _GEN_5136 = 8'h7 < length_1 ? _GEN_4976 : _GEN_4816; // @[executor.scala 308:60]
  wire [7:0] _GEN_5137 = 8'h7 < length_1 ? _GEN_4977 : _GEN_4817; // @[executor.scala 308:60]
  wire [7:0] _GEN_5138 = 8'h7 < length_1 ? _GEN_4978 : _GEN_4818; // @[executor.scala 308:60]
  wire [7:0] _GEN_5139 = 8'h7 < length_1 ? _GEN_4979 : _GEN_4819; // @[executor.scala 308:60]
  wire [7:0] _GEN_5140 = 8'h7 < length_1 ? _GEN_4980 : _GEN_4820; // @[executor.scala 308:60]
  wire [7:0] _GEN_5141 = 8'h7 < length_1 ? _GEN_4981 : _GEN_4821; // @[executor.scala 308:60]
  wire [7:0] _GEN_5142 = 8'h7 < length_1 ? _GEN_4982 : _GEN_4822; // @[executor.scala 308:60]
  wire [7:0] _GEN_5143 = 8'h7 < length_1 ? _GEN_4983 : _GEN_4823; // @[executor.scala 308:60]
  wire [7:0] _GEN_5144 = 8'h7 < length_1 ? _GEN_4984 : _GEN_4824; // @[executor.scala 308:60]
  wire [7:0] _GEN_5145 = 8'h7 < length_1 ? _GEN_4985 : _GEN_4825; // @[executor.scala 308:60]
  wire [7:0] _GEN_5146 = 8'h7 < length_1 ? _GEN_4986 : _GEN_4826; // @[executor.scala 308:60]
  wire [7:0] _GEN_5147 = 8'h7 < length_1 ? _GEN_4987 : _GEN_4827; // @[executor.scala 308:60]
  wire [7:0] _GEN_5148 = 8'h7 < length_1 ? _GEN_4988 : _GEN_4828; // @[executor.scala 308:60]
  wire [7:0] _GEN_5149 = 8'h7 < length_1 ? _GEN_4989 : _GEN_4829; // @[executor.scala 308:60]
  wire [7:0] _GEN_5150 = 8'h7 < length_1 ? _GEN_4990 : _GEN_4830; // @[executor.scala 308:60]
  wire [7:0] _GEN_5151 = 8'h7 < length_1 ? _GEN_4991 : _GEN_4831; // @[executor.scala 308:60]
  wire [7:0] _GEN_5152 = 8'h7 < length_1 ? _GEN_4992 : _GEN_4832; // @[executor.scala 308:60]
  wire [7:0] _GEN_5153 = 8'h7 < length_1 ? _GEN_4993 : _GEN_4833; // @[executor.scala 308:60]
  wire [7:0] _GEN_5154 = 8'h7 < length_1 ? _GEN_4994 : _GEN_4834; // @[executor.scala 308:60]
  wire [7:0] _GEN_5155 = 8'h7 < length_1 ? _GEN_4995 : _GEN_4835; // @[executor.scala 308:60]
  wire [7:0] _GEN_5156 = 8'h7 < length_1 ? _GEN_4996 : _GEN_4836; // @[executor.scala 308:60]
  wire [7:0] _GEN_5157 = 8'h7 < length_1 ? _GEN_4997 : _GEN_4837; // @[executor.scala 308:60]
  wire [7:0] _GEN_5158 = 8'h7 < length_1 ? _GEN_4998 : _GEN_4838; // @[executor.scala 308:60]
  wire [7:0] _GEN_5159 = 8'h7 < length_1 ? _GEN_4999 : _GEN_4839; // @[executor.scala 308:60]
  wire [7:0] _GEN_5160 = 8'h7 < length_1 ? _GEN_5000 : _GEN_4840; // @[executor.scala 308:60]
  wire [7:0] _GEN_5161 = 8'h7 < length_1 ? _GEN_5001 : _GEN_4841; // @[executor.scala 308:60]
  wire [7:0] _GEN_5162 = 8'h7 < length_1 ? _GEN_5002 : _GEN_4842; // @[executor.scala 308:60]
  wire [7:0] _GEN_5163 = 8'h7 < length_1 ? _GEN_5003 : _GEN_4843; // @[executor.scala 308:60]
  wire [7:0] _GEN_5164 = 8'h7 < length_1 ? _GEN_5004 : _GEN_4844; // @[executor.scala 308:60]
  wire [7:0] _GEN_5165 = 8'h7 < length_1 ? _GEN_5005 : _GEN_4845; // @[executor.scala 308:60]
  wire [7:0] _GEN_5166 = 8'h7 < length_1 ? _GEN_5006 : _GEN_4846; // @[executor.scala 308:60]
  wire [7:0] _GEN_5167 = 8'h7 < length_1 ? _GEN_5007 : _GEN_4847; // @[executor.scala 308:60]
  wire [7:0] _GEN_5168 = 8'h7 < length_1 ? _GEN_5008 : _GEN_4848; // @[executor.scala 308:60]
  wire [7:0] _GEN_5169 = 8'h7 < length_1 ? _GEN_5009 : _GEN_4849; // @[executor.scala 308:60]
  wire [7:0] _GEN_5170 = 8'h7 < length_1 ? _GEN_5010 : _GEN_4850; // @[executor.scala 308:60]
  wire [7:0] _GEN_5171 = 8'h7 < length_1 ? _GEN_5011 : _GEN_4851; // @[executor.scala 308:60]
  wire [7:0] _GEN_5172 = 8'h7 < length_1 ? _GEN_5012 : _GEN_4852; // @[executor.scala 308:60]
  wire [7:0] _GEN_5173 = 8'h7 < length_1 ? _GEN_5013 : _GEN_4853; // @[executor.scala 308:60]
  wire [7:0] _GEN_5174 = 8'h7 < length_1 ? _GEN_5014 : _GEN_4854; // @[executor.scala 308:60]
  wire [7:0] _GEN_5175 = 8'h7 < length_1 ? _GEN_5015 : _GEN_4855; // @[executor.scala 308:60]
  wire [7:0] _GEN_5176 = 8'h7 < length_1 ? _GEN_5016 : _GEN_4856; // @[executor.scala 308:60]
  wire [7:0] _GEN_5177 = 8'h7 < length_1 ? _GEN_5017 : _GEN_4857; // @[executor.scala 308:60]
  wire [7:0] _GEN_5178 = 8'h7 < length_1 ? _GEN_5018 : _GEN_4858; // @[executor.scala 308:60]
  wire [7:0] _GEN_5179 = 8'h7 < length_1 ? _GEN_5019 : _GEN_4859; // @[executor.scala 308:60]
  wire [7:0] _GEN_5180 = 8'h7 < length_1 ? _GEN_5020 : _GEN_4860; // @[executor.scala 308:60]
  wire [7:0] _GEN_5181 = 8'h7 < length_1 ? _GEN_5021 : _GEN_4861; // @[executor.scala 308:60]
  wire [7:0] _GEN_5182 = 8'h7 < length_1 ? _GEN_5022 : _GEN_4862; // @[executor.scala 308:60]
  wire [7:0] _GEN_5183 = 8'h7 < length_1 ? _GEN_5023 : _GEN_4863; // @[executor.scala 308:60]
  wire [7:0] _GEN_5184 = 8'h7 < length_1 ? _GEN_5024 : _GEN_4864; // @[executor.scala 308:60]
  wire [7:0] _GEN_5185 = 8'h7 < length_1 ? _GEN_5025 : _GEN_4865; // @[executor.scala 308:60]
  wire [7:0] _GEN_5186 = 8'h7 < length_1 ? _GEN_5026 : _GEN_4866; // @[executor.scala 308:60]
  wire [7:0] _GEN_5187 = 8'h7 < length_1 ? _GEN_5027 : _GEN_4867; // @[executor.scala 308:60]
  wire [7:0] _GEN_5188 = 8'h7 < length_1 ? _GEN_5028 : _GEN_4868; // @[executor.scala 308:60]
  wire [7:0] _GEN_5189 = 8'h7 < length_1 ? _GEN_5029 : _GEN_4869; // @[executor.scala 308:60]
  wire [7:0] _GEN_5190 = 8'h7 < length_1 ? _GEN_5030 : _GEN_4870; // @[executor.scala 308:60]
  wire [7:0] _GEN_5191 = 8'h7 < length_1 ? _GEN_5031 : _GEN_4871; // @[executor.scala 308:60]
  wire [7:0] _GEN_5192 = 8'h7 < length_1 ? _GEN_5032 : _GEN_4872; // @[executor.scala 308:60]
  wire [7:0] _GEN_5193 = 8'h7 < length_1 ? _GEN_5033 : _GEN_4873; // @[executor.scala 308:60]
  wire [7:0] _GEN_5194 = 8'h7 < length_1 ? _GEN_5034 : _GEN_4874; // @[executor.scala 308:60]
  wire [7:0] _GEN_5195 = 8'h7 < length_1 ? _GEN_5035 : _GEN_4875; // @[executor.scala 308:60]
  wire [7:0] _GEN_5196 = 8'h7 < length_1 ? _GEN_5036 : _GEN_4876; // @[executor.scala 308:60]
  wire [7:0] _GEN_5197 = 8'h7 < length_1 ? _GEN_5037 : _GEN_4877; // @[executor.scala 308:60]
  wire [7:0] _GEN_5198 = 8'h7 < length_1 ? _GEN_5038 : _GEN_4878; // @[executor.scala 308:60]
  wire [7:0] _GEN_5199 = 8'h7 < length_1 ? _GEN_5039 : _GEN_4879; // @[executor.scala 308:60]
  wire [7:0] _GEN_5200 = 8'h7 < length_1 ? _GEN_5040 : _GEN_4880; // @[executor.scala 308:60]
  wire [7:0] _GEN_5201 = 8'h7 < length_1 ? _GEN_5041 : _GEN_4881; // @[executor.scala 308:60]
  wire [7:0] _GEN_5202 = 8'h7 < length_1 ? _GEN_5042 : _GEN_4882; // @[executor.scala 308:60]
  wire [7:0] _GEN_5203 = 8'h7 < length_1 ? _GEN_5043 : _GEN_4883; // @[executor.scala 308:60]
  wire [7:0] _GEN_5204 = 8'h7 < length_1 ? _GEN_5044 : _GEN_4884; // @[executor.scala 308:60]
  wire [7:0] _GEN_5205 = 8'h7 < length_1 ? _GEN_5045 : _GEN_4885; // @[executor.scala 308:60]
  wire [7:0] _GEN_5206 = 8'h7 < length_1 ? _GEN_5046 : _GEN_4886; // @[executor.scala 308:60]
  wire [7:0] _GEN_5207 = 8'h7 < length_1 ? _GEN_5047 : _GEN_4887; // @[executor.scala 308:60]
  wire [7:0] _GEN_5208 = 8'h7 < length_1 ? _GEN_5048 : _GEN_4888; // @[executor.scala 308:60]
  wire [7:0] _GEN_5209 = 8'h7 < length_1 ? _GEN_5049 : _GEN_4889; // @[executor.scala 308:60]
  wire [7:0] _GEN_5210 = 8'h7 < length_1 ? _GEN_5050 : _GEN_4890; // @[executor.scala 308:60]
  wire [7:0] _GEN_5211 = 8'h7 < length_1 ? _GEN_5051 : _GEN_4891; // @[executor.scala 308:60]
  wire [7:0] _GEN_5212 = 8'h7 < length_1 ? _GEN_5052 : _GEN_4892; // @[executor.scala 308:60]
  wire [7:0] _GEN_5213 = 8'h7 < length_1 ? _GEN_5053 : _GEN_4893; // @[executor.scala 308:60]
  wire [7:0] _GEN_5214 = 8'h7 < length_1 ? _GEN_5054 : _GEN_4894; // @[executor.scala 308:60]
  wire [7:0] _GEN_5215 = 8'h7 < length_1 ? _GEN_5055 : _GEN_4895; // @[executor.scala 308:60]
  wire [7:0] _GEN_5216 = 8'h7 < length_1 ? _GEN_5056 : _GEN_4896; // @[executor.scala 308:60]
  wire [7:0] _GEN_5217 = 8'h7 < length_1 ? _GEN_5057 : _GEN_4897; // @[executor.scala 308:60]
  wire [7:0] _GEN_5218 = 8'h7 < length_1 ? _GEN_5058 : _GEN_4898; // @[executor.scala 308:60]
  wire [7:0] _GEN_5219 = 8'h7 < length_1 ? _GEN_5059 : _GEN_4899; // @[executor.scala 308:60]
  wire [7:0] _GEN_5220 = 8'h7 < length_1 ? _GEN_5060 : _GEN_4900; // @[executor.scala 308:60]
  wire [7:0] _GEN_5221 = 8'h7 < length_1 ? _GEN_5061 : _GEN_4901; // @[executor.scala 308:60]
  wire [7:0] _GEN_5222 = 8'h7 < length_1 ? _GEN_5062 : _GEN_4902; // @[executor.scala 308:60]
  wire [7:0] _GEN_5223 = 8'h7 < length_1 ? _GEN_5063 : _GEN_4903; // @[executor.scala 308:60]
  wire [7:0] _GEN_5224 = 8'h7 < length_1 ? _GEN_5064 : _GEN_4904; // @[executor.scala 308:60]
  wire [7:0] _GEN_5225 = 8'h7 < length_1 ? _GEN_5065 : _GEN_4905; // @[executor.scala 308:60]
  wire [7:0] _GEN_5226 = 8'h7 < length_1 ? _GEN_5066 : _GEN_4906; // @[executor.scala 308:60]
  wire [7:0] _GEN_5227 = 8'h7 < length_1 ? _GEN_5067 : _GEN_4907; // @[executor.scala 308:60]
  wire [7:0] _GEN_5228 = 8'h7 < length_1 ? _GEN_5068 : _GEN_4908; // @[executor.scala 308:60]
  wire [7:0] _GEN_5229 = 8'h7 < length_1 ? _GEN_5069 : _GEN_4909; // @[executor.scala 308:60]
  wire [7:0] _GEN_5230 = 8'h7 < length_1 ? _GEN_5070 : _GEN_4910; // @[executor.scala 308:60]
  wire [7:0] _GEN_5231 = 8'h7 < length_1 ? _GEN_5071 : _GEN_4911; // @[executor.scala 308:60]
  wire [7:0] _GEN_5232 = 8'h7 < length_1 ? _GEN_5072 : _GEN_4912; // @[executor.scala 308:60]
  wire [7:0] _GEN_5233 = 8'h7 < length_1 ? _GEN_5073 : _GEN_4913; // @[executor.scala 308:60]
  wire [7:0] _GEN_5234 = 8'h7 < length_1 ? _GEN_5074 : _GEN_4914; // @[executor.scala 308:60]
  wire [7:0] _GEN_5235 = 8'h7 < length_1 ? _GEN_5075 : _GEN_4915; // @[executor.scala 308:60]
  wire [7:0] _GEN_5236 = 8'h7 < length_1 ? _GEN_5076 : _GEN_4916; // @[executor.scala 308:60]
  wire [7:0] _GEN_5237 = 8'h7 < length_1 ? _GEN_5077 : _GEN_4917; // @[executor.scala 308:60]
  wire [7:0] _GEN_5238 = 8'h7 < length_1 ? _GEN_5078 : _GEN_4918; // @[executor.scala 308:60]
  wire [7:0] _GEN_5239 = 8'h7 < length_1 ? _GEN_5079 : _GEN_4919; // @[executor.scala 308:60]
  wire [7:0] _GEN_5240 = 8'h7 < length_1 ? _GEN_5080 : _GEN_4920; // @[executor.scala 308:60]
  wire [7:0] _GEN_5241 = 8'h7 < length_1 ? _GEN_5081 : _GEN_4921; // @[executor.scala 308:60]
  wire [7:0] _GEN_5242 = 8'h7 < length_1 ? _GEN_5082 : _GEN_4922; // @[executor.scala 308:60]
  wire [7:0] _GEN_5243 = 8'h7 < length_1 ? _GEN_5083 : _GEN_4923; // @[executor.scala 308:60]
  wire [7:0] _GEN_5244 = 8'h7 < length_1 ? _GEN_5084 : _GEN_4924; // @[executor.scala 308:60]
  wire [7:0] _GEN_5245 = 8'h7 < length_1 ? _GEN_5085 : _GEN_4925; // @[executor.scala 308:60]
  wire [7:0] _GEN_5246 = 8'h7 < length_1 ? _GEN_5086 : _GEN_4926; // @[executor.scala 308:60]
  wire [7:0] _GEN_5247 = 8'h7 < length_1 ? _GEN_5087 : _GEN_4927; // @[executor.scala 308:60]
  wire [7:0] _GEN_5248 = 8'h7 < length_1 ? _GEN_5088 : _GEN_4928; // @[executor.scala 308:60]
  wire [7:0] _GEN_5249 = 8'h7 < length_1 ? _GEN_5089 : _GEN_4929; // @[executor.scala 308:60]
  wire [7:0] _GEN_5250 = 8'h7 < length_1 ? _GEN_5090 : _GEN_4930; // @[executor.scala 308:60]
  wire [7:0] _GEN_5251 = 8'h7 < length_1 ? _GEN_5091 : _GEN_4931; // @[executor.scala 308:60]
  wire [7:0] _GEN_5252 = 8'h7 < length_1 ? _GEN_5092 : _GEN_4932; // @[executor.scala 308:60]
  wire [7:0] _GEN_5253 = 8'h7 < length_1 ? _GEN_5093 : _GEN_4933; // @[executor.scala 308:60]
  wire [7:0] _GEN_5254 = 8'h7 < length_1 ? _GEN_5094 : _GEN_4934; // @[executor.scala 308:60]
  wire [7:0] _GEN_5255 = 8'h7 < length_1 ? _GEN_5095 : _GEN_4935; // @[executor.scala 308:60]
  wire [7:0] _GEN_5256 = 8'h7 < length_1 ? _GEN_5096 : _GEN_4936; // @[executor.scala 308:60]
  wire [7:0] _GEN_5257 = 8'h7 < length_1 ? _GEN_5097 : _GEN_4937; // @[executor.scala 308:60]
  wire [7:0] _GEN_5258 = 8'h7 < length_1 ? _GEN_5098 : _GEN_4938; // @[executor.scala 308:60]
  wire [7:0] _GEN_5259 = 8'h7 < length_1 ? _GEN_5099 : _GEN_4939; // @[executor.scala 308:60]
  wire [7:0] _GEN_5260 = 8'h7 < length_1 ? _GEN_5100 : _GEN_4940; // @[executor.scala 308:60]
  wire [7:0] _GEN_5261 = 8'h7 < length_1 ? _GEN_5101 : _GEN_4941; // @[executor.scala 308:60]
  wire [7:0] _GEN_5262 = 8'h7 < length_1 ? _GEN_5102 : _GEN_4942; // @[executor.scala 308:60]
  wire [7:0] _GEN_5263 = 8'h7 < length_1 ? _GEN_5103 : _GEN_4943; // @[executor.scala 308:60]
  wire [7:0] _GEN_5264 = 8'h7 < length_1 ? _GEN_5104 : _GEN_4944; // @[executor.scala 308:60]
  wire [7:0] _GEN_5265 = 8'h7 < length_1 ? _GEN_5105 : _GEN_4945; // @[executor.scala 308:60]
  wire [7:0] _GEN_5266 = 8'h7 < length_1 ? _GEN_5106 : _GEN_4946; // @[executor.scala 308:60]
  wire [7:0] _GEN_5267 = 8'h7 < length_1 ? _GEN_5107 : _GEN_4947; // @[executor.scala 308:60]
  wire [7:0] _GEN_5268 = 8'h7 < length_1 ? _GEN_5108 : _GEN_4948; // @[executor.scala 308:60]
  wire [7:0] _GEN_5269 = 8'h7 < length_1 ? _GEN_5109 : _GEN_4949; // @[executor.scala 308:60]
  wire [7:0] _GEN_5270 = 8'h7 < length_1 ? _GEN_5110 : _GEN_4950; // @[executor.scala 308:60]
  wire [7:0] _GEN_5271 = 8'h7 < length_1 ? _GEN_5111 : _GEN_4951; // @[executor.scala 308:60]
  wire [7:0] _GEN_5272 = 8'h7 < length_1 ? _GEN_5112 : _GEN_4952; // @[executor.scala 308:60]
  wire [7:0] _GEN_5273 = 8'h7 < length_1 ? _GEN_5113 : _GEN_4953; // @[executor.scala 308:60]
  wire [7:0] _GEN_5274 = 8'h7 < length_1 ? _GEN_5114 : _GEN_4954; // @[executor.scala 308:60]
  wire [7:0] _GEN_5275 = 8'h7 < length_1 ? _GEN_5115 : _GEN_4955; // @[executor.scala 308:60]
  wire [7:0] _GEN_5276 = 8'h7 < length_1 ? _GEN_5116 : _GEN_4956; // @[executor.scala 308:60]
  wire [7:0] _GEN_5277 = 8'h7 < length_1 ? _GEN_5117 : _GEN_4957; // @[executor.scala 308:60]
  wire [7:0] _GEN_5278 = 8'h7 < length_1 ? _GEN_5118 : _GEN_4958; // @[executor.scala 308:60]
  wire [7:0] _GEN_5279 = 8'h7 < length_1 ? _GEN_5119 : _GEN_4959; // @[executor.scala 308:60]
  wire [7:0] _GEN_5280 = 8'h7 < length_1 ? _GEN_5120 : _GEN_4960; // @[executor.scala 308:60]
  wire [7:0] _GEN_5281 = 8'h7 < length_1 ? _GEN_5121 : _GEN_4961; // @[executor.scala 308:60]
  wire [3:0] _GEN_5282 = length_1 == 8'h0 ? field_1[13:10] : _GEN_2560; // @[executor.scala 300:71 executor.scala 301:55]
  wire  _GEN_5283 = length_1 == 8'h0 ? field_1[0] : _GEN_2561; // @[executor.scala 300:71 executor.scala 302:55]
  wire [7:0] _GEN_5284 = length_1 == 8'h0 ? _GEN_2562 : _GEN_5122; // @[executor.scala 300:71]
  wire [7:0] _GEN_5285 = length_1 == 8'h0 ? _GEN_2563 : _GEN_5123; // @[executor.scala 300:71]
  wire [7:0] _GEN_5286 = length_1 == 8'h0 ? _GEN_2564 : _GEN_5124; // @[executor.scala 300:71]
  wire [7:0] _GEN_5287 = length_1 == 8'h0 ? _GEN_2565 : _GEN_5125; // @[executor.scala 300:71]
  wire [7:0] _GEN_5288 = length_1 == 8'h0 ? _GEN_2566 : _GEN_5126; // @[executor.scala 300:71]
  wire [7:0] _GEN_5289 = length_1 == 8'h0 ? _GEN_2567 : _GEN_5127; // @[executor.scala 300:71]
  wire [7:0] _GEN_5290 = length_1 == 8'h0 ? _GEN_2568 : _GEN_5128; // @[executor.scala 300:71]
  wire [7:0] _GEN_5291 = length_1 == 8'h0 ? _GEN_2569 : _GEN_5129; // @[executor.scala 300:71]
  wire [7:0] _GEN_5292 = length_1 == 8'h0 ? _GEN_2570 : _GEN_5130; // @[executor.scala 300:71]
  wire [7:0] _GEN_5293 = length_1 == 8'h0 ? _GEN_2571 : _GEN_5131; // @[executor.scala 300:71]
  wire [7:0] _GEN_5294 = length_1 == 8'h0 ? _GEN_2572 : _GEN_5132; // @[executor.scala 300:71]
  wire [7:0] _GEN_5295 = length_1 == 8'h0 ? _GEN_2573 : _GEN_5133; // @[executor.scala 300:71]
  wire [7:0] _GEN_5296 = length_1 == 8'h0 ? _GEN_2574 : _GEN_5134; // @[executor.scala 300:71]
  wire [7:0] _GEN_5297 = length_1 == 8'h0 ? _GEN_2575 : _GEN_5135; // @[executor.scala 300:71]
  wire [7:0] _GEN_5298 = length_1 == 8'h0 ? _GEN_2576 : _GEN_5136; // @[executor.scala 300:71]
  wire [7:0] _GEN_5299 = length_1 == 8'h0 ? _GEN_2577 : _GEN_5137; // @[executor.scala 300:71]
  wire [7:0] _GEN_5300 = length_1 == 8'h0 ? _GEN_2578 : _GEN_5138; // @[executor.scala 300:71]
  wire [7:0] _GEN_5301 = length_1 == 8'h0 ? _GEN_2579 : _GEN_5139; // @[executor.scala 300:71]
  wire [7:0] _GEN_5302 = length_1 == 8'h0 ? _GEN_2580 : _GEN_5140; // @[executor.scala 300:71]
  wire [7:0] _GEN_5303 = length_1 == 8'h0 ? _GEN_2581 : _GEN_5141; // @[executor.scala 300:71]
  wire [7:0] _GEN_5304 = length_1 == 8'h0 ? _GEN_2582 : _GEN_5142; // @[executor.scala 300:71]
  wire [7:0] _GEN_5305 = length_1 == 8'h0 ? _GEN_2583 : _GEN_5143; // @[executor.scala 300:71]
  wire [7:0] _GEN_5306 = length_1 == 8'h0 ? _GEN_2584 : _GEN_5144; // @[executor.scala 300:71]
  wire [7:0] _GEN_5307 = length_1 == 8'h0 ? _GEN_2585 : _GEN_5145; // @[executor.scala 300:71]
  wire [7:0] _GEN_5308 = length_1 == 8'h0 ? _GEN_2586 : _GEN_5146; // @[executor.scala 300:71]
  wire [7:0] _GEN_5309 = length_1 == 8'h0 ? _GEN_2587 : _GEN_5147; // @[executor.scala 300:71]
  wire [7:0] _GEN_5310 = length_1 == 8'h0 ? _GEN_2588 : _GEN_5148; // @[executor.scala 300:71]
  wire [7:0] _GEN_5311 = length_1 == 8'h0 ? _GEN_2589 : _GEN_5149; // @[executor.scala 300:71]
  wire [7:0] _GEN_5312 = length_1 == 8'h0 ? _GEN_2590 : _GEN_5150; // @[executor.scala 300:71]
  wire [7:0] _GEN_5313 = length_1 == 8'h0 ? _GEN_2591 : _GEN_5151; // @[executor.scala 300:71]
  wire [7:0] _GEN_5314 = length_1 == 8'h0 ? _GEN_2592 : _GEN_5152; // @[executor.scala 300:71]
  wire [7:0] _GEN_5315 = length_1 == 8'h0 ? _GEN_2593 : _GEN_5153; // @[executor.scala 300:71]
  wire [7:0] _GEN_5316 = length_1 == 8'h0 ? _GEN_2594 : _GEN_5154; // @[executor.scala 300:71]
  wire [7:0] _GEN_5317 = length_1 == 8'h0 ? _GEN_2595 : _GEN_5155; // @[executor.scala 300:71]
  wire [7:0] _GEN_5318 = length_1 == 8'h0 ? _GEN_2596 : _GEN_5156; // @[executor.scala 300:71]
  wire [7:0] _GEN_5319 = length_1 == 8'h0 ? _GEN_2597 : _GEN_5157; // @[executor.scala 300:71]
  wire [7:0] _GEN_5320 = length_1 == 8'h0 ? _GEN_2598 : _GEN_5158; // @[executor.scala 300:71]
  wire [7:0] _GEN_5321 = length_1 == 8'h0 ? _GEN_2599 : _GEN_5159; // @[executor.scala 300:71]
  wire [7:0] _GEN_5322 = length_1 == 8'h0 ? _GEN_2600 : _GEN_5160; // @[executor.scala 300:71]
  wire [7:0] _GEN_5323 = length_1 == 8'h0 ? _GEN_2601 : _GEN_5161; // @[executor.scala 300:71]
  wire [7:0] _GEN_5324 = length_1 == 8'h0 ? _GEN_2602 : _GEN_5162; // @[executor.scala 300:71]
  wire [7:0] _GEN_5325 = length_1 == 8'h0 ? _GEN_2603 : _GEN_5163; // @[executor.scala 300:71]
  wire [7:0] _GEN_5326 = length_1 == 8'h0 ? _GEN_2604 : _GEN_5164; // @[executor.scala 300:71]
  wire [7:0] _GEN_5327 = length_1 == 8'h0 ? _GEN_2605 : _GEN_5165; // @[executor.scala 300:71]
  wire [7:0] _GEN_5328 = length_1 == 8'h0 ? _GEN_2606 : _GEN_5166; // @[executor.scala 300:71]
  wire [7:0] _GEN_5329 = length_1 == 8'h0 ? _GEN_2607 : _GEN_5167; // @[executor.scala 300:71]
  wire [7:0] _GEN_5330 = length_1 == 8'h0 ? _GEN_2608 : _GEN_5168; // @[executor.scala 300:71]
  wire [7:0] _GEN_5331 = length_1 == 8'h0 ? _GEN_2609 : _GEN_5169; // @[executor.scala 300:71]
  wire [7:0] _GEN_5332 = length_1 == 8'h0 ? _GEN_2610 : _GEN_5170; // @[executor.scala 300:71]
  wire [7:0] _GEN_5333 = length_1 == 8'h0 ? _GEN_2611 : _GEN_5171; // @[executor.scala 300:71]
  wire [7:0] _GEN_5334 = length_1 == 8'h0 ? _GEN_2612 : _GEN_5172; // @[executor.scala 300:71]
  wire [7:0] _GEN_5335 = length_1 == 8'h0 ? _GEN_2613 : _GEN_5173; // @[executor.scala 300:71]
  wire [7:0] _GEN_5336 = length_1 == 8'h0 ? _GEN_2614 : _GEN_5174; // @[executor.scala 300:71]
  wire [7:0] _GEN_5337 = length_1 == 8'h0 ? _GEN_2615 : _GEN_5175; // @[executor.scala 300:71]
  wire [7:0] _GEN_5338 = length_1 == 8'h0 ? _GEN_2616 : _GEN_5176; // @[executor.scala 300:71]
  wire [7:0] _GEN_5339 = length_1 == 8'h0 ? _GEN_2617 : _GEN_5177; // @[executor.scala 300:71]
  wire [7:0] _GEN_5340 = length_1 == 8'h0 ? _GEN_2618 : _GEN_5178; // @[executor.scala 300:71]
  wire [7:0] _GEN_5341 = length_1 == 8'h0 ? _GEN_2619 : _GEN_5179; // @[executor.scala 300:71]
  wire [7:0] _GEN_5342 = length_1 == 8'h0 ? _GEN_2620 : _GEN_5180; // @[executor.scala 300:71]
  wire [7:0] _GEN_5343 = length_1 == 8'h0 ? _GEN_2621 : _GEN_5181; // @[executor.scala 300:71]
  wire [7:0] _GEN_5344 = length_1 == 8'h0 ? _GEN_2622 : _GEN_5182; // @[executor.scala 300:71]
  wire [7:0] _GEN_5345 = length_1 == 8'h0 ? _GEN_2623 : _GEN_5183; // @[executor.scala 300:71]
  wire [7:0] _GEN_5346 = length_1 == 8'h0 ? _GEN_2624 : _GEN_5184; // @[executor.scala 300:71]
  wire [7:0] _GEN_5347 = length_1 == 8'h0 ? _GEN_2625 : _GEN_5185; // @[executor.scala 300:71]
  wire [7:0] _GEN_5348 = length_1 == 8'h0 ? _GEN_2626 : _GEN_5186; // @[executor.scala 300:71]
  wire [7:0] _GEN_5349 = length_1 == 8'h0 ? _GEN_2627 : _GEN_5187; // @[executor.scala 300:71]
  wire [7:0] _GEN_5350 = length_1 == 8'h0 ? _GEN_2628 : _GEN_5188; // @[executor.scala 300:71]
  wire [7:0] _GEN_5351 = length_1 == 8'h0 ? _GEN_2629 : _GEN_5189; // @[executor.scala 300:71]
  wire [7:0] _GEN_5352 = length_1 == 8'h0 ? _GEN_2630 : _GEN_5190; // @[executor.scala 300:71]
  wire [7:0] _GEN_5353 = length_1 == 8'h0 ? _GEN_2631 : _GEN_5191; // @[executor.scala 300:71]
  wire [7:0] _GEN_5354 = length_1 == 8'h0 ? _GEN_2632 : _GEN_5192; // @[executor.scala 300:71]
  wire [7:0] _GEN_5355 = length_1 == 8'h0 ? _GEN_2633 : _GEN_5193; // @[executor.scala 300:71]
  wire [7:0] _GEN_5356 = length_1 == 8'h0 ? _GEN_2634 : _GEN_5194; // @[executor.scala 300:71]
  wire [7:0] _GEN_5357 = length_1 == 8'h0 ? _GEN_2635 : _GEN_5195; // @[executor.scala 300:71]
  wire [7:0] _GEN_5358 = length_1 == 8'h0 ? _GEN_2636 : _GEN_5196; // @[executor.scala 300:71]
  wire [7:0] _GEN_5359 = length_1 == 8'h0 ? _GEN_2637 : _GEN_5197; // @[executor.scala 300:71]
  wire [7:0] _GEN_5360 = length_1 == 8'h0 ? _GEN_2638 : _GEN_5198; // @[executor.scala 300:71]
  wire [7:0] _GEN_5361 = length_1 == 8'h0 ? _GEN_2639 : _GEN_5199; // @[executor.scala 300:71]
  wire [7:0] _GEN_5362 = length_1 == 8'h0 ? _GEN_2640 : _GEN_5200; // @[executor.scala 300:71]
  wire [7:0] _GEN_5363 = length_1 == 8'h0 ? _GEN_2641 : _GEN_5201; // @[executor.scala 300:71]
  wire [7:0] _GEN_5364 = length_1 == 8'h0 ? _GEN_2642 : _GEN_5202; // @[executor.scala 300:71]
  wire [7:0] _GEN_5365 = length_1 == 8'h0 ? _GEN_2643 : _GEN_5203; // @[executor.scala 300:71]
  wire [7:0] _GEN_5366 = length_1 == 8'h0 ? _GEN_2644 : _GEN_5204; // @[executor.scala 300:71]
  wire [7:0] _GEN_5367 = length_1 == 8'h0 ? _GEN_2645 : _GEN_5205; // @[executor.scala 300:71]
  wire [7:0] _GEN_5368 = length_1 == 8'h0 ? _GEN_2646 : _GEN_5206; // @[executor.scala 300:71]
  wire [7:0] _GEN_5369 = length_1 == 8'h0 ? _GEN_2647 : _GEN_5207; // @[executor.scala 300:71]
  wire [7:0] _GEN_5370 = length_1 == 8'h0 ? _GEN_2648 : _GEN_5208; // @[executor.scala 300:71]
  wire [7:0] _GEN_5371 = length_1 == 8'h0 ? _GEN_2649 : _GEN_5209; // @[executor.scala 300:71]
  wire [7:0] _GEN_5372 = length_1 == 8'h0 ? _GEN_2650 : _GEN_5210; // @[executor.scala 300:71]
  wire [7:0] _GEN_5373 = length_1 == 8'h0 ? _GEN_2651 : _GEN_5211; // @[executor.scala 300:71]
  wire [7:0] _GEN_5374 = length_1 == 8'h0 ? _GEN_2652 : _GEN_5212; // @[executor.scala 300:71]
  wire [7:0] _GEN_5375 = length_1 == 8'h0 ? _GEN_2653 : _GEN_5213; // @[executor.scala 300:71]
  wire [7:0] _GEN_5376 = length_1 == 8'h0 ? _GEN_2654 : _GEN_5214; // @[executor.scala 300:71]
  wire [7:0] _GEN_5377 = length_1 == 8'h0 ? _GEN_2655 : _GEN_5215; // @[executor.scala 300:71]
  wire [7:0] _GEN_5378 = length_1 == 8'h0 ? _GEN_2656 : _GEN_5216; // @[executor.scala 300:71]
  wire [7:0] _GEN_5379 = length_1 == 8'h0 ? _GEN_2657 : _GEN_5217; // @[executor.scala 300:71]
  wire [7:0] _GEN_5380 = length_1 == 8'h0 ? _GEN_2658 : _GEN_5218; // @[executor.scala 300:71]
  wire [7:0] _GEN_5381 = length_1 == 8'h0 ? _GEN_2659 : _GEN_5219; // @[executor.scala 300:71]
  wire [7:0] _GEN_5382 = length_1 == 8'h0 ? _GEN_2660 : _GEN_5220; // @[executor.scala 300:71]
  wire [7:0] _GEN_5383 = length_1 == 8'h0 ? _GEN_2661 : _GEN_5221; // @[executor.scala 300:71]
  wire [7:0] _GEN_5384 = length_1 == 8'h0 ? _GEN_2662 : _GEN_5222; // @[executor.scala 300:71]
  wire [7:0] _GEN_5385 = length_1 == 8'h0 ? _GEN_2663 : _GEN_5223; // @[executor.scala 300:71]
  wire [7:0] _GEN_5386 = length_1 == 8'h0 ? _GEN_2664 : _GEN_5224; // @[executor.scala 300:71]
  wire [7:0] _GEN_5387 = length_1 == 8'h0 ? _GEN_2665 : _GEN_5225; // @[executor.scala 300:71]
  wire [7:0] _GEN_5388 = length_1 == 8'h0 ? _GEN_2666 : _GEN_5226; // @[executor.scala 300:71]
  wire [7:0] _GEN_5389 = length_1 == 8'h0 ? _GEN_2667 : _GEN_5227; // @[executor.scala 300:71]
  wire [7:0] _GEN_5390 = length_1 == 8'h0 ? _GEN_2668 : _GEN_5228; // @[executor.scala 300:71]
  wire [7:0] _GEN_5391 = length_1 == 8'h0 ? _GEN_2669 : _GEN_5229; // @[executor.scala 300:71]
  wire [7:0] _GEN_5392 = length_1 == 8'h0 ? _GEN_2670 : _GEN_5230; // @[executor.scala 300:71]
  wire [7:0] _GEN_5393 = length_1 == 8'h0 ? _GEN_2671 : _GEN_5231; // @[executor.scala 300:71]
  wire [7:0] _GEN_5394 = length_1 == 8'h0 ? _GEN_2672 : _GEN_5232; // @[executor.scala 300:71]
  wire [7:0] _GEN_5395 = length_1 == 8'h0 ? _GEN_2673 : _GEN_5233; // @[executor.scala 300:71]
  wire [7:0] _GEN_5396 = length_1 == 8'h0 ? _GEN_2674 : _GEN_5234; // @[executor.scala 300:71]
  wire [7:0] _GEN_5397 = length_1 == 8'h0 ? _GEN_2675 : _GEN_5235; // @[executor.scala 300:71]
  wire [7:0] _GEN_5398 = length_1 == 8'h0 ? _GEN_2676 : _GEN_5236; // @[executor.scala 300:71]
  wire [7:0] _GEN_5399 = length_1 == 8'h0 ? _GEN_2677 : _GEN_5237; // @[executor.scala 300:71]
  wire [7:0] _GEN_5400 = length_1 == 8'h0 ? _GEN_2678 : _GEN_5238; // @[executor.scala 300:71]
  wire [7:0] _GEN_5401 = length_1 == 8'h0 ? _GEN_2679 : _GEN_5239; // @[executor.scala 300:71]
  wire [7:0] _GEN_5402 = length_1 == 8'h0 ? _GEN_2680 : _GEN_5240; // @[executor.scala 300:71]
  wire [7:0] _GEN_5403 = length_1 == 8'h0 ? _GEN_2681 : _GEN_5241; // @[executor.scala 300:71]
  wire [7:0] _GEN_5404 = length_1 == 8'h0 ? _GEN_2682 : _GEN_5242; // @[executor.scala 300:71]
  wire [7:0] _GEN_5405 = length_1 == 8'h0 ? _GEN_2683 : _GEN_5243; // @[executor.scala 300:71]
  wire [7:0] _GEN_5406 = length_1 == 8'h0 ? _GEN_2684 : _GEN_5244; // @[executor.scala 300:71]
  wire [7:0] _GEN_5407 = length_1 == 8'h0 ? _GEN_2685 : _GEN_5245; // @[executor.scala 300:71]
  wire [7:0] _GEN_5408 = length_1 == 8'h0 ? _GEN_2686 : _GEN_5246; // @[executor.scala 300:71]
  wire [7:0] _GEN_5409 = length_1 == 8'h0 ? _GEN_2687 : _GEN_5247; // @[executor.scala 300:71]
  wire [7:0] _GEN_5410 = length_1 == 8'h0 ? _GEN_2688 : _GEN_5248; // @[executor.scala 300:71]
  wire [7:0] _GEN_5411 = length_1 == 8'h0 ? _GEN_2689 : _GEN_5249; // @[executor.scala 300:71]
  wire [7:0] _GEN_5412 = length_1 == 8'h0 ? _GEN_2690 : _GEN_5250; // @[executor.scala 300:71]
  wire [7:0] _GEN_5413 = length_1 == 8'h0 ? _GEN_2691 : _GEN_5251; // @[executor.scala 300:71]
  wire [7:0] _GEN_5414 = length_1 == 8'h0 ? _GEN_2692 : _GEN_5252; // @[executor.scala 300:71]
  wire [7:0] _GEN_5415 = length_1 == 8'h0 ? _GEN_2693 : _GEN_5253; // @[executor.scala 300:71]
  wire [7:0] _GEN_5416 = length_1 == 8'h0 ? _GEN_2694 : _GEN_5254; // @[executor.scala 300:71]
  wire [7:0] _GEN_5417 = length_1 == 8'h0 ? _GEN_2695 : _GEN_5255; // @[executor.scala 300:71]
  wire [7:0] _GEN_5418 = length_1 == 8'h0 ? _GEN_2696 : _GEN_5256; // @[executor.scala 300:71]
  wire [7:0] _GEN_5419 = length_1 == 8'h0 ? _GEN_2697 : _GEN_5257; // @[executor.scala 300:71]
  wire [7:0] _GEN_5420 = length_1 == 8'h0 ? _GEN_2698 : _GEN_5258; // @[executor.scala 300:71]
  wire [7:0] _GEN_5421 = length_1 == 8'h0 ? _GEN_2699 : _GEN_5259; // @[executor.scala 300:71]
  wire [7:0] _GEN_5422 = length_1 == 8'h0 ? _GEN_2700 : _GEN_5260; // @[executor.scala 300:71]
  wire [7:0] _GEN_5423 = length_1 == 8'h0 ? _GEN_2701 : _GEN_5261; // @[executor.scala 300:71]
  wire [7:0] _GEN_5424 = length_1 == 8'h0 ? _GEN_2702 : _GEN_5262; // @[executor.scala 300:71]
  wire [7:0] _GEN_5425 = length_1 == 8'h0 ? _GEN_2703 : _GEN_5263; // @[executor.scala 300:71]
  wire [7:0] _GEN_5426 = length_1 == 8'h0 ? _GEN_2704 : _GEN_5264; // @[executor.scala 300:71]
  wire [7:0] _GEN_5427 = length_1 == 8'h0 ? _GEN_2705 : _GEN_5265; // @[executor.scala 300:71]
  wire [7:0] _GEN_5428 = length_1 == 8'h0 ? _GEN_2706 : _GEN_5266; // @[executor.scala 300:71]
  wire [7:0] _GEN_5429 = length_1 == 8'h0 ? _GEN_2707 : _GEN_5267; // @[executor.scala 300:71]
  wire [7:0] _GEN_5430 = length_1 == 8'h0 ? _GEN_2708 : _GEN_5268; // @[executor.scala 300:71]
  wire [7:0] _GEN_5431 = length_1 == 8'h0 ? _GEN_2709 : _GEN_5269; // @[executor.scala 300:71]
  wire [7:0] _GEN_5432 = length_1 == 8'h0 ? _GEN_2710 : _GEN_5270; // @[executor.scala 300:71]
  wire [7:0] _GEN_5433 = length_1 == 8'h0 ? _GEN_2711 : _GEN_5271; // @[executor.scala 300:71]
  wire [7:0] _GEN_5434 = length_1 == 8'h0 ? _GEN_2712 : _GEN_5272; // @[executor.scala 300:71]
  wire [7:0] _GEN_5435 = length_1 == 8'h0 ? _GEN_2713 : _GEN_5273; // @[executor.scala 300:71]
  wire [7:0] _GEN_5436 = length_1 == 8'h0 ? _GEN_2714 : _GEN_5274; // @[executor.scala 300:71]
  wire [7:0] _GEN_5437 = length_1 == 8'h0 ? _GEN_2715 : _GEN_5275; // @[executor.scala 300:71]
  wire [7:0] _GEN_5438 = length_1 == 8'h0 ? _GEN_2716 : _GEN_5276; // @[executor.scala 300:71]
  wire [7:0] _GEN_5439 = length_1 == 8'h0 ? _GEN_2717 : _GEN_5277; // @[executor.scala 300:71]
  wire [7:0] _GEN_5440 = length_1 == 8'h0 ? _GEN_2718 : _GEN_5278; // @[executor.scala 300:71]
  wire [7:0] _GEN_5441 = length_1 == 8'h0 ? _GEN_2719 : _GEN_5279; // @[executor.scala 300:71]
  wire [7:0] _GEN_5442 = length_1 == 8'h0 ? _GEN_2720 : _GEN_5280; // @[executor.scala 300:71]
  wire [7:0] _GEN_5443 = length_1 == 8'h0 ? _GEN_2721 : _GEN_5281; // @[executor.scala 300:71]
  wire [7:0] field_byte_16 = field_2[63:56]; // @[executor.scala 305:57]
  wire [8:0] _total_offset_T_16 = {{1'd0}, offset_2}; // @[executor.scala 307:57]
  wire [7:0] total_offset_16 = _total_offset_T_16[7:0]; // @[executor.scala 307:57]
  wire [7:0] _GEN_5444 = 8'h0 == total_offset_16 ? field_byte_16 : _GEN_5284; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5445 = 8'h1 == total_offset_16 ? field_byte_16 : _GEN_5285; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5446 = 8'h2 == total_offset_16 ? field_byte_16 : _GEN_5286; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5447 = 8'h3 == total_offset_16 ? field_byte_16 : _GEN_5287; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5448 = 8'h4 == total_offset_16 ? field_byte_16 : _GEN_5288; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5449 = 8'h5 == total_offset_16 ? field_byte_16 : _GEN_5289; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5450 = 8'h6 == total_offset_16 ? field_byte_16 : _GEN_5290; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5451 = 8'h7 == total_offset_16 ? field_byte_16 : _GEN_5291; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5452 = 8'h8 == total_offset_16 ? field_byte_16 : _GEN_5292; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5453 = 8'h9 == total_offset_16 ? field_byte_16 : _GEN_5293; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5454 = 8'ha == total_offset_16 ? field_byte_16 : _GEN_5294; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5455 = 8'hb == total_offset_16 ? field_byte_16 : _GEN_5295; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5456 = 8'hc == total_offset_16 ? field_byte_16 : _GEN_5296; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5457 = 8'hd == total_offset_16 ? field_byte_16 : _GEN_5297; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5458 = 8'he == total_offset_16 ? field_byte_16 : _GEN_5298; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5459 = 8'hf == total_offset_16 ? field_byte_16 : _GEN_5299; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5460 = 8'h10 == total_offset_16 ? field_byte_16 : _GEN_5300; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5461 = 8'h11 == total_offset_16 ? field_byte_16 : _GEN_5301; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5462 = 8'h12 == total_offset_16 ? field_byte_16 : _GEN_5302; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5463 = 8'h13 == total_offset_16 ? field_byte_16 : _GEN_5303; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5464 = 8'h14 == total_offset_16 ? field_byte_16 : _GEN_5304; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5465 = 8'h15 == total_offset_16 ? field_byte_16 : _GEN_5305; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5466 = 8'h16 == total_offset_16 ? field_byte_16 : _GEN_5306; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5467 = 8'h17 == total_offset_16 ? field_byte_16 : _GEN_5307; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5468 = 8'h18 == total_offset_16 ? field_byte_16 : _GEN_5308; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5469 = 8'h19 == total_offset_16 ? field_byte_16 : _GEN_5309; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5470 = 8'h1a == total_offset_16 ? field_byte_16 : _GEN_5310; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5471 = 8'h1b == total_offset_16 ? field_byte_16 : _GEN_5311; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5472 = 8'h1c == total_offset_16 ? field_byte_16 : _GEN_5312; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5473 = 8'h1d == total_offset_16 ? field_byte_16 : _GEN_5313; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5474 = 8'h1e == total_offset_16 ? field_byte_16 : _GEN_5314; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5475 = 8'h1f == total_offset_16 ? field_byte_16 : _GEN_5315; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5476 = 8'h20 == total_offset_16 ? field_byte_16 : _GEN_5316; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5477 = 8'h21 == total_offset_16 ? field_byte_16 : _GEN_5317; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5478 = 8'h22 == total_offset_16 ? field_byte_16 : _GEN_5318; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5479 = 8'h23 == total_offset_16 ? field_byte_16 : _GEN_5319; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5480 = 8'h24 == total_offset_16 ? field_byte_16 : _GEN_5320; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5481 = 8'h25 == total_offset_16 ? field_byte_16 : _GEN_5321; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5482 = 8'h26 == total_offset_16 ? field_byte_16 : _GEN_5322; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5483 = 8'h27 == total_offset_16 ? field_byte_16 : _GEN_5323; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5484 = 8'h28 == total_offset_16 ? field_byte_16 : _GEN_5324; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5485 = 8'h29 == total_offset_16 ? field_byte_16 : _GEN_5325; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5486 = 8'h2a == total_offset_16 ? field_byte_16 : _GEN_5326; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5487 = 8'h2b == total_offset_16 ? field_byte_16 : _GEN_5327; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5488 = 8'h2c == total_offset_16 ? field_byte_16 : _GEN_5328; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5489 = 8'h2d == total_offset_16 ? field_byte_16 : _GEN_5329; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5490 = 8'h2e == total_offset_16 ? field_byte_16 : _GEN_5330; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5491 = 8'h2f == total_offset_16 ? field_byte_16 : _GEN_5331; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5492 = 8'h30 == total_offset_16 ? field_byte_16 : _GEN_5332; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5493 = 8'h31 == total_offset_16 ? field_byte_16 : _GEN_5333; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5494 = 8'h32 == total_offset_16 ? field_byte_16 : _GEN_5334; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5495 = 8'h33 == total_offset_16 ? field_byte_16 : _GEN_5335; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5496 = 8'h34 == total_offset_16 ? field_byte_16 : _GEN_5336; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5497 = 8'h35 == total_offset_16 ? field_byte_16 : _GEN_5337; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5498 = 8'h36 == total_offset_16 ? field_byte_16 : _GEN_5338; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5499 = 8'h37 == total_offset_16 ? field_byte_16 : _GEN_5339; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5500 = 8'h38 == total_offset_16 ? field_byte_16 : _GEN_5340; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5501 = 8'h39 == total_offset_16 ? field_byte_16 : _GEN_5341; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5502 = 8'h3a == total_offset_16 ? field_byte_16 : _GEN_5342; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5503 = 8'h3b == total_offset_16 ? field_byte_16 : _GEN_5343; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5504 = 8'h3c == total_offset_16 ? field_byte_16 : _GEN_5344; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5505 = 8'h3d == total_offset_16 ? field_byte_16 : _GEN_5345; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5506 = 8'h3e == total_offset_16 ? field_byte_16 : _GEN_5346; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5507 = 8'h3f == total_offset_16 ? field_byte_16 : _GEN_5347; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5508 = 8'h40 == total_offset_16 ? field_byte_16 : _GEN_5348; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5509 = 8'h41 == total_offset_16 ? field_byte_16 : _GEN_5349; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5510 = 8'h42 == total_offset_16 ? field_byte_16 : _GEN_5350; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5511 = 8'h43 == total_offset_16 ? field_byte_16 : _GEN_5351; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5512 = 8'h44 == total_offset_16 ? field_byte_16 : _GEN_5352; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5513 = 8'h45 == total_offset_16 ? field_byte_16 : _GEN_5353; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5514 = 8'h46 == total_offset_16 ? field_byte_16 : _GEN_5354; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5515 = 8'h47 == total_offset_16 ? field_byte_16 : _GEN_5355; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5516 = 8'h48 == total_offset_16 ? field_byte_16 : _GEN_5356; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5517 = 8'h49 == total_offset_16 ? field_byte_16 : _GEN_5357; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5518 = 8'h4a == total_offset_16 ? field_byte_16 : _GEN_5358; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5519 = 8'h4b == total_offset_16 ? field_byte_16 : _GEN_5359; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5520 = 8'h4c == total_offset_16 ? field_byte_16 : _GEN_5360; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5521 = 8'h4d == total_offset_16 ? field_byte_16 : _GEN_5361; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5522 = 8'h4e == total_offset_16 ? field_byte_16 : _GEN_5362; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5523 = 8'h4f == total_offset_16 ? field_byte_16 : _GEN_5363; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5524 = 8'h50 == total_offset_16 ? field_byte_16 : _GEN_5364; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5525 = 8'h51 == total_offset_16 ? field_byte_16 : _GEN_5365; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5526 = 8'h52 == total_offset_16 ? field_byte_16 : _GEN_5366; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5527 = 8'h53 == total_offset_16 ? field_byte_16 : _GEN_5367; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5528 = 8'h54 == total_offset_16 ? field_byte_16 : _GEN_5368; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5529 = 8'h55 == total_offset_16 ? field_byte_16 : _GEN_5369; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5530 = 8'h56 == total_offset_16 ? field_byte_16 : _GEN_5370; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5531 = 8'h57 == total_offset_16 ? field_byte_16 : _GEN_5371; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5532 = 8'h58 == total_offset_16 ? field_byte_16 : _GEN_5372; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5533 = 8'h59 == total_offset_16 ? field_byte_16 : _GEN_5373; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5534 = 8'h5a == total_offset_16 ? field_byte_16 : _GEN_5374; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5535 = 8'h5b == total_offset_16 ? field_byte_16 : _GEN_5375; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5536 = 8'h5c == total_offset_16 ? field_byte_16 : _GEN_5376; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5537 = 8'h5d == total_offset_16 ? field_byte_16 : _GEN_5377; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5538 = 8'h5e == total_offset_16 ? field_byte_16 : _GEN_5378; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5539 = 8'h5f == total_offset_16 ? field_byte_16 : _GEN_5379; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5540 = 8'h60 == total_offset_16 ? field_byte_16 : _GEN_5380; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5541 = 8'h61 == total_offset_16 ? field_byte_16 : _GEN_5381; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5542 = 8'h62 == total_offset_16 ? field_byte_16 : _GEN_5382; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5543 = 8'h63 == total_offset_16 ? field_byte_16 : _GEN_5383; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5544 = 8'h64 == total_offset_16 ? field_byte_16 : _GEN_5384; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5545 = 8'h65 == total_offset_16 ? field_byte_16 : _GEN_5385; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5546 = 8'h66 == total_offset_16 ? field_byte_16 : _GEN_5386; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5547 = 8'h67 == total_offset_16 ? field_byte_16 : _GEN_5387; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5548 = 8'h68 == total_offset_16 ? field_byte_16 : _GEN_5388; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5549 = 8'h69 == total_offset_16 ? field_byte_16 : _GEN_5389; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5550 = 8'h6a == total_offset_16 ? field_byte_16 : _GEN_5390; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5551 = 8'h6b == total_offset_16 ? field_byte_16 : _GEN_5391; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5552 = 8'h6c == total_offset_16 ? field_byte_16 : _GEN_5392; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5553 = 8'h6d == total_offset_16 ? field_byte_16 : _GEN_5393; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5554 = 8'h6e == total_offset_16 ? field_byte_16 : _GEN_5394; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5555 = 8'h6f == total_offset_16 ? field_byte_16 : _GEN_5395; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5556 = 8'h70 == total_offset_16 ? field_byte_16 : _GEN_5396; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5557 = 8'h71 == total_offset_16 ? field_byte_16 : _GEN_5397; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5558 = 8'h72 == total_offset_16 ? field_byte_16 : _GEN_5398; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5559 = 8'h73 == total_offset_16 ? field_byte_16 : _GEN_5399; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5560 = 8'h74 == total_offset_16 ? field_byte_16 : _GEN_5400; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5561 = 8'h75 == total_offset_16 ? field_byte_16 : _GEN_5401; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5562 = 8'h76 == total_offset_16 ? field_byte_16 : _GEN_5402; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5563 = 8'h77 == total_offset_16 ? field_byte_16 : _GEN_5403; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5564 = 8'h78 == total_offset_16 ? field_byte_16 : _GEN_5404; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5565 = 8'h79 == total_offset_16 ? field_byte_16 : _GEN_5405; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5566 = 8'h7a == total_offset_16 ? field_byte_16 : _GEN_5406; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5567 = 8'h7b == total_offset_16 ? field_byte_16 : _GEN_5407; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5568 = 8'h7c == total_offset_16 ? field_byte_16 : _GEN_5408; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5569 = 8'h7d == total_offset_16 ? field_byte_16 : _GEN_5409; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5570 = 8'h7e == total_offset_16 ? field_byte_16 : _GEN_5410; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5571 = 8'h7f == total_offset_16 ? field_byte_16 : _GEN_5411; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5572 = 8'h80 == total_offset_16 ? field_byte_16 : _GEN_5412; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5573 = 8'h81 == total_offset_16 ? field_byte_16 : _GEN_5413; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5574 = 8'h82 == total_offset_16 ? field_byte_16 : _GEN_5414; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5575 = 8'h83 == total_offset_16 ? field_byte_16 : _GEN_5415; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5576 = 8'h84 == total_offset_16 ? field_byte_16 : _GEN_5416; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5577 = 8'h85 == total_offset_16 ? field_byte_16 : _GEN_5417; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5578 = 8'h86 == total_offset_16 ? field_byte_16 : _GEN_5418; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5579 = 8'h87 == total_offset_16 ? field_byte_16 : _GEN_5419; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5580 = 8'h88 == total_offset_16 ? field_byte_16 : _GEN_5420; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5581 = 8'h89 == total_offset_16 ? field_byte_16 : _GEN_5421; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5582 = 8'h8a == total_offset_16 ? field_byte_16 : _GEN_5422; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5583 = 8'h8b == total_offset_16 ? field_byte_16 : _GEN_5423; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5584 = 8'h8c == total_offset_16 ? field_byte_16 : _GEN_5424; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5585 = 8'h8d == total_offset_16 ? field_byte_16 : _GEN_5425; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5586 = 8'h8e == total_offset_16 ? field_byte_16 : _GEN_5426; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5587 = 8'h8f == total_offset_16 ? field_byte_16 : _GEN_5427; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5588 = 8'h90 == total_offset_16 ? field_byte_16 : _GEN_5428; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5589 = 8'h91 == total_offset_16 ? field_byte_16 : _GEN_5429; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5590 = 8'h92 == total_offset_16 ? field_byte_16 : _GEN_5430; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5591 = 8'h93 == total_offset_16 ? field_byte_16 : _GEN_5431; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5592 = 8'h94 == total_offset_16 ? field_byte_16 : _GEN_5432; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5593 = 8'h95 == total_offset_16 ? field_byte_16 : _GEN_5433; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5594 = 8'h96 == total_offset_16 ? field_byte_16 : _GEN_5434; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5595 = 8'h97 == total_offset_16 ? field_byte_16 : _GEN_5435; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5596 = 8'h98 == total_offset_16 ? field_byte_16 : _GEN_5436; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5597 = 8'h99 == total_offset_16 ? field_byte_16 : _GEN_5437; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5598 = 8'h9a == total_offset_16 ? field_byte_16 : _GEN_5438; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5599 = 8'h9b == total_offset_16 ? field_byte_16 : _GEN_5439; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5600 = 8'h9c == total_offset_16 ? field_byte_16 : _GEN_5440; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5601 = 8'h9d == total_offset_16 ? field_byte_16 : _GEN_5441; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5602 = 8'h9e == total_offset_16 ? field_byte_16 : _GEN_5442; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5603 = 8'h9f == total_offset_16 ? field_byte_16 : _GEN_5443; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5604 = 8'h0 < length_2 ? _GEN_5444 : _GEN_5284; // @[executor.scala 308:60]
  wire [7:0] _GEN_5605 = 8'h0 < length_2 ? _GEN_5445 : _GEN_5285; // @[executor.scala 308:60]
  wire [7:0] _GEN_5606 = 8'h0 < length_2 ? _GEN_5446 : _GEN_5286; // @[executor.scala 308:60]
  wire [7:0] _GEN_5607 = 8'h0 < length_2 ? _GEN_5447 : _GEN_5287; // @[executor.scala 308:60]
  wire [7:0] _GEN_5608 = 8'h0 < length_2 ? _GEN_5448 : _GEN_5288; // @[executor.scala 308:60]
  wire [7:0] _GEN_5609 = 8'h0 < length_2 ? _GEN_5449 : _GEN_5289; // @[executor.scala 308:60]
  wire [7:0] _GEN_5610 = 8'h0 < length_2 ? _GEN_5450 : _GEN_5290; // @[executor.scala 308:60]
  wire [7:0] _GEN_5611 = 8'h0 < length_2 ? _GEN_5451 : _GEN_5291; // @[executor.scala 308:60]
  wire [7:0] _GEN_5612 = 8'h0 < length_2 ? _GEN_5452 : _GEN_5292; // @[executor.scala 308:60]
  wire [7:0] _GEN_5613 = 8'h0 < length_2 ? _GEN_5453 : _GEN_5293; // @[executor.scala 308:60]
  wire [7:0] _GEN_5614 = 8'h0 < length_2 ? _GEN_5454 : _GEN_5294; // @[executor.scala 308:60]
  wire [7:0] _GEN_5615 = 8'h0 < length_2 ? _GEN_5455 : _GEN_5295; // @[executor.scala 308:60]
  wire [7:0] _GEN_5616 = 8'h0 < length_2 ? _GEN_5456 : _GEN_5296; // @[executor.scala 308:60]
  wire [7:0] _GEN_5617 = 8'h0 < length_2 ? _GEN_5457 : _GEN_5297; // @[executor.scala 308:60]
  wire [7:0] _GEN_5618 = 8'h0 < length_2 ? _GEN_5458 : _GEN_5298; // @[executor.scala 308:60]
  wire [7:0] _GEN_5619 = 8'h0 < length_2 ? _GEN_5459 : _GEN_5299; // @[executor.scala 308:60]
  wire [7:0] _GEN_5620 = 8'h0 < length_2 ? _GEN_5460 : _GEN_5300; // @[executor.scala 308:60]
  wire [7:0] _GEN_5621 = 8'h0 < length_2 ? _GEN_5461 : _GEN_5301; // @[executor.scala 308:60]
  wire [7:0] _GEN_5622 = 8'h0 < length_2 ? _GEN_5462 : _GEN_5302; // @[executor.scala 308:60]
  wire [7:0] _GEN_5623 = 8'h0 < length_2 ? _GEN_5463 : _GEN_5303; // @[executor.scala 308:60]
  wire [7:0] _GEN_5624 = 8'h0 < length_2 ? _GEN_5464 : _GEN_5304; // @[executor.scala 308:60]
  wire [7:0] _GEN_5625 = 8'h0 < length_2 ? _GEN_5465 : _GEN_5305; // @[executor.scala 308:60]
  wire [7:0] _GEN_5626 = 8'h0 < length_2 ? _GEN_5466 : _GEN_5306; // @[executor.scala 308:60]
  wire [7:0] _GEN_5627 = 8'h0 < length_2 ? _GEN_5467 : _GEN_5307; // @[executor.scala 308:60]
  wire [7:0] _GEN_5628 = 8'h0 < length_2 ? _GEN_5468 : _GEN_5308; // @[executor.scala 308:60]
  wire [7:0] _GEN_5629 = 8'h0 < length_2 ? _GEN_5469 : _GEN_5309; // @[executor.scala 308:60]
  wire [7:0] _GEN_5630 = 8'h0 < length_2 ? _GEN_5470 : _GEN_5310; // @[executor.scala 308:60]
  wire [7:0] _GEN_5631 = 8'h0 < length_2 ? _GEN_5471 : _GEN_5311; // @[executor.scala 308:60]
  wire [7:0] _GEN_5632 = 8'h0 < length_2 ? _GEN_5472 : _GEN_5312; // @[executor.scala 308:60]
  wire [7:0] _GEN_5633 = 8'h0 < length_2 ? _GEN_5473 : _GEN_5313; // @[executor.scala 308:60]
  wire [7:0] _GEN_5634 = 8'h0 < length_2 ? _GEN_5474 : _GEN_5314; // @[executor.scala 308:60]
  wire [7:0] _GEN_5635 = 8'h0 < length_2 ? _GEN_5475 : _GEN_5315; // @[executor.scala 308:60]
  wire [7:0] _GEN_5636 = 8'h0 < length_2 ? _GEN_5476 : _GEN_5316; // @[executor.scala 308:60]
  wire [7:0] _GEN_5637 = 8'h0 < length_2 ? _GEN_5477 : _GEN_5317; // @[executor.scala 308:60]
  wire [7:0] _GEN_5638 = 8'h0 < length_2 ? _GEN_5478 : _GEN_5318; // @[executor.scala 308:60]
  wire [7:0] _GEN_5639 = 8'h0 < length_2 ? _GEN_5479 : _GEN_5319; // @[executor.scala 308:60]
  wire [7:0] _GEN_5640 = 8'h0 < length_2 ? _GEN_5480 : _GEN_5320; // @[executor.scala 308:60]
  wire [7:0] _GEN_5641 = 8'h0 < length_2 ? _GEN_5481 : _GEN_5321; // @[executor.scala 308:60]
  wire [7:0] _GEN_5642 = 8'h0 < length_2 ? _GEN_5482 : _GEN_5322; // @[executor.scala 308:60]
  wire [7:0] _GEN_5643 = 8'h0 < length_2 ? _GEN_5483 : _GEN_5323; // @[executor.scala 308:60]
  wire [7:0] _GEN_5644 = 8'h0 < length_2 ? _GEN_5484 : _GEN_5324; // @[executor.scala 308:60]
  wire [7:0] _GEN_5645 = 8'h0 < length_2 ? _GEN_5485 : _GEN_5325; // @[executor.scala 308:60]
  wire [7:0] _GEN_5646 = 8'h0 < length_2 ? _GEN_5486 : _GEN_5326; // @[executor.scala 308:60]
  wire [7:0] _GEN_5647 = 8'h0 < length_2 ? _GEN_5487 : _GEN_5327; // @[executor.scala 308:60]
  wire [7:0] _GEN_5648 = 8'h0 < length_2 ? _GEN_5488 : _GEN_5328; // @[executor.scala 308:60]
  wire [7:0] _GEN_5649 = 8'h0 < length_2 ? _GEN_5489 : _GEN_5329; // @[executor.scala 308:60]
  wire [7:0] _GEN_5650 = 8'h0 < length_2 ? _GEN_5490 : _GEN_5330; // @[executor.scala 308:60]
  wire [7:0] _GEN_5651 = 8'h0 < length_2 ? _GEN_5491 : _GEN_5331; // @[executor.scala 308:60]
  wire [7:0] _GEN_5652 = 8'h0 < length_2 ? _GEN_5492 : _GEN_5332; // @[executor.scala 308:60]
  wire [7:0] _GEN_5653 = 8'h0 < length_2 ? _GEN_5493 : _GEN_5333; // @[executor.scala 308:60]
  wire [7:0] _GEN_5654 = 8'h0 < length_2 ? _GEN_5494 : _GEN_5334; // @[executor.scala 308:60]
  wire [7:0] _GEN_5655 = 8'h0 < length_2 ? _GEN_5495 : _GEN_5335; // @[executor.scala 308:60]
  wire [7:0] _GEN_5656 = 8'h0 < length_2 ? _GEN_5496 : _GEN_5336; // @[executor.scala 308:60]
  wire [7:0] _GEN_5657 = 8'h0 < length_2 ? _GEN_5497 : _GEN_5337; // @[executor.scala 308:60]
  wire [7:0] _GEN_5658 = 8'h0 < length_2 ? _GEN_5498 : _GEN_5338; // @[executor.scala 308:60]
  wire [7:0] _GEN_5659 = 8'h0 < length_2 ? _GEN_5499 : _GEN_5339; // @[executor.scala 308:60]
  wire [7:0] _GEN_5660 = 8'h0 < length_2 ? _GEN_5500 : _GEN_5340; // @[executor.scala 308:60]
  wire [7:0] _GEN_5661 = 8'h0 < length_2 ? _GEN_5501 : _GEN_5341; // @[executor.scala 308:60]
  wire [7:0] _GEN_5662 = 8'h0 < length_2 ? _GEN_5502 : _GEN_5342; // @[executor.scala 308:60]
  wire [7:0] _GEN_5663 = 8'h0 < length_2 ? _GEN_5503 : _GEN_5343; // @[executor.scala 308:60]
  wire [7:0] _GEN_5664 = 8'h0 < length_2 ? _GEN_5504 : _GEN_5344; // @[executor.scala 308:60]
  wire [7:0] _GEN_5665 = 8'h0 < length_2 ? _GEN_5505 : _GEN_5345; // @[executor.scala 308:60]
  wire [7:0] _GEN_5666 = 8'h0 < length_2 ? _GEN_5506 : _GEN_5346; // @[executor.scala 308:60]
  wire [7:0] _GEN_5667 = 8'h0 < length_2 ? _GEN_5507 : _GEN_5347; // @[executor.scala 308:60]
  wire [7:0] _GEN_5668 = 8'h0 < length_2 ? _GEN_5508 : _GEN_5348; // @[executor.scala 308:60]
  wire [7:0] _GEN_5669 = 8'h0 < length_2 ? _GEN_5509 : _GEN_5349; // @[executor.scala 308:60]
  wire [7:0] _GEN_5670 = 8'h0 < length_2 ? _GEN_5510 : _GEN_5350; // @[executor.scala 308:60]
  wire [7:0] _GEN_5671 = 8'h0 < length_2 ? _GEN_5511 : _GEN_5351; // @[executor.scala 308:60]
  wire [7:0] _GEN_5672 = 8'h0 < length_2 ? _GEN_5512 : _GEN_5352; // @[executor.scala 308:60]
  wire [7:0] _GEN_5673 = 8'h0 < length_2 ? _GEN_5513 : _GEN_5353; // @[executor.scala 308:60]
  wire [7:0] _GEN_5674 = 8'h0 < length_2 ? _GEN_5514 : _GEN_5354; // @[executor.scala 308:60]
  wire [7:0] _GEN_5675 = 8'h0 < length_2 ? _GEN_5515 : _GEN_5355; // @[executor.scala 308:60]
  wire [7:0] _GEN_5676 = 8'h0 < length_2 ? _GEN_5516 : _GEN_5356; // @[executor.scala 308:60]
  wire [7:0] _GEN_5677 = 8'h0 < length_2 ? _GEN_5517 : _GEN_5357; // @[executor.scala 308:60]
  wire [7:0] _GEN_5678 = 8'h0 < length_2 ? _GEN_5518 : _GEN_5358; // @[executor.scala 308:60]
  wire [7:0] _GEN_5679 = 8'h0 < length_2 ? _GEN_5519 : _GEN_5359; // @[executor.scala 308:60]
  wire [7:0] _GEN_5680 = 8'h0 < length_2 ? _GEN_5520 : _GEN_5360; // @[executor.scala 308:60]
  wire [7:0] _GEN_5681 = 8'h0 < length_2 ? _GEN_5521 : _GEN_5361; // @[executor.scala 308:60]
  wire [7:0] _GEN_5682 = 8'h0 < length_2 ? _GEN_5522 : _GEN_5362; // @[executor.scala 308:60]
  wire [7:0] _GEN_5683 = 8'h0 < length_2 ? _GEN_5523 : _GEN_5363; // @[executor.scala 308:60]
  wire [7:0] _GEN_5684 = 8'h0 < length_2 ? _GEN_5524 : _GEN_5364; // @[executor.scala 308:60]
  wire [7:0] _GEN_5685 = 8'h0 < length_2 ? _GEN_5525 : _GEN_5365; // @[executor.scala 308:60]
  wire [7:0] _GEN_5686 = 8'h0 < length_2 ? _GEN_5526 : _GEN_5366; // @[executor.scala 308:60]
  wire [7:0] _GEN_5687 = 8'h0 < length_2 ? _GEN_5527 : _GEN_5367; // @[executor.scala 308:60]
  wire [7:0] _GEN_5688 = 8'h0 < length_2 ? _GEN_5528 : _GEN_5368; // @[executor.scala 308:60]
  wire [7:0] _GEN_5689 = 8'h0 < length_2 ? _GEN_5529 : _GEN_5369; // @[executor.scala 308:60]
  wire [7:0] _GEN_5690 = 8'h0 < length_2 ? _GEN_5530 : _GEN_5370; // @[executor.scala 308:60]
  wire [7:0] _GEN_5691 = 8'h0 < length_2 ? _GEN_5531 : _GEN_5371; // @[executor.scala 308:60]
  wire [7:0] _GEN_5692 = 8'h0 < length_2 ? _GEN_5532 : _GEN_5372; // @[executor.scala 308:60]
  wire [7:0] _GEN_5693 = 8'h0 < length_2 ? _GEN_5533 : _GEN_5373; // @[executor.scala 308:60]
  wire [7:0] _GEN_5694 = 8'h0 < length_2 ? _GEN_5534 : _GEN_5374; // @[executor.scala 308:60]
  wire [7:0] _GEN_5695 = 8'h0 < length_2 ? _GEN_5535 : _GEN_5375; // @[executor.scala 308:60]
  wire [7:0] _GEN_5696 = 8'h0 < length_2 ? _GEN_5536 : _GEN_5376; // @[executor.scala 308:60]
  wire [7:0] _GEN_5697 = 8'h0 < length_2 ? _GEN_5537 : _GEN_5377; // @[executor.scala 308:60]
  wire [7:0] _GEN_5698 = 8'h0 < length_2 ? _GEN_5538 : _GEN_5378; // @[executor.scala 308:60]
  wire [7:0] _GEN_5699 = 8'h0 < length_2 ? _GEN_5539 : _GEN_5379; // @[executor.scala 308:60]
  wire [7:0] _GEN_5700 = 8'h0 < length_2 ? _GEN_5540 : _GEN_5380; // @[executor.scala 308:60]
  wire [7:0] _GEN_5701 = 8'h0 < length_2 ? _GEN_5541 : _GEN_5381; // @[executor.scala 308:60]
  wire [7:0] _GEN_5702 = 8'h0 < length_2 ? _GEN_5542 : _GEN_5382; // @[executor.scala 308:60]
  wire [7:0] _GEN_5703 = 8'h0 < length_2 ? _GEN_5543 : _GEN_5383; // @[executor.scala 308:60]
  wire [7:0] _GEN_5704 = 8'h0 < length_2 ? _GEN_5544 : _GEN_5384; // @[executor.scala 308:60]
  wire [7:0] _GEN_5705 = 8'h0 < length_2 ? _GEN_5545 : _GEN_5385; // @[executor.scala 308:60]
  wire [7:0] _GEN_5706 = 8'h0 < length_2 ? _GEN_5546 : _GEN_5386; // @[executor.scala 308:60]
  wire [7:0] _GEN_5707 = 8'h0 < length_2 ? _GEN_5547 : _GEN_5387; // @[executor.scala 308:60]
  wire [7:0] _GEN_5708 = 8'h0 < length_2 ? _GEN_5548 : _GEN_5388; // @[executor.scala 308:60]
  wire [7:0] _GEN_5709 = 8'h0 < length_2 ? _GEN_5549 : _GEN_5389; // @[executor.scala 308:60]
  wire [7:0] _GEN_5710 = 8'h0 < length_2 ? _GEN_5550 : _GEN_5390; // @[executor.scala 308:60]
  wire [7:0] _GEN_5711 = 8'h0 < length_2 ? _GEN_5551 : _GEN_5391; // @[executor.scala 308:60]
  wire [7:0] _GEN_5712 = 8'h0 < length_2 ? _GEN_5552 : _GEN_5392; // @[executor.scala 308:60]
  wire [7:0] _GEN_5713 = 8'h0 < length_2 ? _GEN_5553 : _GEN_5393; // @[executor.scala 308:60]
  wire [7:0] _GEN_5714 = 8'h0 < length_2 ? _GEN_5554 : _GEN_5394; // @[executor.scala 308:60]
  wire [7:0] _GEN_5715 = 8'h0 < length_2 ? _GEN_5555 : _GEN_5395; // @[executor.scala 308:60]
  wire [7:0] _GEN_5716 = 8'h0 < length_2 ? _GEN_5556 : _GEN_5396; // @[executor.scala 308:60]
  wire [7:0] _GEN_5717 = 8'h0 < length_2 ? _GEN_5557 : _GEN_5397; // @[executor.scala 308:60]
  wire [7:0] _GEN_5718 = 8'h0 < length_2 ? _GEN_5558 : _GEN_5398; // @[executor.scala 308:60]
  wire [7:0] _GEN_5719 = 8'h0 < length_2 ? _GEN_5559 : _GEN_5399; // @[executor.scala 308:60]
  wire [7:0] _GEN_5720 = 8'h0 < length_2 ? _GEN_5560 : _GEN_5400; // @[executor.scala 308:60]
  wire [7:0] _GEN_5721 = 8'h0 < length_2 ? _GEN_5561 : _GEN_5401; // @[executor.scala 308:60]
  wire [7:0] _GEN_5722 = 8'h0 < length_2 ? _GEN_5562 : _GEN_5402; // @[executor.scala 308:60]
  wire [7:0] _GEN_5723 = 8'h0 < length_2 ? _GEN_5563 : _GEN_5403; // @[executor.scala 308:60]
  wire [7:0] _GEN_5724 = 8'h0 < length_2 ? _GEN_5564 : _GEN_5404; // @[executor.scala 308:60]
  wire [7:0] _GEN_5725 = 8'h0 < length_2 ? _GEN_5565 : _GEN_5405; // @[executor.scala 308:60]
  wire [7:0] _GEN_5726 = 8'h0 < length_2 ? _GEN_5566 : _GEN_5406; // @[executor.scala 308:60]
  wire [7:0] _GEN_5727 = 8'h0 < length_2 ? _GEN_5567 : _GEN_5407; // @[executor.scala 308:60]
  wire [7:0] _GEN_5728 = 8'h0 < length_2 ? _GEN_5568 : _GEN_5408; // @[executor.scala 308:60]
  wire [7:0] _GEN_5729 = 8'h0 < length_2 ? _GEN_5569 : _GEN_5409; // @[executor.scala 308:60]
  wire [7:0] _GEN_5730 = 8'h0 < length_2 ? _GEN_5570 : _GEN_5410; // @[executor.scala 308:60]
  wire [7:0] _GEN_5731 = 8'h0 < length_2 ? _GEN_5571 : _GEN_5411; // @[executor.scala 308:60]
  wire [7:0] _GEN_5732 = 8'h0 < length_2 ? _GEN_5572 : _GEN_5412; // @[executor.scala 308:60]
  wire [7:0] _GEN_5733 = 8'h0 < length_2 ? _GEN_5573 : _GEN_5413; // @[executor.scala 308:60]
  wire [7:0] _GEN_5734 = 8'h0 < length_2 ? _GEN_5574 : _GEN_5414; // @[executor.scala 308:60]
  wire [7:0] _GEN_5735 = 8'h0 < length_2 ? _GEN_5575 : _GEN_5415; // @[executor.scala 308:60]
  wire [7:0] _GEN_5736 = 8'h0 < length_2 ? _GEN_5576 : _GEN_5416; // @[executor.scala 308:60]
  wire [7:0] _GEN_5737 = 8'h0 < length_2 ? _GEN_5577 : _GEN_5417; // @[executor.scala 308:60]
  wire [7:0] _GEN_5738 = 8'h0 < length_2 ? _GEN_5578 : _GEN_5418; // @[executor.scala 308:60]
  wire [7:0] _GEN_5739 = 8'h0 < length_2 ? _GEN_5579 : _GEN_5419; // @[executor.scala 308:60]
  wire [7:0] _GEN_5740 = 8'h0 < length_2 ? _GEN_5580 : _GEN_5420; // @[executor.scala 308:60]
  wire [7:0] _GEN_5741 = 8'h0 < length_2 ? _GEN_5581 : _GEN_5421; // @[executor.scala 308:60]
  wire [7:0] _GEN_5742 = 8'h0 < length_2 ? _GEN_5582 : _GEN_5422; // @[executor.scala 308:60]
  wire [7:0] _GEN_5743 = 8'h0 < length_2 ? _GEN_5583 : _GEN_5423; // @[executor.scala 308:60]
  wire [7:0] _GEN_5744 = 8'h0 < length_2 ? _GEN_5584 : _GEN_5424; // @[executor.scala 308:60]
  wire [7:0] _GEN_5745 = 8'h0 < length_2 ? _GEN_5585 : _GEN_5425; // @[executor.scala 308:60]
  wire [7:0] _GEN_5746 = 8'h0 < length_2 ? _GEN_5586 : _GEN_5426; // @[executor.scala 308:60]
  wire [7:0] _GEN_5747 = 8'h0 < length_2 ? _GEN_5587 : _GEN_5427; // @[executor.scala 308:60]
  wire [7:0] _GEN_5748 = 8'h0 < length_2 ? _GEN_5588 : _GEN_5428; // @[executor.scala 308:60]
  wire [7:0] _GEN_5749 = 8'h0 < length_2 ? _GEN_5589 : _GEN_5429; // @[executor.scala 308:60]
  wire [7:0] _GEN_5750 = 8'h0 < length_2 ? _GEN_5590 : _GEN_5430; // @[executor.scala 308:60]
  wire [7:0] _GEN_5751 = 8'h0 < length_2 ? _GEN_5591 : _GEN_5431; // @[executor.scala 308:60]
  wire [7:0] _GEN_5752 = 8'h0 < length_2 ? _GEN_5592 : _GEN_5432; // @[executor.scala 308:60]
  wire [7:0] _GEN_5753 = 8'h0 < length_2 ? _GEN_5593 : _GEN_5433; // @[executor.scala 308:60]
  wire [7:0] _GEN_5754 = 8'h0 < length_2 ? _GEN_5594 : _GEN_5434; // @[executor.scala 308:60]
  wire [7:0] _GEN_5755 = 8'h0 < length_2 ? _GEN_5595 : _GEN_5435; // @[executor.scala 308:60]
  wire [7:0] _GEN_5756 = 8'h0 < length_2 ? _GEN_5596 : _GEN_5436; // @[executor.scala 308:60]
  wire [7:0] _GEN_5757 = 8'h0 < length_2 ? _GEN_5597 : _GEN_5437; // @[executor.scala 308:60]
  wire [7:0] _GEN_5758 = 8'h0 < length_2 ? _GEN_5598 : _GEN_5438; // @[executor.scala 308:60]
  wire [7:0] _GEN_5759 = 8'h0 < length_2 ? _GEN_5599 : _GEN_5439; // @[executor.scala 308:60]
  wire [7:0] _GEN_5760 = 8'h0 < length_2 ? _GEN_5600 : _GEN_5440; // @[executor.scala 308:60]
  wire [7:0] _GEN_5761 = 8'h0 < length_2 ? _GEN_5601 : _GEN_5441; // @[executor.scala 308:60]
  wire [7:0] _GEN_5762 = 8'h0 < length_2 ? _GEN_5602 : _GEN_5442; // @[executor.scala 308:60]
  wire [7:0] _GEN_5763 = 8'h0 < length_2 ? _GEN_5603 : _GEN_5443; // @[executor.scala 308:60]
  wire [7:0] field_byte_17 = field_2[55:48]; // @[executor.scala 305:57]
  wire [7:0] total_offset_17 = offset_2 + 8'h1; // @[executor.scala 307:57]
  wire [7:0] _GEN_5764 = 8'h0 == total_offset_17 ? field_byte_17 : _GEN_5604; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5765 = 8'h1 == total_offset_17 ? field_byte_17 : _GEN_5605; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5766 = 8'h2 == total_offset_17 ? field_byte_17 : _GEN_5606; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5767 = 8'h3 == total_offset_17 ? field_byte_17 : _GEN_5607; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5768 = 8'h4 == total_offset_17 ? field_byte_17 : _GEN_5608; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5769 = 8'h5 == total_offset_17 ? field_byte_17 : _GEN_5609; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5770 = 8'h6 == total_offset_17 ? field_byte_17 : _GEN_5610; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5771 = 8'h7 == total_offset_17 ? field_byte_17 : _GEN_5611; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5772 = 8'h8 == total_offset_17 ? field_byte_17 : _GEN_5612; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5773 = 8'h9 == total_offset_17 ? field_byte_17 : _GEN_5613; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5774 = 8'ha == total_offset_17 ? field_byte_17 : _GEN_5614; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5775 = 8'hb == total_offset_17 ? field_byte_17 : _GEN_5615; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5776 = 8'hc == total_offset_17 ? field_byte_17 : _GEN_5616; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5777 = 8'hd == total_offset_17 ? field_byte_17 : _GEN_5617; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5778 = 8'he == total_offset_17 ? field_byte_17 : _GEN_5618; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5779 = 8'hf == total_offset_17 ? field_byte_17 : _GEN_5619; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5780 = 8'h10 == total_offset_17 ? field_byte_17 : _GEN_5620; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5781 = 8'h11 == total_offset_17 ? field_byte_17 : _GEN_5621; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5782 = 8'h12 == total_offset_17 ? field_byte_17 : _GEN_5622; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5783 = 8'h13 == total_offset_17 ? field_byte_17 : _GEN_5623; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5784 = 8'h14 == total_offset_17 ? field_byte_17 : _GEN_5624; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5785 = 8'h15 == total_offset_17 ? field_byte_17 : _GEN_5625; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5786 = 8'h16 == total_offset_17 ? field_byte_17 : _GEN_5626; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5787 = 8'h17 == total_offset_17 ? field_byte_17 : _GEN_5627; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5788 = 8'h18 == total_offset_17 ? field_byte_17 : _GEN_5628; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5789 = 8'h19 == total_offset_17 ? field_byte_17 : _GEN_5629; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5790 = 8'h1a == total_offset_17 ? field_byte_17 : _GEN_5630; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5791 = 8'h1b == total_offset_17 ? field_byte_17 : _GEN_5631; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5792 = 8'h1c == total_offset_17 ? field_byte_17 : _GEN_5632; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5793 = 8'h1d == total_offset_17 ? field_byte_17 : _GEN_5633; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5794 = 8'h1e == total_offset_17 ? field_byte_17 : _GEN_5634; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5795 = 8'h1f == total_offset_17 ? field_byte_17 : _GEN_5635; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5796 = 8'h20 == total_offset_17 ? field_byte_17 : _GEN_5636; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5797 = 8'h21 == total_offset_17 ? field_byte_17 : _GEN_5637; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5798 = 8'h22 == total_offset_17 ? field_byte_17 : _GEN_5638; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5799 = 8'h23 == total_offset_17 ? field_byte_17 : _GEN_5639; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5800 = 8'h24 == total_offset_17 ? field_byte_17 : _GEN_5640; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5801 = 8'h25 == total_offset_17 ? field_byte_17 : _GEN_5641; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5802 = 8'h26 == total_offset_17 ? field_byte_17 : _GEN_5642; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5803 = 8'h27 == total_offset_17 ? field_byte_17 : _GEN_5643; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5804 = 8'h28 == total_offset_17 ? field_byte_17 : _GEN_5644; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5805 = 8'h29 == total_offset_17 ? field_byte_17 : _GEN_5645; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5806 = 8'h2a == total_offset_17 ? field_byte_17 : _GEN_5646; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5807 = 8'h2b == total_offset_17 ? field_byte_17 : _GEN_5647; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5808 = 8'h2c == total_offset_17 ? field_byte_17 : _GEN_5648; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5809 = 8'h2d == total_offset_17 ? field_byte_17 : _GEN_5649; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5810 = 8'h2e == total_offset_17 ? field_byte_17 : _GEN_5650; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5811 = 8'h2f == total_offset_17 ? field_byte_17 : _GEN_5651; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5812 = 8'h30 == total_offset_17 ? field_byte_17 : _GEN_5652; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5813 = 8'h31 == total_offset_17 ? field_byte_17 : _GEN_5653; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5814 = 8'h32 == total_offset_17 ? field_byte_17 : _GEN_5654; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5815 = 8'h33 == total_offset_17 ? field_byte_17 : _GEN_5655; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5816 = 8'h34 == total_offset_17 ? field_byte_17 : _GEN_5656; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5817 = 8'h35 == total_offset_17 ? field_byte_17 : _GEN_5657; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5818 = 8'h36 == total_offset_17 ? field_byte_17 : _GEN_5658; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5819 = 8'h37 == total_offset_17 ? field_byte_17 : _GEN_5659; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5820 = 8'h38 == total_offset_17 ? field_byte_17 : _GEN_5660; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5821 = 8'h39 == total_offset_17 ? field_byte_17 : _GEN_5661; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5822 = 8'h3a == total_offset_17 ? field_byte_17 : _GEN_5662; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5823 = 8'h3b == total_offset_17 ? field_byte_17 : _GEN_5663; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5824 = 8'h3c == total_offset_17 ? field_byte_17 : _GEN_5664; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5825 = 8'h3d == total_offset_17 ? field_byte_17 : _GEN_5665; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5826 = 8'h3e == total_offset_17 ? field_byte_17 : _GEN_5666; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5827 = 8'h3f == total_offset_17 ? field_byte_17 : _GEN_5667; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5828 = 8'h40 == total_offset_17 ? field_byte_17 : _GEN_5668; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5829 = 8'h41 == total_offset_17 ? field_byte_17 : _GEN_5669; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5830 = 8'h42 == total_offset_17 ? field_byte_17 : _GEN_5670; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5831 = 8'h43 == total_offset_17 ? field_byte_17 : _GEN_5671; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5832 = 8'h44 == total_offset_17 ? field_byte_17 : _GEN_5672; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5833 = 8'h45 == total_offset_17 ? field_byte_17 : _GEN_5673; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5834 = 8'h46 == total_offset_17 ? field_byte_17 : _GEN_5674; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5835 = 8'h47 == total_offset_17 ? field_byte_17 : _GEN_5675; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5836 = 8'h48 == total_offset_17 ? field_byte_17 : _GEN_5676; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5837 = 8'h49 == total_offset_17 ? field_byte_17 : _GEN_5677; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5838 = 8'h4a == total_offset_17 ? field_byte_17 : _GEN_5678; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5839 = 8'h4b == total_offset_17 ? field_byte_17 : _GEN_5679; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5840 = 8'h4c == total_offset_17 ? field_byte_17 : _GEN_5680; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5841 = 8'h4d == total_offset_17 ? field_byte_17 : _GEN_5681; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5842 = 8'h4e == total_offset_17 ? field_byte_17 : _GEN_5682; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5843 = 8'h4f == total_offset_17 ? field_byte_17 : _GEN_5683; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5844 = 8'h50 == total_offset_17 ? field_byte_17 : _GEN_5684; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5845 = 8'h51 == total_offset_17 ? field_byte_17 : _GEN_5685; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5846 = 8'h52 == total_offset_17 ? field_byte_17 : _GEN_5686; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5847 = 8'h53 == total_offset_17 ? field_byte_17 : _GEN_5687; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5848 = 8'h54 == total_offset_17 ? field_byte_17 : _GEN_5688; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5849 = 8'h55 == total_offset_17 ? field_byte_17 : _GEN_5689; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5850 = 8'h56 == total_offset_17 ? field_byte_17 : _GEN_5690; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5851 = 8'h57 == total_offset_17 ? field_byte_17 : _GEN_5691; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5852 = 8'h58 == total_offset_17 ? field_byte_17 : _GEN_5692; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5853 = 8'h59 == total_offset_17 ? field_byte_17 : _GEN_5693; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5854 = 8'h5a == total_offset_17 ? field_byte_17 : _GEN_5694; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5855 = 8'h5b == total_offset_17 ? field_byte_17 : _GEN_5695; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5856 = 8'h5c == total_offset_17 ? field_byte_17 : _GEN_5696; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5857 = 8'h5d == total_offset_17 ? field_byte_17 : _GEN_5697; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5858 = 8'h5e == total_offset_17 ? field_byte_17 : _GEN_5698; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5859 = 8'h5f == total_offset_17 ? field_byte_17 : _GEN_5699; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5860 = 8'h60 == total_offset_17 ? field_byte_17 : _GEN_5700; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5861 = 8'h61 == total_offset_17 ? field_byte_17 : _GEN_5701; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5862 = 8'h62 == total_offset_17 ? field_byte_17 : _GEN_5702; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5863 = 8'h63 == total_offset_17 ? field_byte_17 : _GEN_5703; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5864 = 8'h64 == total_offset_17 ? field_byte_17 : _GEN_5704; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5865 = 8'h65 == total_offset_17 ? field_byte_17 : _GEN_5705; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5866 = 8'h66 == total_offset_17 ? field_byte_17 : _GEN_5706; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5867 = 8'h67 == total_offset_17 ? field_byte_17 : _GEN_5707; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5868 = 8'h68 == total_offset_17 ? field_byte_17 : _GEN_5708; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5869 = 8'h69 == total_offset_17 ? field_byte_17 : _GEN_5709; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5870 = 8'h6a == total_offset_17 ? field_byte_17 : _GEN_5710; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5871 = 8'h6b == total_offset_17 ? field_byte_17 : _GEN_5711; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5872 = 8'h6c == total_offset_17 ? field_byte_17 : _GEN_5712; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5873 = 8'h6d == total_offset_17 ? field_byte_17 : _GEN_5713; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5874 = 8'h6e == total_offset_17 ? field_byte_17 : _GEN_5714; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5875 = 8'h6f == total_offset_17 ? field_byte_17 : _GEN_5715; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5876 = 8'h70 == total_offset_17 ? field_byte_17 : _GEN_5716; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5877 = 8'h71 == total_offset_17 ? field_byte_17 : _GEN_5717; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5878 = 8'h72 == total_offset_17 ? field_byte_17 : _GEN_5718; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5879 = 8'h73 == total_offset_17 ? field_byte_17 : _GEN_5719; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5880 = 8'h74 == total_offset_17 ? field_byte_17 : _GEN_5720; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5881 = 8'h75 == total_offset_17 ? field_byte_17 : _GEN_5721; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5882 = 8'h76 == total_offset_17 ? field_byte_17 : _GEN_5722; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5883 = 8'h77 == total_offset_17 ? field_byte_17 : _GEN_5723; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5884 = 8'h78 == total_offset_17 ? field_byte_17 : _GEN_5724; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5885 = 8'h79 == total_offset_17 ? field_byte_17 : _GEN_5725; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5886 = 8'h7a == total_offset_17 ? field_byte_17 : _GEN_5726; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5887 = 8'h7b == total_offset_17 ? field_byte_17 : _GEN_5727; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5888 = 8'h7c == total_offset_17 ? field_byte_17 : _GEN_5728; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5889 = 8'h7d == total_offset_17 ? field_byte_17 : _GEN_5729; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5890 = 8'h7e == total_offset_17 ? field_byte_17 : _GEN_5730; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5891 = 8'h7f == total_offset_17 ? field_byte_17 : _GEN_5731; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5892 = 8'h80 == total_offset_17 ? field_byte_17 : _GEN_5732; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5893 = 8'h81 == total_offset_17 ? field_byte_17 : _GEN_5733; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5894 = 8'h82 == total_offset_17 ? field_byte_17 : _GEN_5734; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5895 = 8'h83 == total_offset_17 ? field_byte_17 : _GEN_5735; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5896 = 8'h84 == total_offset_17 ? field_byte_17 : _GEN_5736; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5897 = 8'h85 == total_offset_17 ? field_byte_17 : _GEN_5737; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5898 = 8'h86 == total_offset_17 ? field_byte_17 : _GEN_5738; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5899 = 8'h87 == total_offset_17 ? field_byte_17 : _GEN_5739; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5900 = 8'h88 == total_offset_17 ? field_byte_17 : _GEN_5740; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5901 = 8'h89 == total_offset_17 ? field_byte_17 : _GEN_5741; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5902 = 8'h8a == total_offset_17 ? field_byte_17 : _GEN_5742; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5903 = 8'h8b == total_offset_17 ? field_byte_17 : _GEN_5743; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5904 = 8'h8c == total_offset_17 ? field_byte_17 : _GEN_5744; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5905 = 8'h8d == total_offset_17 ? field_byte_17 : _GEN_5745; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5906 = 8'h8e == total_offset_17 ? field_byte_17 : _GEN_5746; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5907 = 8'h8f == total_offset_17 ? field_byte_17 : _GEN_5747; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5908 = 8'h90 == total_offset_17 ? field_byte_17 : _GEN_5748; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5909 = 8'h91 == total_offset_17 ? field_byte_17 : _GEN_5749; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5910 = 8'h92 == total_offset_17 ? field_byte_17 : _GEN_5750; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5911 = 8'h93 == total_offset_17 ? field_byte_17 : _GEN_5751; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5912 = 8'h94 == total_offset_17 ? field_byte_17 : _GEN_5752; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5913 = 8'h95 == total_offset_17 ? field_byte_17 : _GEN_5753; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5914 = 8'h96 == total_offset_17 ? field_byte_17 : _GEN_5754; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5915 = 8'h97 == total_offset_17 ? field_byte_17 : _GEN_5755; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5916 = 8'h98 == total_offset_17 ? field_byte_17 : _GEN_5756; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5917 = 8'h99 == total_offset_17 ? field_byte_17 : _GEN_5757; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5918 = 8'h9a == total_offset_17 ? field_byte_17 : _GEN_5758; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5919 = 8'h9b == total_offset_17 ? field_byte_17 : _GEN_5759; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5920 = 8'h9c == total_offset_17 ? field_byte_17 : _GEN_5760; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5921 = 8'h9d == total_offset_17 ? field_byte_17 : _GEN_5761; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5922 = 8'h9e == total_offset_17 ? field_byte_17 : _GEN_5762; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5923 = 8'h9f == total_offset_17 ? field_byte_17 : _GEN_5763; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_5924 = 8'h1 < length_2 ? _GEN_5764 : _GEN_5604; // @[executor.scala 308:60]
  wire [7:0] _GEN_5925 = 8'h1 < length_2 ? _GEN_5765 : _GEN_5605; // @[executor.scala 308:60]
  wire [7:0] _GEN_5926 = 8'h1 < length_2 ? _GEN_5766 : _GEN_5606; // @[executor.scala 308:60]
  wire [7:0] _GEN_5927 = 8'h1 < length_2 ? _GEN_5767 : _GEN_5607; // @[executor.scala 308:60]
  wire [7:0] _GEN_5928 = 8'h1 < length_2 ? _GEN_5768 : _GEN_5608; // @[executor.scala 308:60]
  wire [7:0] _GEN_5929 = 8'h1 < length_2 ? _GEN_5769 : _GEN_5609; // @[executor.scala 308:60]
  wire [7:0] _GEN_5930 = 8'h1 < length_2 ? _GEN_5770 : _GEN_5610; // @[executor.scala 308:60]
  wire [7:0] _GEN_5931 = 8'h1 < length_2 ? _GEN_5771 : _GEN_5611; // @[executor.scala 308:60]
  wire [7:0] _GEN_5932 = 8'h1 < length_2 ? _GEN_5772 : _GEN_5612; // @[executor.scala 308:60]
  wire [7:0] _GEN_5933 = 8'h1 < length_2 ? _GEN_5773 : _GEN_5613; // @[executor.scala 308:60]
  wire [7:0] _GEN_5934 = 8'h1 < length_2 ? _GEN_5774 : _GEN_5614; // @[executor.scala 308:60]
  wire [7:0] _GEN_5935 = 8'h1 < length_2 ? _GEN_5775 : _GEN_5615; // @[executor.scala 308:60]
  wire [7:0] _GEN_5936 = 8'h1 < length_2 ? _GEN_5776 : _GEN_5616; // @[executor.scala 308:60]
  wire [7:0] _GEN_5937 = 8'h1 < length_2 ? _GEN_5777 : _GEN_5617; // @[executor.scala 308:60]
  wire [7:0] _GEN_5938 = 8'h1 < length_2 ? _GEN_5778 : _GEN_5618; // @[executor.scala 308:60]
  wire [7:0] _GEN_5939 = 8'h1 < length_2 ? _GEN_5779 : _GEN_5619; // @[executor.scala 308:60]
  wire [7:0] _GEN_5940 = 8'h1 < length_2 ? _GEN_5780 : _GEN_5620; // @[executor.scala 308:60]
  wire [7:0] _GEN_5941 = 8'h1 < length_2 ? _GEN_5781 : _GEN_5621; // @[executor.scala 308:60]
  wire [7:0] _GEN_5942 = 8'h1 < length_2 ? _GEN_5782 : _GEN_5622; // @[executor.scala 308:60]
  wire [7:0] _GEN_5943 = 8'h1 < length_2 ? _GEN_5783 : _GEN_5623; // @[executor.scala 308:60]
  wire [7:0] _GEN_5944 = 8'h1 < length_2 ? _GEN_5784 : _GEN_5624; // @[executor.scala 308:60]
  wire [7:0] _GEN_5945 = 8'h1 < length_2 ? _GEN_5785 : _GEN_5625; // @[executor.scala 308:60]
  wire [7:0] _GEN_5946 = 8'h1 < length_2 ? _GEN_5786 : _GEN_5626; // @[executor.scala 308:60]
  wire [7:0] _GEN_5947 = 8'h1 < length_2 ? _GEN_5787 : _GEN_5627; // @[executor.scala 308:60]
  wire [7:0] _GEN_5948 = 8'h1 < length_2 ? _GEN_5788 : _GEN_5628; // @[executor.scala 308:60]
  wire [7:0] _GEN_5949 = 8'h1 < length_2 ? _GEN_5789 : _GEN_5629; // @[executor.scala 308:60]
  wire [7:0] _GEN_5950 = 8'h1 < length_2 ? _GEN_5790 : _GEN_5630; // @[executor.scala 308:60]
  wire [7:0] _GEN_5951 = 8'h1 < length_2 ? _GEN_5791 : _GEN_5631; // @[executor.scala 308:60]
  wire [7:0] _GEN_5952 = 8'h1 < length_2 ? _GEN_5792 : _GEN_5632; // @[executor.scala 308:60]
  wire [7:0] _GEN_5953 = 8'h1 < length_2 ? _GEN_5793 : _GEN_5633; // @[executor.scala 308:60]
  wire [7:0] _GEN_5954 = 8'h1 < length_2 ? _GEN_5794 : _GEN_5634; // @[executor.scala 308:60]
  wire [7:0] _GEN_5955 = 8'h1 < length_2 ? _GEN_5795 : _GEN_5635; // @[executor.scala 308:60]
  wire [7:0] _GEN_5956 = 8'h1 < length_2 ? _GEN_5796 : _GEN_5636; // @[executor.scala 308:60]
  wire [7:0] _GEN_5957 = 8'h1 < length_2 ? _GEN_5797 : _GEN_5637; // @[executor.scala 308:60]
  wire [7:0] _GEN_5958 = 8'h1 < length_2 ? _GEN_5798 : _GEN_5638; // @[executor.scala 308:60]
  wire [7:0] _GEN_5959 = 8'h1 < length_2 ? _GEN_5799 : _GEN_5639; // @[executor.scala 308:60]
  wire [7:0] _GEN_5960 = 8'h1 < length_2 ? _GEN_5800 : _GEN_5640; // @[executor.scala 308:60]
  wire [7:0] _GEN_5961 = 8'h1 < length_2 ? _GEN_5801 : _GEN_5641; // @[executor.scala 308:60]
  wire [7:0] _GEN_5962 = 8'h1 < length_2 ? _GEN_5802 : _GEN_5642; // @[executor.scala 308:60]
  wire [7:0] _GEN_5963 = 8'h1 < length_2 ? _GEN_5803 : _GEN_5643; // @[executor.scala 308:60]
  wire [7:0] _GEN_5964 = 8'h1 < length_2 ? _GEN_5804 : _GEN_5644; // @[executor.scala 308:60]
  wire [7:0] _GEN_5965 = 8'h1 < length_2 ? _GEN_5805 : _GEN_5645; // @[executor.scala 308:60]
  wire [7:0] _GEN_5966 = 8'h1 < length_2 ? _GEN_5806 : _GEN_5646; // @[executor.scala 308:60]
  wire [7:0] _GEN_5967 = 8'h1 < length_2 ? _GEN_5807 : _GEN_5647; // @[executor.scala 308:60]
  wire [7:0] _GEN_5968 = 8'h1 < length_2 ? _GEN_5808 : _GEN_5648; // @[executor.scala 308:60]
  wire [7:0] _GEN_5969 = 8'h1 < length_2 ? _GEN_5809 : _GEN_5649; // @[executor.scala 308:60]
  wire [7:0] _GEN_5970 = 8'h1 < length_2 ? _GEN_5810 : _GEN_5650; // @[executor.scala 308:60]
  wire [7:0] _GEN_5971 = 8'h1 < length_2 ? _GEN_5811 : _GEN_5651; // @[executor.scala 308:60]
  wire [7:0] _GEN_5972 = 8'h1 < length_2 ? _GEN_5812 : _GEN_5652; // @[executor.scala 308:60]
  wire [7:0] _GEN_5973 = 8'h1 < length_2 ? _GEN_5813 : _GEN_5653; // @[executor.scala 308:60]
  wire [7:0] _GEN_5974 = 8'h1 < length_2 ? _GEN_5814 : _GEN_5654; // @[executor.scala 308:60]
  wire [7:0] _GEN_5975 = 8'h1 < length_2 ? _GEN_5815 : _GEN_5655; // @[executor.scala 308:60]
  wire [7:0] _GEN_5976 = 8'h1 < length_2 ? _GEN_5816 : _GEN_5656; // @[executor.scala 308:60]
  wire [7:0] _GEN_5977 = 8'h1 < length_2 ? _GEN_5817 : _GEN_5657; // @[executor.scala 308:60]
  wire [7:0] _GEN_5978 = 8'h1 < length_2 ? _GEN_5818 : _GEN_5658; // @[executor.scala 308:60]
  wire [7:0] _GEN_5979 = 8'h1 < length_2 ? _GEN_5819 : _GEN_5659; // @[executor.scala 308:60]
  wire [7:0] _GEN_5980 = 8'h1 < length_2 ? _GEN_5820 : _GEN_5660; // @[executor.scala 308:60]
  wire [7:0] _GEN_5981 = 8'h1 < length_2 ? _GEN_5821 : _GEN_5661; // @[executor.scala 308:60]
  wire [7:0] _GEN_5982 = 8'h1 < length_2 ? _GEN_5822 : _GEN_5662; // @[executor.scala 308:60]
  wire [7:0] _GEN_5983 = 8'h1 < length_2 ? _GEN_5823 : _GEN_5663; // @[executor.scala 308:60]
  wire [7:0] _GEN_5984 = 8'h1 < length_2 ? _GEN_5824 : _GEN_5664; // @[executor.scala 308:60]
  wire [7:0] _GEN_5985 = 8'h1 < length_2 ? _GEN_5825 : _GEN_5665; // @[executor.scala 308:60]
  wire [7:0] _GEN_5986 = 8'h1 < length_2 ? _GEN_5826 : _GEN_5666; // @[executor.scala 308:60]
  wire [7:0] _GEN_5987 = 8'h1 < length_2 ? _GEN_5827 : _GEN_5667; // @[executor.scala 308:60]
  wire [7:0] _GEN_5988 = 8'h1 < length_2 ? _GEN_5828 : _GEN_5668; // @[executor.scala 308:60]
  wire [7:0] _GEN_5989 = 8'h1 < length_2 ? _GEN_5829 : _GEN_5669; // @[executor.scala 308:60]
  wire [7:0] _GEN_5990 = 8'h1 < length_2 ? _GEN_5830 : _GEN_5670; // @[executor.scala 308:60]
  wire [7:0] _GEN_5991 = 8'h1 < length_2 ? _GEN_5831 : _GEN_5671; // @[executor.scala 308:60]
  wire [7:0] _GEN_5992 = 8'h1 < length_2 ? _GEN_5832 : _GEN_5672; // @[executor.scala 308:60]
  wire [7:0] _GEN_5993 = 8'h1 < length_2 ? _GEN_5833 : _GEN_5673; // @[executor.scala 308:60]
  wire [7:0] _GEN_5994 = 8'h1 < length_2 ? _GEN_5834 : _GEN_5674; // @[executor.scala 308:60]
  wire [7:0] _GEN_5995 = 8'h1 < length_2 ? _GEN_5835 : _GEN_5675; // @[executor.scala 308:60]
  wire [7:0] _GEN_5996 = 8'h1 < length_2 ? _GEN_5836 : _GEN_5676; // @[executor.scala 308:60]
  wire [7:0] _GEN_5997 = 8'h1 < length_2 ? _GEN_5837 : _GEN_5677; // @[executor.scala 308:60]
  wire [7:0] _GEN_5998 = 8'h1 < length_2 ? _GEN_5838 : _GEN_5678; // @[executor.scala 308:60]
  wire [7:0] _GEN_5999 = 8'h1 < length_2 ? _GEN_5839 : _GEN_5679; // @[executor.scala 308:60]
  wire [7:0] _GEN_6000 = 8'h1 < length_2 ? _GEN_5840 : _GEN_5680; // @[executor.scala 308:60]
  wire [7:0] _GEN_6001 = 8'h1 < length_2 ? _GEN_5841 : _GEN_5681; // @[executor.scala 308:60]
  wire [7:0] _GEN_6002 = 8'h1 < length_2 ? _GEN_5842 : _GEN_5682; // @[executor.scala 308:60]
  wire [7:0] _GEN_6003 = 8'h1 < length_2 ? _GEN_5843 : _GEN_5683; // @[executor.scala 308:60]
  wire [7:0] _GEN_6004 = 8'h1 < length_2 ? _GEN_5844 : _GEN_5684; // @[executor.scala 308:60]
  wire [7:0] _GEN_6005 = 8'h1 < length_2 ? _GEN_5845 : _GEN_5685; // @[executor.scala 308:60]
  wire [7:0] _GEN_6006 = 8'h1 < length_2 ? _GEN_5846 : _GEN_5686; // @[executor.scala 308:60]
  wire [7:0] _GEN_6007 = 8'h1 < length_2 ? _GEN_5847 : _GEN_5687; // @[executor.scala 308:60]
  wire [7:0] _GEN_6008 = 8'h1 < length_2 ? _GEN_5848 : _GEN_5688; // @[executor.scala 308:60]
  wire [7:0] _GEN_6009 = 8'h1 < length_2 ? _GEN_5849 : _GEN_5689; // @[executor.scala 308:60]
  wire [7:0] _GEN_6010 = 8'h1 < length_2 ? _GEN_5850 : _GEN_5690; // @[executor.scala 308:60]
  wire [7:0] _GEN_6011 = 8'h1 < length_2 ? _GEN_5851 : _GEN_5691; // @[executor.scala 308:60]
  wire [7:0] _GEN_6012 = 8'h1 < length_2 ? _GEN_5852 : _GEN_5692; // @[executor.scala 308:60]
  wire [7:0] _GEN_6013 = 8'h1 < length_2 ? _GEN_5853 : _GEN_5693; // @[executor.scala 308:60]
  wire [7:0] _GEN_6014 = 8'h1 < length_2 ? _GEN_5854 : _GEN_5694; // @[executor.scala 308:60]
  wire [7:0] _GEN_6015 = 8'h1 < length_2 ? _GEN_5855 : _GEN_5695; // @[executor.scala 308:60]
  wire [7:0] _GEN_6016 = 8'h1 < length_2 ? _GEN_5856 : _GEN_5696; // @[executor.scala 308:60]
  wire [7:0] _GEN_6017 = 8'h1 < length_2 ? _GEN_5857 : _GEN_5697; // @[executor.scala 308:60]
  wire [7:0] _GEN_6018 = 8'h1 < length_2 ? _GEN_5858 : _GEN_5698; // @[executor.scala 308:60]
  wire [7:0] _GEN_6019 = 8'h1 < length_2 ? _GEN_5859 : _GEN_5699; // @[executor.scala 308:60]
  wire [7:0] _GEN_6020 = 8'h1 < length_2 ? _GEN_5860 : _GEN_5700; // @[executor.scala 308:60]
  wire [7:0] _GEN_6021 = 8'h1 < length_2 ? _GEN_5861 : _GEN_5701; // @[executor.scala 308:60]
  wire [7:0] _GEN_6022 = 8'h1 < length_2 ? _GEN_5862 : _GEN_5702; // @[executor.scala 308:60]
  wire [7:0] _GEN_6023 = 8'h1 < length_2 ? _GEN_5863 : _GEN_5703; // @[executor.scala 308:60]
  wire [7:0] _GEN_6024 = 8'h1 < length_2 ? _GEN_5864 : _GEN_5704; // @[executor.scala 308:60]
  wire [7:0] _GEN_6025 = 8'h1 < length_2 ? _GEN_5865 : _GEN_5705; // @[executor.scala 308:60]
  wire [7:0] _GEN_6026 = 8'h1 < length_2 ? _GEN_5866 : _GEN_5706; // @[executor.scala 308:60]
  wire [7:0] _GEN_6027 = 8'h1 < length_2 ? _GEN_5867 : _GEN_5707; // @[executor.scala 308:60]
  wire [7:0] _GEN_6028 = 8'h1 < length_2 ? _GEN_5868 : _GEN_5708; // @[executor.scala 308:60]
  wire [7:0] _GEN_6029 = 8'h1 < length_2 ? _GEN_5869 : _GEN_5709; // @[executor.scala 308:60]
  wire [7:0] _GEN_6030 = 8'h1 < length_2 ? _GEN_5870 : _GEN_5710; // @[executor.scala 308:60]
  wire [7:0] _GEN_6031 = 8'h1 < length_2 ? _GEN_5871 : _GEN_5711; // @[executor.scala 308:60]
  wire [7:0] _GEN_6032 = 8'h1 < length_2 ? _GEN_5872 : _GEN_5712; // @[executor.scala 308:60]
  wire [7:0] _GEN_6033 = 8'h1 < length_2 ? _GEN_5873 : _GEN_5713; // @[executor.scala 308:60]
  wire [7:0] _GEN_6034 = 8'h1 < length_2 ? _GEN_5874 : _GEN_5714; // @[executor.scala 308:60]
  wire [7:0] _GEN_6035 = 8'h1 < length_2 ? _GEN_5875 : _GEN_5715; // @[executor.scala 308:60]
  wire [7:0] _GEN_6036 = 8'h1 < length_2 ? _GEN_5876 : _GEN_5716; // @[executor.scala 308:60]
  wire [7:0] _GEN_6037 = 8'h1 < length_2 ? _GEN_5877 : _GEN_5717; // @[executor.scala 308:60]
  wire [7:0] _GEN_6038 = 8'h1 < length_2 ? _GEN_5878 : _GEN_5718; // @[executor.scala 308:60]
  wire [7:0] _GEN_6039 = 8'h1 < length_2 ? _GEN_5879 : _GEN_5719; // @[executor.scala 308:60]
  wire [7:0] _GEN_6040 = 8'h1 < length_2 ? _GEN_5880 : _GEN_5720; // @[executor.scala 308:60]
  wire [7:0] _GEN_6041 = 8'h1 < length_2 ? _GEN_5881 : _GEN_5721; // @[executor.scala 308:60]
  wire [7:0] _GEN_6042 = 8'h1 < length_2 ? _GEN_5882 : _GEN_5722; // @[executor.scala 308:60]
  wire [7:0] _GEN_6043 = 8'h1 < length_2 ? _GEN_5883 : _GEN_5723; // @[executor.scala 308:60]
  wire [7:0] _GEN_6044 = 8'h1 < length_2 ? _GEN_5884 : _GEN_5724; // @[executor.scala 308:60]
  wire [7:0] _GEN_6045 = 8'h1 < length_2 ? _GEN_5885 : _GEN_5725; // @[executor.scala 308:60]
  wire [7:0] _GEN_6046 = 8'h1 < length_2 ? _GEN_5886 : _GEN_5726; // @[executor.scala 308:60]
  wire [7:0] _GEN_6047 = 8'h1 < length_2 ? _GEN_5887 : _GEN_5727; // @[executor.scala 308:60]
  wire [7:0] _GEN_6048 = 8'h1 < length_2 ? _GEN_5888 : _GEN_5728; // @[executor.scala 308:60]
  wire [7:0] _GEN_6049 = 8'h1 < length_2 ? _GEN_5889 : _GEN_5729; // @[executor.scala 308:60]
  wire [7:0] _GEN_6050 = 8'h1 < length_2 ? _GEN_5890 : _GEN_5730; // @[executor.scala 308:60]
  wire [7:0] _GEN_6051 = 8'h1 < length_2 ? _GEN_5891 : _GEN_5731; // @[executor.scala 308:60]
  wire [7:0] _GEN_6052 = 8'h1 < length_2 ? _GEN_5892 : _GEN_5732; // @[executor.scala 308:60]
  wire [7:0] _GEN_6053 = 8'h1 < length_2 ? _GEN_5893 : _GEN_5733; // @[executor.scala 308:60]
  wire [7:0] _GEN_6054 = 8'h1 < length_2 ? _GEN_5894 : _GEN_5734; // @[executor.scala 308:60]
  wire [7:0] _GEN_6055 = 8'h1 < length_2 ? _GEN_5895 : _GEN_5735; // @[executor.scala 308:60]
  wire [7:0] _GEN_6056 = 8'h1 < length_2 ? _GEN_5896 : _GEN_5736; // @[executor.scala 308:60]
  wire [7:0] _GEN_6057 = 8'h1 < length_2 ? _GEN_5897 : _GEN_5737; // @[executor.scala 308:60]
  wire [7:0] _GEN_6058 = 8'h1 < length_2 ? _GEN_5898 : _GEN_5738; // @[executor.scala 308:60]
  wire [7:0] _GEN_6059 = 8'h1 < length_2 ? _GEN_5899 : _GEN_5739; // @[executor.scala 308:60]
  wire [7:0] _GEN_6060 = 8'h1 < length_2 ? _GEN_5900 : _GEN_5740; // @[executor.scala 308:60]
  wire [7:0] _GEN_6061 = 8'h1 < length_2 ? _GEN_5901 : _GEN_5741; // @[executor.scala 308:60]
  wire [7:0] _GEN_6062 = 8'h1 < length_2 ? _GEN_5902 : _GEN_5742; // @[executor.scala 308:60]
  wire [7:0] _GEN_6063 = 8'h1 < length_2 ? _GEN_5903 : _GEN_5743; // @[executor.scala 308:60]
  wire [7:0] _GEN_6064 = 8'h1 < length_2 ? _GEN_5904 : _GEN_5744; // @[executor.scala 308:60]
  wire [7:0] _GEN_6065 = 8'h1 < length_2 ? _GEN_5905 : _GEN_5745; // @[executor.scala 308:60]
  wire [7:0] _GEN_6066 = 8'h1 < length_2 ? _GEN_5906 : _GEN_5746; // @[executor.scala 308:60]
  wire [7:0] _GEN_6067 = 8'h1 < length_2 ? _GEN_5907 : _GEN_5747; // @[executor.scala 308:60]
  wire [7:0] _GEN_6068 = 8'h1 < length_2 ? _GEN_5908 : _GEN_5748; // @[executor.scala 308:60]
  wire [7:0] _GEN_6069 = 8'h1 < length_2 ? _GEN_5909 : _GEN_5749; // @[executor.scala 308:60]
  wire [7:0] _GEN_6070 = 8'h1 < length_2 ? _GEN_5910 : _GEN_5750; // @[executor.scala 308:60]
  wire [7:0] _GEN_6071 = 8'h1 < length_2 ? _GEN_5911 : _GEN_5751; // @[executor.scala 308:60]
  wire [7:0] _GEN_6072 = 8'h1 < length_2 ? _GEN_5912 : _GEN_5752; // @[executor.scala 308:60]
  wire [7:0] _GEN_6073 = 8'h1 < length_2 ? _GEN_5913 : _GEN_5753; // @[executor.scala 308:60]
  wire [7:0] _GEN_6074 = 8'h1 < length_2 ? _GEN_5914 : _GEN_5754; // @[executor.scala 308:60]
  wire [7:0] _GEN_6075 = 8'h1 < length_2 ? _GEN_5915 : _GEN_5755; // @[executor.scala 308:60]
  wire [7:0] _GEN_6076 = 8'h1 < length_2 ? _GEN_5916 : _GEN_5756; // @[executor.scala 308:60]
  wire [7:0] _GEN_6077 = 8'h1 < length_2 ? _GEN_5917 : _GEN_5757; // @[executor.scala 308:60]
  wire [7:0] _GEN_6078 = 8'h1 < length_2 ? _GEN_5918 : _GEN_5758; // @[executor.scala 308:60]
  wire [7:0] _GEN_6079 = 8'h1 < length_2 ? _GEN_5919 : _GEN_5759; // @[executor.scala 308:60]
  wire [7:0] _GEN_6080 = 8'h1 < length_2 ? _GEN_5920 : _GEN_5760; // @[executor.scala 308:60]
  wire [7:0] _GEN_6081 = 8'h1 < length_2 ? _GEN_5921 : _GEN_5761; // @[executor.scala 308:60]
  wire [7:0] _GEN_6082 = 8'h1 < length_2 ? _GEN_5922 : _GEN_5762; // @[executor.scala 308:60]
  wire [7:0] _GEN_6083 = 8'h1 < length_2 ? _GEN_5923 : _GEN_5763; // @[executor.scala 308:60]
  wire [7:0] field_byte_18 = field_2[47:40]; // @[executor.scala 305:57]
  wire [7:0] total_offset_18 = offset_2 + 8'h2; // @[executor.scala 307:57]
  wire [7:0] _GEN_6084 = 8'h0 == total_offset_18 ? field_byte_18 : _GEN_5924; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6085 = 8'h1 == total_offset_18 ? field_byte_18 : _GEN_5925; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6086 = 8'h2 == total_offset_18 ? field_byte_18 : _GEN_5926; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6087 = 8'h3 == total_offset_18 ? field_byte_18 : _GEN_5927; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6088 = 8'h4 == total_offset_18 ? field_byte_18 : _GEN_5928; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6089 = 8'h5 == total_offset_18 ? field_byte_18 : _GEN_5929; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6090 = 8'h6 == total_offset_18 ? field_byte_18 : _GEN_5930; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6091 = 8'h7 == total_offset_18 ? field_byte_18 : _GEN_5931; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6092 = 8'h8 == total_offset_18 ? field_byte_18 : _GEN_5932; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6093 = 8'h9 == total_offset_18 ? field_byte_18 : _GEN_5933; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6094 = 8'ha == total_offset_18 ? field_byte_18 : _GEN_5934; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6095 = 8'hb == total_offset_18 ? field_byte_18 : _GEN_5935; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6096 = 8'hc == total_offset_18 ? field_byte_18 : _GEN_5936; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6097 = 8'hd == total_offset_18 ? field_byte_18 : _GEN_5937; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6098 = 8'he == total_offset_18 ? field_byte_18 : _GEN_5938; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6099 = 8'hf == total_offset_18 ? field_byte_18 : _GEN_5939; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6100 = 8'h10 == total_offset_18 ? field_byte_18 : _GEN_5940; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6101 = 8'h11 == total_offset_18 ? field_byte_18 : _GEN_5941; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6102 = 8'h12 == total_offset_18 ? field_byte_18 : _GEN_5942; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6103 = 8'h13 == total_offset_18 ? field_byte_18 : _GEN_5943; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6104 = 8'h14 == total_offset_18 ? field_byte_18 : _GEN_5944; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6105 = 8'h15 == total_offset_18 ? field_byte_18 : _GEN_5945; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6106 = 8'h16 == total_offset_18 ? field_byte_18 : _GEN_5946; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6107 = 8'h17 == total_offset_18 ? field_byte_18 : _GEN_5947; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6108 = 8'h18 == total_offset_18 ? field_byte_18 : _GEN_5948; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6109 = 8'h19 == total_offset_18 ? field_byte_18 : _GEN_5949; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6110 = 8'h1a == total_offset_18 ? field_byte_18 : _GEN_5950; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6111 = 8'h1b == total_offset_18 ? field_byte_18 : _GEN_5951; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6112 = 8'h1c == total_offset_18 ? field_byte_18 : _GEN_5952; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6113 = 8'h1d == total_offset_18 ? field_byte_18 : _GEN_5953; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6114 = 8'h1e == total_offset_18 ? field_byte_18 : _GEN_5954; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6115 = 8'h1f == total_offset_18 ? field_byte_18 : _GEN_5955; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6116 = 8'h20 == total_offset_18 ? field_byte_18 : _GEN_5956; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6117 = 8'h21 == total_offset_18 ? field_byte_18 : _GEN_5957; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6118 = 8'h22 == total_offset_18 ? field_byte_18 : _GEN_5958; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6119 = 8'h23 == total_offset_18 ? field_byte_18 : _GEN_5959; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6120 = 8'h24 == total_offset_18 ? field_byte_18 : _GEN_5960; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6121 = 8'h25 == total_offset_18 ? field_byte_18 : _GEN_5961; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6122 = 8'h26 == total_offset_18 ? field_byte_18 : _GEN_5962; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6123 = 8'h27 == total_offset_18 ? field_byte_18 : _GEN_5963; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6124 = 8'h28 == total_offset_18 ? field_byte_18 : _GEN_5964; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6125 = 8'h29 == total_offset_18 ? field_byte_18 : _GEN_5965; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6126 = 8'h2a == total_offset_18 ? field_byte_18 : _GEN_5966; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6127 = 8'h2b == total_offset_18 ? field_byte_18 : _GEN_5967; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6128 = 8'h2c == total_offset_18 ? field_byte_18 : _GEN_5968; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6129 = 8'h2d == total_offset_18 ? field_byte_18 : _GEN_5969; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6130 = 8'h2e == total_offset_18 ? field_byte_18 : _GEN_5970; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6131 = 8'h2f == total_offset_18 ? field_byte_18 : _GEN_5971; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6132 = 8'h30 == total_offset_18 ? field_byte_18 : _GEN_5972; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6133 = 8'h31 == total_offset_18 ? field_byte_18 : _GEN_5973; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6134 = 8'h32 == total_offset_18 ? field_byte_18 : _GEN_5974; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6135 = 8'h33 == total_offset_18 ? field_byte_18 : _GEN_5975; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6136 = 8'h34 == total_offset_18 ? field_byte_18 : _GEN_5976; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6137 = 8'h35 == total_offset_18 ? field_byte_18 : _GEN_5977; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6138 = 8'h36 == total_offset_18 ? field_byte_18 : _GEN_5978; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6139 = 8'h37 == total_offset_18 ? field_byte_18 : _GEN_5979; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6140 = 8'h38 == total_offset_18 ? field_byte_18 : _GEN_5980; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6141 = 8'h39 == total_offset_18 ? field_byte_18 : _GEN_5981; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6142 = 8'h3a == total_offset_18 ? field_byte_18 : _GEN_5982; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6143 = 8'h3b == total_offset_18 ? field_byte_18 : _GEN_5983; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6144 = 8'h3c == total_offset_18 ? field_byte_18 : _GEN_5984; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6145 = 8'h3d == total_offset_18 ? field_byte_18 : _GEN_5985; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6146 = 8'h3e == total_offset_18 ? field_byte_18 : _GEN_5986; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6147 = 8'h3f == total_offset_18 ? field_byte_18 : _GEN_5987; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6148 = 8'h40 == total_offset_18 ? field_byte_18 : _GEN_5988; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6149 = 8'h41 == total_offset_18 ? field_byte_18 : _GEN_5989; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6150 = 8'h42 == total_offset_18 ? field_byte_18 : _GEN_5990; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6151 = 8'h43 == total_offset_18 ? field_byte_18 : _GEN_5991; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6152 = 8'h44 == total_offset_18 ? field_byte_18 : _GEN_5992; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6153 = 8'h45 == total_offset_18 ? field_byte_18 : _GEN_5993; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6154 = 8'h46 == total_offset_18 ? field_byte_18 : _GEN_5994; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6155 = 8'h47 == total_offset_18 ? field_byte_18 : _GEN_5995; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6156 = 8'h48 == total_offset_18 ? field_byte_18 : _GEN_5996; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6157 = 8'h49 == total_offset_18 ? field_byte_18 : _GEN_5997; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6158 = 8'h4a == total_offset_18 ? field_byte_18 : _GEN_5998; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6159 = 8'h4b == total_offset_18 ? field_byte_18 : _GEN_5999; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6160 = 8'h4c == total_offset_18 ? field_byte_18 : _GEN_6000; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6161 = 8'h4d == total_offset_18 ? field_byte_18 : _GEN_6001; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6162 = 8'h4e == total_offset_18 ? field_byte_18 : _GEN_6002; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6163 = 8'h4f == total_offset_18 ? field_byte_18 : _GEN_6003; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6164 = 8'h50 == total_offset_18 ? field_byte_18 : _GEN_6004; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6165 = 8'h51 == total_offset_18 ? field_byte_18 : _GEN_6005; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6166 = 8'h52 == total_offset_18 ? field_byte_18 : _GEN_6006; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6167 = 8'h53 == total_offset_18 ? field_byte_18 : _GEN_6007; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6168 = 8'h54 == total_offset_18 ? field_byte_18 : _GEN_6008; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6169 = 8'h55 == total_offset_18 ? field_byte_18 : _GEN_6009; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6170 = 8'h56 == total_offset_18 ? field_byte_18 : _GEN_6010; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6171 = 8'h57 == total_offset_18 ? field_byte_18 : _GEN_6011; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6172 = 8'h58 == total_offset_18 ? field_byte_18 : _GEN_6012; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6173 = 8'h59 == total_offset_18 ? field_byte_18 : _GEN_6013; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6174 = 8'h5a == total_offset_18 ? field_byte_18 : _GEN_6014; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6175 = 8'h5b == total_offset_18 ? field_byte_18 : _GEN_6015; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6176 = 8'h5c == total_offset_18 ? field_byte_18 : _GEN_6016; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6177 = 8'h5d == total_offset_18 ? field_byte_18 : _GEN_6017; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6178 = 8'h5e == total_offset_18 ? field_byte_18 : _GEN_6018; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6179 = 8'h5f == total_offset_18 ? field_byte_18 : _GEN_6019; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6180 = 8'h60 == total_offset_18 ? field_byte_18 : _GEN_6020; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6181 = 8'h61 == total_offset_18 ? field_byte_18 : _GEN_6021; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6182 = 8'h62 == total_offset_18 ? field_byte_18 : _GEN_6022; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6183 = 8'h63 == total_offset_18 ? field_byte_18 : _GEN_6023; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6184 = 8'h64 == total_offset_18 ? field_byte_18 : _GEN_6024; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6185 = 8'h65 == total_offset_18 ? field_byte_18 : _GEN_6025; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6186 = 8'h66 == total_offset_18 ? field_byte_18 : _GEN_6026; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6187 = 8'h67 == total_offset_18 ? field_byte_18 : _GEN_6027; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6188 = 8'h68 == total_offset_18 ? field_byte_18 : _GEN_6028; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6189 = 8'h69 == total_offset_18 ? field_byte_18 : _GEN_6029; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6190 = 8'h6a == total_offset_18 ? field_byte_18 : _GEN_6030; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6191 = 8'h6b == total_offset_18 ? field_byte_18 : _GEN_6031; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6192 = 8'h6c == total_offset_18 ? field_byte_18 : _GEN_6032; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6193 = 8'h6d == total_offset_18 ? field_byte_18 : _GEN_6033; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6194 = 8'h6e == total_offset_18 ? field_byte_18 : _GEN_6034; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6195 = 8'h6f == total_offset_18 ? field_byte_18 : _GEN_6035; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6196 = 8'h70 == total_offset_18 ? field_byte_18 : _GEN_6036; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6197 = 8'h71 == total_offset_18 ? field_byte_18 : _GEN_6037; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6198 = 8'h72 == total_offset_18 ? field_byte_18 : _GEN_6038; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6199 = 8'h73 == total_offset_18 ? field_byte_18 : _GEN_6039; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6200 = 8'h74 == total_offset_18 ? field_byte_18 : _GEN_6040; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6201 = 8'h75 == total_offset_18 ? field_byte_18 : _GEN_6041; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6202 = 8'h76 == total_offset_18 ? field_byte_18 : _GEN_6042; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6203 = 8'h77 == total_offset_18 ? field_byte_18 : _GEN_6043; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6204 = 8'h78 == total_offset_18 ? field_byte_18 : _GEN_6044; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6205 = 8'h79 == total_offset_18 ? field_byte_18 : _GEN_6045; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6206 = 8'h7a == total_offset_18 ? field_byte_18 : _GEN_6046; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6207 = 8'h7b == total_offset_18 ? field_byte_18 : _GEN_6047; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6208 = 8'h7c == total_offset_18 ? field_byte_18 : _GEN_6048; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6209 = 8'h7d == total_offset_18 ? field_byte_18 : _GEN_6049; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6210 = 8'h7e == total_offset_18 ? field_byte_18 : _GEN_6050; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6211 = 8'h7f == total_offset_18 ? field_byte_18 : _GEN_6051; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6212 = 8'h80 == total_offset_18 ? field_byte_18 : _GEN_6052; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6213 = 8'h81 == total_offset_18 ? field_byte_18 : _GEN_6053; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6214 = 8'h82 == total_offset_18 ? field_byte_18 : _GEN_6054; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6215 = 8'h83 == total_offset_18 ? field_byte_18 : _GEN_6055; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6216 = 8'h84 == total_offset_18 ? field_byte_18 : _GEN_6056; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6217 = 8'h85 == total_offset_18 ? field_byte_18 : _GEN_6057; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6218 = 8'h86 == total_offset_18 ? field_byte_18 : _GEN_6058; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6219 = 8'h87 == total_offset_18 ? field_byte_18 : _GEN_6059; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6220 = 8'h88 == total_offset_18 ? field_byte_18 : _GEN_6060; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6221 = 8'h89 == total_offset_18 ? field_byte_18 : _GEN_6061; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6222 = 8'h8a == total_offset_18 ? field_byte_18 : _GEN_6062; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6223 = 8'h8b == total_offset_18 ? field_byte_18 : _GEN_6063; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6224 = 8'h8c == total_offset_18 ? field_byte_18 : _GEN_6064; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6225 = 8'h8d == total_offset_18 ? field_byte_18 : _GEN_6065; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6226 = 8'h8e == total_offset_18 ? field_byte_18 : _GEN_6066; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6227 = 8'h8f == total_offset_18 ? field_byte_18 : _GEN_6067; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6228 = 8'h90 == total_offset_18 ? field_byte_18 : _GEN_6068; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6229 = 8'h91 == total_offset_18 ? field_byte_18 : _GEN_6069; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6230 = 8'h92 == total_offset_18 ? field_byte_18 : _GEN_6070; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6231 = 8'h93 == total_offset_18 ? field_byte_18 : _GEN_6071; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6232 = 8'h94 == total_offset_18 ? field_byte_18 : _GEN_6072; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6233 = 8'h95 == total_offset_18 ? field_byte_18 : _GEN_6073; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6234 = 8'h96 == total_offset_18 ? field_byte_18 : _GEN_6074; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6235 = 8'h97 == total_offset_18 ? field_byte_18 : _GEN_6075; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6236 = 8'h98 == total_offset_18 ? field_byte_18 : _GEN_6076; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6237 = 8'h99 == total_offset_18 ? field_byte_18 : _GEN_6077; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6238 = 8'h9a == total_offset_18 ? field_byte_18 : _GEN_6078; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6239 = 8'h9b == total_offset_18 ? field_byte_18 : _GEN_6079; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6240 = 8'h9c == total_offset_18 ? field_byte_18 : _GEN_6080; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6241 = 8'h9d == total_offset_18 ? field_byte_18 : _GEN_6081; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6242 = 8'h9e == total_offset_18 ? field_byte_18 : _GEN_6082; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6243 = 8'h9f == total_offset_18 ? field_byte_18 : _GEN_6083; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6244 = 8'h2 < length_2 ? _GEN_6084 : _GEN_5924; // @[executor.scala 308:60]
  wire [7:0] _GEN_6245 = 8'h2 < length_2 ? _GEN_6085 : _GEN_5925; // @[executor.scala 308:60]
  wire [7:0] _GEN_6246 = 8'h2 < length_2 ? _GEN_6086 : _GEN_5926; // @[executor.scala 308:60]
  wire [7:0] _GEN_6247 = 8'h2 < length_2 ? _GEN_6087 : _GEN_5927; // @[executor.scala 308:60]
  wire [7:0] _GEN_6248 = 8'h2 < length_2 ? _GEN_6088 : _GEN_5928; // @[executor.scala 308:60]
  wire [7:0] _GEN_6249 = 8'h2 < length_2 ? _GEN_6089 : _GEN_5929; // @[executor.scala 308:60]
  wire [7:0] _GEN_6250 = 8'h2 < length_2 ? _GEN_6090 : _GEN_5930; // @[executor.scala 308:60]
  wire [7:0] _GEN_6251 = 8'h2 < length_2 ? _GEN_6091 : _GEN_5931; // @[executor.scala 308:60]
  wire [7:0] _GEN_6252 = 8'h2 < length_2 ? _GEN_6092 : _GEN_5932; // @[executor.scala 308:60]
  wire [7:0] _GEN_6253 = 8'h2 < length_2 ? _GEN_6093 : _GEN_5933; // @[executor.scala 308:60]
  wire [7:0] _GEN_6254 = 8'h2 < length_2 ? _GEN_6094 : _GEN_5934; // @[executor.scala 308:60]
  wire [7:0] _GEN_6255 = 8'h2 < length_2 ? _GEN_6095 : _GEN_5935; // @[executor.scala 308:60]
  wire [7:0] _GEN_6256 = 8'h2 < length_2 ? _GEN_6096 : _GEN_5936; // @[executor.scala 308:60]
  wire [7:0] _GEN_6257 = 8'h2 < length_2 ? _GEN_6097 : _GEN_5937; // @[executor.scala 308:60]
  wire [7:0] _GEN_6258 = 8'h2 < length_2 ? _GEN_6098 : _GEN_5938; // @[executor.scala 308:60]
  wire [7:0] _GEN_6259 = 8'h2 < length_2 ? _GEN_6099 : _GEN_5939; // @[executor.scala 308:60]
  wire [7:0] _GEN_6260 = 8'h2 < length_2 ? _GEN_6100 : _GEN_5940; // @[executor.scala 308:60]
  wire [7:0] _GEN_6261 = 8'h2 < length_2 ? _GEN_6101 : _GEN_5941; // @[executor.scala 308:60]
  wire [7:0] _GEN_6262 = 8'h2 < length_2 ? _GEN_6102 : _GEN_5942; // @[executor.scala 308:60]
  wire [7:0] _GEN_6263 = 8'h2 < length_2 ? _GEN_6103 : _GEN_5943; // @[executor.scala 308:60]
  wire [7:0] _GEN_6264 = 8'h2 < length_2 ? _GEN_6104 : _GEN_5944; // @[executor.scala 308:60]
  wire [7:0] _GEN_6265 = 8'h2 < length_2 ? _GEN_6105 : _GEN_5945; // @[executor.scala 308:60]
  wire [7:0] _GEN_6266 = 8'h2 < length_2 ? _GEN_6106 : _GEN_5946; // @[executor.scala 308:60]
  wire [7:0] _GEN_6267 = 8'h2 < length_2 ? _GEN_6107 : _GEN_5947; // @[executor.scala 308:60]
  wire [7:0] _GEN_6268 = 8'h2 < length_2 ? _GEN_6108 : _GEN_5948; // @[executor.scala 308:60]
  wire [7:0] _GEN_6269 = 8'h2 < length_2 ? _GEN_6109 : _GEN_5949; // @[executor.scala 308:60]
  wire [7:0] _GEN_6270 = 8'h2 < length_2 ? _GEN_6110 : _GEN_5950; // @[executor.scala 308:60]
  wire [7:0] _GEN_6271 = 8'h2 < length_2 ? _GEN_6111 : _GEN_5951; // @[executor.scala 308:60]
  wire [7:0] _GEN_6272 = 8'h2 < length_2 ? _GEN_6112 : _GEN_5952; // @[executor.scala 308:60]
  wire [7:0] _GEN_6273 = 8'h2 < length_2 ? _GEN_6113 : _GEN_5953; // @[executor.scala 308:60]
  wire [7:0] _GEN_6274 = 8'h2 < length_2 ? _GEN_6114 : _GEN_5954; // @[executor.scala 308:60]
  wire [7:0] _GEN_6275 = 8'h2 < length_2 ? _GEN_6115 : _GEN_5955; // @[executor.scala 308:60]
  wire [7:0] _GEN_6276 = 8'h2 < length_2 ? _GEN_6116 : _GEN_5956; // @[executor.scala 308:60]
  wire [7:0] _GEN_6277 = 8'h2 < length_2 ? _GEN_6117 : _GEN_5957; // @[executor.scala 308:60]
  wire [7:0] _GEN_6278 = 8'h2 < length_2 ? _GEN_6118 : _GEN_5958; // @[executor.scala 308:60]
  wire [7:0] _GEN_6279 = 8'h2 < length_2 ? _GEN_6119 : _GEN_5959; // @[executor.scala 308:60]
  wire [7:0] _GEN_6280 = 8'h2 < length_2 ? _GEN_6120 : _GEN_5960; // @[executor.scala 308:60]
  wire [7:0] _GEN_6281 = 8'h2 < length_2 ? _GEN_6121 : _GEN_5961; // @[executor.scala 308:60]
  wire [7:0] _GEN_6282 = 8'h2 < length_2 ? _GEN_6122 : _GEN_5962; // @[executor.scala 308:60]
  wire [7:0] _GEN_6283 = 8'h2 < length_2 ? _GEN_6123 : _GEN_5963; // @[executor.scala 308:60]
  wire [7:0] _GEN_6284 = 8'h2 < length_2 ? _GEN_6124 : _GEN_5964; // @[executor.scala 308:60]
  wire [7:0] _GEN_6285 = 8'h2 < length_2 ? _GEN_6125 : _GEN_5965; // @[executor.scala 308:60]
  wire [7:0] _GEN_6286 = 8'h2 < length_2 ? _GEN_6126 : _GEN_5966; // @[executor.scala 308:60]
  wire [7:0] _GEN_6287 = 8'h2 < length_2 ? _GEN_6127 : _GEN_5967; // @[executor.scala 308:60]
  wire [7:0] _GEN_6288 = 8'h2 < length_2 ? _GEN_6128 : _GEN_5968; // @[executor.scala 308:60]
  wire [7:0] _GEN_6289 = 8'h2 < length_2 ? _GEN_6129 : _GEN_5969; // @[executor.scala 308:60]
  wire [7:0] _GEN_6290 = 8'h2 < length_2 ? _GEN_6130 : _GEN_5970; // @[executor.scala 308:60]
  wire [7:0] _GEN_6291 = 8'h2 < length_2 ? _GEN_6131 : _GEN_5971; // @[executor.scala 308:60]
  wire [7:0] _GEN_6292 = 8'h2 < length_2 ? _GEN_6132 : _GEN_5972; // @[executor.scala 308:60]
  wire [7:0] _GEN_6293 = 8'h2 < length_2 ? _GEN_6133 : _GEN_5973; // @[executor.scala 308:60]
  wire [7:0] _GEN_6294 = 8'h2 < length_2 ? _GEN_6134 : _GEN_5974; // @[executor.scala 308:60]
  wire [7:0] _GEN_6295 = 8'h2 < length_2 ? _GEN_6135 : _GEN_5975; // @[executor.scala 308:60]
  wire [7:0] _GEN_6296 = 8'h2 < length_2 ? _GEN_6136 : _GEN_5976; // @[executor.scala 308:60]
  wire [7:0] _GEN_6297 = 8'h2 < length_2 ? _GEN_6137 : _GEN_5977; // @[executor.scala 308:60]
  wire [7:0] _GEN_6298 = 8'h2 < length_2 ? _GEN_6138 : _GEN_5978; // @[executor.scala 308:60]
  wire [7:0] _GEN_6299 = 8'h2 < length_2 ? _GEN_6139 : _GEN_5979; // @[executor.scala 308:60]
  wire [7:0] _GEN_6300 = 8'h2 < length_2 ? _GEN_6140 : _GEN_5980; // @[executor.scala 308:60]
  wire [7:0] _GEN_6301 = 8'h2 < length_2 ? _GEN_6141 : _GEN_5981; // @[executor.scala 308:60]
  wire [7:0] _GEN_6302 = 8'h2 < length_2 ? _GEN_6142 : _GEN_5982; // @[executor.scala 308:60]
  wire [7:0] _GEN_6303 = 8'h2 < length_2 ? _GEN_6143 : _GEN_5983; // @[executor.scala 308:60]
  wire [7:0] _GEN_6304 = 8'h2 < length_2 ? _GEN_6144 : _GEN_5984; // @[executor.scala 308:60]
  wire [7:0] _GEN_6305 = 8'h2 < length_2 ? _GEN_6145 : _GEN_5985; // @[executor.scala 308:60]
  wire [7:0] _GEN_6306 = 8'h2 < length_2 ? _GEN_6146 : _GEN_5986; // @[executor.scala 308:60]
  wire [7:0] _GEN_6307 = 8'h2 < length_2 ? _GEN_6147 : _GEN_5987; // @[executor.scala 308:60]
  wire [7:0] _GEN_6308 = 8'h2 < length_2 ? _GEN_6148 : _GEN_5988; // @[executor.scala 308:60]
  wire [7:0] _GEN_6309 = 8'h2 < length_2 ? _GEN_6149 : _GEN_5989; // @[executor.scala 308:60]
  wire [7:0] _GEN_6310 = 8'h2 < length_2 ? _GEN_6150 : _GEN_5990; // @[executor.scala 308:60]
  wire [7:0] _GEN_6311 = 8'h2 < length_2 ? _GEN_6151 : _GEN_5991; // @[executor.scala 308:60]
  wire [7:0] _GEN_6312 = 8'h2 < length_2 ? _GEN_6152 : _GEN_5992; // @[executor.scala 308:60]
  wire [7:0] _GEN_6313 = 8'h2 < length_2 ? _GEN_6153 : _GEN_5993; // @[executor.scala 308:60]
  wire [7:0] _GEN_6314 = 8'h2 < length_2 ? _GEN_6154 : _GEN_5994; // @[executor.scala 308:60]
  wire [7:0] _GEN_6315 = 8'h2 < length_2 ? _GEN_6155 : _GEN_5995; // @[executor.scala 308:60]
  wire [7:0] _GEN_6316 = 8'h2 < length_2 ? _GEN_6156 : _GEN_5996; // @[executor.scala 308:60]
  wire [7:0] _GEN_6317 = 8'h2 < length_2 ? _GEN_6157 : _GEN_5997; // @[executor.scala 308:60]
  wire [7:0] _GEN_6318 = 8'h2 < length_2 ? _GEN_6158 : _GEN_5998; // @[executor.scala 308:60]
  wire [7:0] _GEN_6319 = 8'h2 < length_2 ? _GEN_6159 : _GEN_5999; // @[executor.scala 308:60]
  wire [7:0] _GEN_6320 = 8'h2 < length_2 ? _GEN_6160 : _GEN_6000; // @[executor.scala 308:60]
  wire [7:0] _GEN_6321 = 8'h2 < length_2 ? _GEN_6161 : _GEN_6001; // @[executor.scala 308:60]
  wire [7:0] _GEN_6322 = 8'h2 < length_2 ? _GEN_6162 : _GEN_6002; // @[executor.scala 308:60]
  wire [7:0] _GEN_6323 = 8'h2 < length_2 ? _GEN_6163 : _GEN_6003; // @[executor.scala 308:60]
  wire [7:0] _GEN_6324 = 8'h2 < length_2 ? _GEN_6164 : _GEN_6004; // @[executor.scala 308:60]
  wire [7:0] _GEN_6325 = 8'h2 < length_2 ? _GEN_6165 : _GEN_6005; // @[executor.scala 308:60]
  wire [7:0] _GEN_6326 = 8'h2 < length_2 ? _GEN_6166 : _GEN_6006; // @[executor.scala 308:60]
  wire [7:0] _GEN_6327 = 8'h2 < length_2 ? _GEN_6167 : _GEN_6007; // @[executor.scala 308:60]
  wire [7:0] _GEN_6328 = 8'h2 < length_2 ? _GEN_6168 : _GEN_6008; // @[executor.scala 308:60]
  wire [7:0] _GEN_6329 = 8'h2 < length_2 ? _GEN_6169 : _GEN_6009; // @[executor.scala 308:60]
  wire [7:0] _GEN_6330 = 8'h2 < length_2 ? _GEN_6170 : _GEN_6010; // @[executor.scala 308:60]
  wire [7:0] _GEN_6331 = 8'h2 < length_2 ? _GEN_6171 : _GEN_6011; // @[executor.scala 308:60]
  wire [7:0] _GEN_6332 = 8'h2 < length_2 ? _GEN_6172 : _GEN_6012; // @[executor.scala 308:60]
  wire [7:0] _GEN_6333 = 8'h2 < length_2 ? _GEN_6173 : _GEN_6013; // @[executor.scala 308:60]
  wire [7:0] _GEN_6334 = 8'h2 < length_2 ? _GEN_6174 : _GEN_6014; // @[executor.scala 308:60]
  wire [7:0] _GEN_6335 = 8'h2 < length_2 ? _GEN_6175 : _GEN_6015; // @[executor.scala 308:60]
  wire [7:0] _GEN_6336 = 8'h2 < length_2 ? _GEN_6176 : _GEN_6016; // @[executor.scala 308:60]
  wire [7:0] _GEN_6337 = 8'h2 < length_2 ? _GEN_6177 : _GEN_6017; // @[executor.scala 308:60]
  wire [7:0] _GEN_6338 = 8'h2 < length_2 ? _GEN_6178 : _GEN_6018; // @[executor.scala 308:60]
  wire [7:0] _GEN_6339 = 8'h2 < length_2 ? _GEN_6179 : _GEN_6019; // @[executor.scala 308:60]
  wire [7:0] _GEN_6340 = 8'h2 < length_2 ? _GEN_6180 : _GEN_6020; // @[executor.scala 308:60]
  wire [7:0] _GEN_6341 = 8'h2 < length_2 ? _GEN_6181 : _GEN_6021; // @[executor.scala 308:60]
  wire [7:0] _GEN_6342 = 8'h2 < length_2 ? _GEN_6182 : _GEN_6022; // @[executor.scala 308:60]
  wire [7:0] _GEN_6343 = 8'h2 < length_2 ? _GEN_6183 : _GEN_6023; // @[executor.scala 308:60]
  wire [7:0] _GEN_6344 = 8'h2 < length_2 ? _GEN_6184 : _GEN_6024; // @[executor.scala 308:60]
  wire [7:0] _GEN_6345 = 8'h2 < length_2 ? _GEN_6185 : _GEN_6025; // @[executor.scala 308:60]
  wire [7:0] _GEN_6346 = 8'h2 < length_2 ? _GEN_6186 : _GEN_6026; // @[executor.scala 308:60]
  wire [7:0] _GEN_6347 = 8'h2 < length_2 ? _GEN_6187 : _GEN_6027; // @[executor.scala 308:60]
  wire [7:0] _GEN_6348 = 8'h2 < length_2 ? _GEN_6188 : _GEN_6028; // @[executor.scala 308:60]
  wire [7:0] _GEN_6349 = 8'h2 < length_2 ? _GEN_6189 : _GEN_6029; // @[executor.scala 308:60]
  wire [7:0] _GEN_6350 = 8'h2 < length_2 ? _GEN_6190 : _GEN_6030; // @[executor.scala 308:60]
  wire [7:0] _GEN_6351 = 8'h2 < length_2 ? _GEN_6191 : _GEN_6031; // @[executor.scala 308:60]
  wire [7:0] _GEN_6352 = 8'h2 < length_2 ? _GEN_6192 : _GEN_6032; // @[executor.scala 308:60]
  wire [7:0] _GEN_6353 = 8'h2 < length_2 ? _GEN_6193 : _GEN_6033; // @[executor.scala 308:60]
  wire [7:0] _GEN_6354 = 8'h2 < length_2 ? _GEN_6194 : _GEN_6034; // @[executor.scala 308:60]
  wire [7:0] _GEN_6355 = 8'h2 < length_2 ? _GEN_6195 : _GEN_6035; // @[executor.scala 308:60]
  wire [7:0] _GEN_6356 = 8'h2 < length_2 ? _GEN_6196 : _GEN_6036; // @[executor.scala 308:60]
  wire [7:0] _GEN_6357 = 8'h2 < length_2 ? _GEN_6197 : _GEN_6037; // @[executor.scala 308:60]
  wire [7:0] _GEN_6358 = 8'h2 < length_2 ? _GEN_6198 : _GEN_6038; // @[executor.scala 308:60]
  wire [7:0] _GEN_6359 = 8'h2 < length_2 ? _GEN_6199 : _GEN_6039; // @[executor.scala 308:60]
  wire [7:0] _GEN_6360 = 8'h2 < length_2 ? _GEN_6200 : _GEN_6040; // @[executor.scala 308:60]
  wire [7:0] _GEN_6361 = 8'h2 < length_2 ? _GEN_6201 : _GEN_6041; // @[executor.scala 308:60]
  wire [7:0] _GEN_6362 = 8'h2 < length_2 ? _GEN_6202 : _GEN_6042; // @[executor.scala 308:60]
  wire [7:0] _GEN_6363 = 8'h2 < length_2 ? _GEN_6203 : _GEN_6043; // @[executor.scala 308:60]
  wire [7:0] _GEN_6364 = 8'h2 < length_2 ? _GEN_6204 : _GEN_6044; // @[executor.scala 308:60]
  wire [7:0] _GEN_6365 = 8'h2 < length_2 ? _GEN_6205 : _GEN_6045; // @[executor.scala 308:60]
  wire [7:0] _GEN_6366 = 8'h2 < length_2 ? _GEN_6206 : _GEN_6046; // @[executor.scala 308:60]
  wire [7:0] _GEN_6367 = 8'h2 < length_2 ? _GEN_6207 : _GEN_6047; // @[executor.scala 308:60]
  wire [7:0] _GEN_6368 = 8'h2 < length_2 ? _GEN_6208 : _GEN_6048; // @[executor.scala 308:60]
  wire [7:0] _GEN_6369 = 8'h2 < length_2 ? _GEN_6209 : _GEN_6049; // @[executor.scala 308:60]
  wire [7:0] _GEN_6370 = 8'h2 < length_2 ? _GEN_6210 : _GEN_6050; // @[executor.scala 308:60]
  wire [7:0] _GEN_6371 = 8'h2 < length_2 ? _GEN_6211 : _GEN_6051; // @[executor.scala 308:60]
  wire [7:0] _GEN_6372 = 8'h2 < length_2 ? _GEN_6212 : _GEN_6052; // @[executor.scala 308:60]
  wire [7:0] _GEN_6373 = 8'h2 < length_2 ? _GEN_6213 : _GEN_6053; // @[executor.scala 308:60]
  wire [7:0] _GEN_6374 = 8'h2 < length_2 ? _GEN_6214 : _GEN_6054; // @[executor.scala 308:60]
  wire [7:0] _GEN_6375 = 8'h2 < length_2 ? _GEN_6215 : _GEN_6055; // @[executor.scala 308:60]
  wire [7:0] _GEN_6376 = 8'h2 < length_2 ? _GEN_6216 : _GEN_6056; // @[executor.scala 308:60]
  wire [7:0] _GEN_6377 = 8'h2 < length_2 ? _GEN_6217 : _GEN_6057; // @[executor.scala 308:60]
  wire [7:0] _GEN_6378 = 8'h2 < length_2 ? _GEN_6218 : _GEN_6058; // @[executor.scala 308:60]
  wire [7:0] _GEN_6379 = 8'h2 < length_2 ? _GEN_6219 : _GEN_6059; // @[executor.scala 308:60]
  wire [7:0] _GEN_6380 = 8'h2 < length_2 ? _GEN_6220 : _GEN_6060; // @[executor.scala 308:60]
  wire [7:0] _GEN_6381 = 8'h2 < length_2 ? _GEN_6221 : _GEN_6061; // @[executor.scala 308:60]
  wire [7:0] _GEN_6382 = 8'h2 < length_2 ? _GEN_6222 : _GEN_6062; // @[executor.scala 308:60]
  wire [7:0] _GEN_6383 = 8'h2 < length_2 ? _GEN_6223 : _GEN_6063; // @[executor.scala 308:60]
  wire [7:0] _GEN_6384 = 8'h2 < length_2 ? _GEN_6224 : _GEN_6064; // @[executor.scala 308:60]
  wire [7:0] _GEN_6385 = 8'h2 < length_2 ? _GEN_6225 : _GEN_6065; // @[executor.scala 308:60]
  wire [7:0] _GEN_6386 = 8'h2 < length_2 ? _GEN_6226 : _GEN_6066; // @[executor.scala 308:60]
  wire [7:0] _GEN_6387 = 8'h2 < length_2 ? _GEN_6227 : _GEN_6067; // @[executor.scala 308:60]
  wire [7:0] _GEN_6388 = 8'h2 < length_2 ? _GEN_6228 : _GEN_6068; // @[executor.scala 308:60]
  wire [7:0] _GEN_6389 = 8'h2 < length_2 ? _GEN_6229 : _GEN_6069; // @[executor.scala 308:60]
  wire [7:0] _GEN_6390 = 8'h2 < length_2 ? _GEN_6230 : _GEN_6070; // @[executor.scala 308:60]
  wire [7:0] _GEN_6391 = 8'h2 < length_2 ? _GEN_6231 : _GEN_6071; // @[executor.scala 308:60]
  wire [7:0] _GEN_6392 = 8'h2 < length_2 ? _GEN_6232 : _GEN_6072; // @[executor.scala 308:60]
  wire [7:0] _GEN_6393 = 8'h2 < length_2 ? _GEN_6233 : _GEN_6073; // @[executor.scala 308:60]
  wire [7:0] _GEN_6394 = 8'h2 < length_2 ? _GEN_6234 : _GEN_6074; // @[executor.scala 308:60]
  wire [7:0] _GEN_6395 = 8'h2 < length_2 ? _GEN_6235 : _GEN_6075; // @[executor.scala 308:60]
  wire [7:0] _GEN_6396 = 8'h2 < length_2 ? _GEN_6236 : _GEN_6076; // @[executor.scala 308:60]
  wire [7:0] _GEN_6397 = 8'h2 < length_2 ? _GEN_6237 : _GEN_6077; // @[executor.scala 308:60]
  wire [7:0] _GEN_6398 = 8'h2 < length_2 ? _GEN_6238 : _GEN_6078; // @[executor.scala 308:60]
  wire [7:0] _GEN_6399 = 8'h2 < length_2 ? _GEN_6239 : _GEN_6079; // @[executor.scala 308:60]
  wire [7:0] _GEN_6400 = 8'h2 < length_2 ? _GEN_6240 : _GEN_6080; // @[executor.scala 308:60]
  wire [7:0] _GEN_6401 = 8'h2 < length_2 ? _GEN_6241 : _GEN_6081; // @[executor.scala 308:60]
  wire [7:0] _GEN_6402 = 8'h2 < length_2 ? _GEN_6242 : _GEN_6082; // @[executor.scala 308:60]
  wire [7:0] _GEN_6403 = 8'h2 < length_2 ? _GEN_6243 : _GEN_6083; // @[executor.scala 308:60]
  wire [7:0] field_byte_19 = field_2[39:32]; // @[executor.scala 305:57]
  wire [7:0] total_offset_19 = offset_2 + 8'h3; // @[executor.scala 307:57]
  wire [7:0] _GEN_6404 = 8'h0 == total_offset_19 ? field_byte_19 : _GEN_6244; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6405 = 8'h1 == total_offset_19 ? field_byte_19 : _GEN_6245; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6406 = 8'h2 == total_offset_19 ? field_byte_19 : _GEN_6246; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6407 = 8'h3 == total_offset_19 ? field_byte_19 : _GEN_6247; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6408 = 8'h4 == total_offset_19 ? field_byte_19 : _GEN_6248; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6409 = 8'h5 == total_offset_19 ? field_byte_19 : _GEN_6249; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6410 = 8'h6 == total_offset_19 ? field_byte_19 : _GEN_6250; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6411 = 8'h7 == total_offset_19 ? field_byte_19 : _GEN_6251; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6412 = 8'h8 == total_offset_19 ? field_byte_19 : _GEN_6252; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6413 = 8'h9 == total_offset_19 ? field_byte_19 : _GEN_6253; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6414 = 8'ha == total_offset_19 ? field_byte_19 : _GEN_6254; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6415 = 8'hb == total_offset_19 ? field_byte_19 : _GEN_6255; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6416 = 8'hc == total_offset_19 ? field_byte_19 : _GEN_6256; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6417 = 8'hd == total_offset_19 ? field_byte_19 : _GEN_6257; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6418 = 8'he == total_offset_19 ? field_byte_19 : _GEN_6258; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6419 = 8'hf == total_offset_19 ? field_byte_19 : _GEN_6259; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6420 = 8'h10 == total_offset_19 ? field_byte_19 : _GEN_6260; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6421 = 8'h11 == total_offset_19 ? field_byte_19 : _GEN_6261; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6422 = 8'h12 == total_offset_19 ? field_byte_19 : _GEN_6262; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6423 = 8'h13 == total_offset_19 ? field_byte_19 : _GEN_6263; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6424 = 8'h14 == total_offset_19 ? field_byte_19 : _GEN_6264; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6425 = 8'h15 == total_offset_19 ? field_byte_19 : _GEN_6265; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6426 = 8'h16 == total_offset_19 ? field_byte_19 : _GEN_6266; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6427 = 8'h17 == total_offset_19 ? field_byte_19 : _GEN_6267; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6428 = 8'h18 == total_offset_19 ? field_byte_19 : _GEN_6268; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6429 = 8'h19 == total_offset_19 ? field_byte_19 : _GEN_6269; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6430 = 8'h1a == total_offset_19 ? field_byte_19 : _GEN_6270; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6431 = 8'h1b == total_offset_19 ? field_byte_19 : _GEN_6271; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6432 = 8'h1c == total_offset_19 ? field_byte_19 : _GEN_6272; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6433 = 8'h1d == total_offset_19 ? field_byte_19 : _GEN_6273; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6434 = 8'h1e == total_offset_19 ? field_byte_19 : _GEN_6274; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6435 = 8'h1f == total_offset_19 ? field_byte_19 : _GEN_6275; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6436 = 8'h20 == total_offset_19 ? field_byte_19 : _GEN_6276; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6437 = 8'h21 == total_offset_19 ? field_byte_19 : _GEN_6277; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6438 = 8'h22 == total_offset_19 ? field_byte_19 : _GEN_6278; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6439 = 8'h23 == total_offset_19 ? field_byte_19 : _GEN_6279; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6440 = 8'h24 == total_offset_19 ? field_byte_19 : _GEN_6280; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6441 = 8'h25 == total_offset_19 ? field_byte_19 : _GEN_6281; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6442 = 8'h26 == total_offset_19 ? field_byte_19 : _GEN_6282; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6443 = 8'h27 == total_offset_19 ? field_byte_19 : _GEN_6283; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6444 = 8'h28 == total_offset_19 ? field_byte_19 : _GEN_6284; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6445 = 8'h29 == total_offset_19 ? field_byte_19 : _GEN_6285; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6446 = 8'h2a == total_offset_19 ? field_byte_19 : _GEN_6286; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6447 = 8'h2b == total_offset_19 ? field_byte_19 : _GEN_6287; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6448 = 8'h2c == total_offset_19 ? field_byte_19 : _GEN_6288; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6449 = 8'h2d == total_offset_19 ? field_byte_19 : _GEN_6289; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6450 = 8'h2e == total_offset_19 ? field_byte_19 : _GEN_6290; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6451 = 8'h2f == total_offset_19 ? field_byte_19 : _GEN_6291; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6452 = 8'h30 == total_offset_19 ? field_byte_19 : _GEN_6292; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6453 = 8'h31 == total_offset_19 ? field_byte_19 : _GEN_6293; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6454 = 8'h32 == total_offset_19 ? field_byte_19 : _GEN_6294; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6455 = 8'h33 == total_offset_19 ? field_byte_19 : _GEN_6295; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6456 = 8'h34 == total_offset_19 ? field_byte_19 : _GEN_6296; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6457 = 8'h35 == total_offset_19 ? field_byte_19 : _GEN_6297; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6458 = 8'h36 == total_offset_19 ? field_byte_19 : _GEN_6298; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6459 = 8'h37 == total_offset_19 ? field_byte_19 : _GEN_6299; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6460 = 8'h38 == total_offset_19 ? field_byte_19 : _GEN_6300; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6461 = 8'h39 == total_offset_19 ? field_byte_19 : _GEN_6301; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6462 = 8'h3a == total_offset_19 ? field_byte_19 : _GEN_6302; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6463 = 8'h3b == total_offset_19 ? field_byte_19 : _GEN_6303; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6464 = 8'h3c == total_offset_19 ? field_byte_19 : _GEN_6304; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6465 = 8'h3d == total_offset_19 ? field_byte_19 : _GEN_6305; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6466 = 8'h3e == total_offset_19 ? field_byte_19 : _GEN_6306; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6467 = 8'h3f == total_offset_19 ? field_byte_19 : _GEN_6307; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6468 = 8'h40 == total_offset_19 ? field_byte_19 : _GEN_6308; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6469 = 8'h41 == total_offset_19 ? field_byte_19 : _GEN_6309; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6470 = 8'h42 == total_offset_19 ? field_byte_19 : _GEN_6310; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6471 = 8'h43 == total_offset_19 ? field_byte_19 : _GEN_6311; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6472 = 8'h44 == total_offset_19 ? field_byte_19 : _GEN_6312; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6473 = 8'h45 == total_offset_19 ? field_byte_19 : _GEN_6313; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6474 = 8'h46 == total_offset_19 ? field_byte_19 : _GEN_6314; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6475 = 8'h47 == total_offset_19 ? field_byte_19 : _GEN_6315; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6476 = 8'h48 == total_offset_19 ? field_byte_19 : _GEN_6316; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6477 = 8'h49 == total_offset_19 ? field_byte_19 : _GEN_6317; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6478 = 8'h4a == total_offset_19 ? field_byte_19 : _GEN_6318; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6479 = 8'h4b == total_offset_19 ? field_byte_19 : _GEN_6319; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6480 = 8'h4c == total_offset_19 ? field_byte_19 : _GEN_6320; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6481 = 8'h4d == total_offset_19 ? field_byte_19 : _GEN_6321; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6482 = 8'h4e == total_offset_19 ? field_byte_19 : _GEN_6322; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6483 = 8'h4f == total_offset_19 ? field_byte_19 : _GEN_6323; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6484 = 8'h50 == total_offset_19 ? field_byte_19 : _GEN_6324; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6485 = 8'h51 == total_offset_19 ? field_byte_19 : _GEN_6325; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6486 = 8'h52 == total_offset_19 ? field_byte_19 : _GEN_6326; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6487 = 8'h53 == total_offset_19 ? field_byte_19 : _GEN_6327; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6488 = 8'h54 == total_offset_19 ? field_byte_19 : _GEN_6328; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6489 = 8'h55 == total_offset_19 ? field_byte_19 : _GEN_6329; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6490 = 8'h56 == total_offset_19 ? field_byte_19 : _GEN_6330; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6491 = 8'h57 == total_offset_19 ? field_byte_19 : _GEN_6331; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6492 = 8'h58 == total_offset_19 ? field_byte_19 : _GEN_6332; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6493 = 8'h59 == total_offset_19 ? field_byte_19 : _GEN_6333; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6494 = 8'h5a == total_offset_19 ? field_byte_19 : _GEN_6334; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6495 = 8'h5b == total_offset_19 ? field_byte_19 : _GEN_6335; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6496 = 8'h5c == total_offset_19 ? field_byte_19 : _GEN_6336; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6497 = 8'h5d == total_offset_19 ? field_byte_19 : _GEN_6337; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6498 = 8'h5e == total_offset_19 ? field_byte_19 : _GEN_6338; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6499 = 8'h5f == total_offset_19 ? field_byte_19 : _GEN_6339; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6500 = 8'h60 == total_offset_19 ? field_byte_19 : _GEN_6340; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6501 = 8'h61 == total_offset_19 ? field_byte_19 : _GEN_6341; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6502 = 8'h62 == total_offset_19 ? field_byte_19 : _GEN_6342; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6503 = 8'h63 == total_offset_19 ? field_byte_19 : _GEN_6343; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6504 = 8'h64 == total_offset_19 ? field_byte_19 : _GEN_6344; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6505 = 8'h65 == total_offset_19 ? field_byte_19 : _GEN_6345; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6506 = 8'h66 == total_offset_19 ? field_byte_19 : _GEN_6346; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6507 = 8'h67 == total_offset_19 ? field_byte_19 : _GEN_6347; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6508 = 8'h68 == total_offset_19 ? field_byte_19 : _GEN_6348; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6509 = 8'h69 == total_offset_19 ? field_byte_19 : _GEN_6349; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6510 = 8'h6a == total_offset_19 ? field_byte_19 : _GEN_6350; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6511 = 8'h6b == total_offset_19 ? field_byte_19 : _GEN_6351; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6512 = 8'h6c == total_offset_19 ? field_byte_19 : _GEN_6352; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6513 = 8'h6d == total_offset_19 ? field_byte_19 : _GEN_6353; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6514 = 8'h6e == total_offset_19 ? field_byte_19 : _GEN_6354; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6515 = 8'h6f == total_offset_19 ? field_byte_19 : _GEN_6355; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6516 = 8'h70 == total_offset_19 ? field_byte_19 : _GEN_6356; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6517 = 8'h71 == total_offset_19 ? field_byte_19 : _GEN_6357; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6518 = 8'h72 == total_offset_19 ? field_byte_19 : _GEN_6358; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6519 = 8'h73 == total_offset_19 ? field_byte_19 : _GEN_6359; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6520 = 8'h74 == total_offset_19 ? field_byte_19 : _GEN_6360; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6521 = 8'h75 == total_offset_19 ? field_byte_19 : _GEN_6361; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6522 = 8'h76 == total_offset_19 ? field_byte_19 : _GEN_6362; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6523 = 8'h77 == total_offset_19 ? field_byte_19 : _GEN_6363; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6524 = 8'h78 == total_offset_19 ? field_byte_19 : _GEN_6364; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6525 = 8'h79 == total_offset_19 ? field_byte_19 : _GEN_6365; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6526 = 8'h7a == total_offset_19 ? field_byte_19 : _GEN_6366; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6527 = 8'h7b == total_offset_19 ? field_byte_19 : _GEN_6367; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6528 = 8'h7c == total_offset_19 ? field_byte_19 : _GEN_6368; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6529 = 8'h7d == total_offset_19 ? field_byte_19 : _GEN_6369; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6530 = 8'h7e == total_offset_19 ? field_byte_19 : _GEN_6370; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6531 = 8'h7f == total_offset_19 ? field_byte_19 : _GEN_6371; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6532 = 8'h80 == total_offset_19 ? field_byte_19 : _GEN_6372; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6533 = 8'h81 == total_offset_19 ? field_byte_19 : _GEN_6373; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6534 = 8'h82 == total_offset_19 ? field_byte_19 : _GEN_6374; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6535 = 8'h83 == total_offset_19 ? field_byte_19 : _GEN_6375; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6536 = 8'h84 == total_offset_19 ? field_byte_19 : _GEN_6376; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6537 = 8'h85 == total_offset_19 ? field_byte_19 : _GEN_6377; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6538 = 8'h86 == total_offset_19 ? field_byte_19 : _GEN_6378; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6539 = 8'h87 == total_offset_19 ? field_byte_19 : _GEN_6379; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6540 = 8'h88 == total_offset_19 ? field_byte_19 : _GEN_6380; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6541 = 8'h89 == total_offset_19 ? field_byte_19 : _GEN_6381; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6542 = 8'h8a == total_offset_19 ? field_byte_19 : _GEN_6382; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6543 = 8'h8b == total_offset_19 ? field_byte_19 : _GEN_6383; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6544 = 8'h8c == total_offset_19 ? field_byte_19 : _GEN_6384; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6545 = 8'h8d == total_offset_19 ? field_byte_19 : _GEN_6385; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6546 = 8'h8e == total_offset_19 ? field_byte_19 : _GEN_6386; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6547 = 8'h8f == total_offset_19 ? field_byte_19 : _GEN_6387; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6548 = 8'h90 == total_offset_19 ? field_byte_19 : _GEN_6388; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6549 = 8'h91 == total_offset_19 ? field_byte_19 : _GEN_6389; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6550 = 8'h92 == total_offset_19 ? field_byte_19 : _GEN_6390; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6551 = 8'h93 == total_offset_19 ? field_byte_19 : _GEN_6391; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6552 = 8'h94 == total_offset_19 ? field_byte_19 : _GEN_6392; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6553 = 8'h95 == total_offset_19 ? field_byte_19 : _GEN_6393; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6554 = 8'h96 == total_offset_19 ? field_byte_19 : _GEN_6394; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6555 = 8'h97 == total_offset_19 ? field_byte_19 : _GEN_6395; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6556 = 8'h98 == total_offset_19 ? field_byte_19 : _GEN_6396; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6557 = 8'h99 == total_offset_19 ? field_byte_19 : _GEN_6397; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6558 = 8'h9a == total_offset_19 ? field_byte_19 : _GEN_6398; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6559 = 8'h9b == total_offset_19 ? field_byte_19 : _GEN_6399; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6560 = 8'h9c == total_offset_19 ? field_byte_19 : _GEN_6400; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6561 = 8'h9d == total_offset_19 ? field_byte_19 : _GEN_6401; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6562 = 8'h9e == total_offset_19 ? field_byte_19 : _GEN_6402; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6563 = 8'h9f == total_offset_19 ? field_byte_19 : _GEN_6403; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6564 = 8'h3 < length_2 ? _GEN_6404 : _GEN_6244; // @[executor.scala 308:60]
  wire [7:0] _GEN_6565 = 8'h3 < length_2 ? _GEN_6405 : _GEN_6245; // @[executor.scala 308:60]
  wire [7:0] _GEN_6566 = 8'h3 < length_2 ? _GEN_6406 : _GEN_6246; // @[executor.scala 308:60]
  wire [7:0] _GEN_6567 = 8'h3 < length_2 ? _GEN_6407 : _GEN_6247; // @[executor.scala 308:60]
  wire [7:0] _GEN_6568 = 8'h3 < length_2 ? _GEN_6408 : _GEN_6248; // @[executor.scala 308:60]
  wire [7:0] _GEN_6569 = 8'h3 < length_2 ? _GEN_6409 : _GEN_6249; // @[executor.scala 308:60]
  wire [7:0] _GEN_6570 = 8'h3 < length_2 ? _GEN_6410 : _GEN_6250; // @[executor.scala 308:60]
  wire [7:0] _GEN_6571 = 8'h3 < length_2 ? _GEN_6411 : _GEN_6251; // @[executor.scala 308:60]
  wire [7:0] _GEN_6572 = 8'h3 < length_2 ? _GEN_6412 : _GEN_6252; // @[executor.scala 308:60]
  wire [7:0] _GEN_6573 = 8'h3 < length_2 ? _GEN_6413 : _GEN_6253; // @[executor.scala 308:60]
  wire [7:0] _GEN_6574 = 8'h3 < length_2 ? _GEN_6414 : _GEN_6254; // @[executor.scala 308:60]
  wire [7:0] _GEN_6575 = 8'h3 < length_2 ? _GEN_6415 : _GEN_6255; // @[executor.scala 308:60]
  wire [7:0] _GEN_6576 = 8'h3 < length_2 ? _GEN_6416 : _GEN_6256; // @[executor.scala 308:60]
  wire [7:0] _GEN_6577 = 8'h3 < length_2 ? _GEN_6417 : _GEN_6257; // @[executor.scala 308:60]
  wire [7:0] _GEN_6578 = 8'h3 < length_2 ? _GEN_6418 : _GEN_6258; // @[executor.scala 308:60]
  wire [7:0] _GEN_6579 = 8'h3 < length_2 ? _GEN_6419 : _GEN_6259; // @[executor.scala 308:60]
  wire [7:0] _GEN_6580 = 8'h3 < length_2 ? _GEN_6420 : _GEN_6260; // @[executor.scala 308:60]
  wire [7:0] _GEN_6581 = 8'h3 < length_2 ? _GEN_6421 : _GEN_6261; // @[executor.scala 308:60]
  wire [7:0] _GEN_6582 = 8'h3 < length_2 ? _GEN_6422 : _GEN_6262; // @[executor.scala 308:60]
  wire [7:0] _GEN_6583 = 8'h3 < length_2 ? _GEN_6423 : _GEN_6263; // @[executor.scala 308:60]
  wire [7:0] _GEN_6584 = 8'h3 < length_2 ? _GEN_6424 : _GEN_6264; // @[executor.scala 308:60]
  wire [7:0] _GEN_6585 = 8'h3 < length_2 ? _GEN_6425 : _GEN_6265; // @[executor.scala 308:60]
  wire [7:0] _GEN_6586 = 8'h3 < length_2 ? _GEN_6426 : _GEN_6266; // @[executor.scala 308:60]
  wire [7:0] _GEN_6587 = 8'h3 < length_2 ? _GEN_6427 : _GEN_6267; // @[executor.scala 308:60]
  wire [7:0] _GEN_6588 = 8'h3 < length_2 ? _GEN_6428 : _GEN_6268; // @[executor.scala 308:60]
  wire [7:0] _GEN_6589 = 8'h3 < length_2 ? _GEN_6429 : _GEN_6269; // @[executor.scala 308:60]
  wire [7:0] _GEN_6590 = 8'h3 < length_2 ? _GEN_6430 : _GEN_6270; // @[executor.scala 308:60]
  wire [7:0] _GEN_6591 = 8'h3 < length_2 ? _GEN_6431 : _GEN_6271; // @[executor.scala 308:60]
  wire [7:0] _GEN_6592 = 8'h3 < length_2 ? _GEN_6432 : _GEN_6272; // @[executor.scala 308:60]
  wire [7:0] _GEN_6593 = 8'h3 < length_2 ? _GEN_6433 : _GEN_6273; // @[executor.scala 308:60]
  wire [7:0] _GEN_6594 = 8'h3 < length_2 ? _GEN_6434 : _GEN_6274; // @[executor.scala 308:60]
  wire [7:0] _GEN_6595 = 8'h3 < length_2 ? _GEN_6435 : _GEN_6275; // @[executor.scala 308:60]
  wire [7:0] _GEN_6596 = 8'h3 < length_2 ? _GEN_6436 : _GEN_6276; // @[executor.scala 308:60]
  wire [7:0] _GEN_6597 = 8'h3 < length_2 ? _GEN_6437 : _GEN_6277; // @[executor.scala 308:60]
  wire [7:0] _GEN_6598 = 8'h3 < length_2 ? _GEN_6438 : _GEN_6278; // @[executor.scala 308:60]
  wire [7:0] _GEN_6599 = 8'h3 < length_2 ? _GEN_6439 : _GEN_6279; // @[executor.scala 308:60]
  wire [7:0] _GEN_6600 = 8'h3 < length_2 ? _GEN_6440 : _GEN_6280; // @[executor.scala 308:60]
  wire [7:0] _GEN_6601 = 8'h3 < length_2 ? _GEN_6441 : _GEN_6281; // @[executor.scala 308:60]
  wire [7:0] _GEN_6602 = 8'h3 < length_2 ? _GEN_6442 : _GEN_6282; // @[executor.scala 308:60]
  wire [7:0] _GEN_6603 = 8'h3 < length_2 ? _GEN_6443 : _GEN_6283; // @[executor.scala 308:60]
  wire [7:0] _GEN_6604 = 8'h3 < length_2 ? _GEN_6444 : _GEN_6284; // @[executor.scala 308:60]
  wire [7:0] _GEN_6605 = 8'h3 < length_2 ? _GEN_6445 : _GEN_6285; // @[executor.scala 308:60]
  wire [7:0] _GEN_6606 = 8'h3 < length_2 ? _GEN_6446 : _GEN_6286; // @[executor.scala 308:60]
  wire [7:0] _GEN_6607 = 8'h3 < length_2 ? _GEN_6447 : _GEN_6287; // @[executor.scala 308:60]
  wire [7:0] _GEN_6608 = 8'h3 < length_2 ? _GEN_6448 : _GEN_6288; // @[executor.scala 308:60]
  wire [7:0] _GEN_6609 = 8'h3 < length_2 ? _GEN_6449 : _GEN_6289; // @[executor.scala 308:60]
  wire [7:0] _GEN_6610 = 8'h3 < length_2 ? _GEN_6450 : _GEN_6290; // @[executor.scala 308:60]
  wire [7:0] _GEN_6611 = 8'h3 < length_2 ? _GEN_6451 : _GEN_6291; // @[executor.scala 308:60]
  wire [7:0] _GEN_6612 = 8'h3 < length_2 ? _GEN_6452 : _GEN_6292; // @[executor.scala 308:60]
  wire [7:0] _GEN_6613 = 8'h3 < length_2 ? _GEN_6453 : _GEN_6293; // @[executor.scala 308:60]
  wire [7:0] _GEN_6614 = 8'h3 < length_2 ? _GEN_6454 : _GEN_6294; // @[executor.scala 308:60]
  wire [7:0] _GEN_6615 = 8'h3 < length_2 ? _GEN_6455 : _GEN_6295; // @[executor.scala 308:60]
  wire [7:0] _GEN_6616 = 8'h3 < length_2 ? _GEN_6456 : _GEN_6296; // @[executor.scala 308:60]
  wire [7:0] _GEN_6617 = 8'h3 < length_2 ? _GEN_6457 : _GEN_6297; // @[executor.scala 308:60]
  wire [7:0] _GEN_6618 = 8'h3 < length_2 ? _GEN_6458 : _GEN_6298; // @[executor.scala 308:60]
  wire [7:0] _GEN_6619 = 8'h3 < length_2 ? _GEN_6459 : _GEN_6299; // @[executor.scala 308:60]
  wire [7:0] _GEN_6620 = 8'h3 < length_2 ? _GEN_6460 : _GEN_6300; // @[executor.scala 308:60]
  wire [7:0] _GEN_6621 = 8'h3 < length_2 ? _GEN_6461 : _GEN_6301; // @[executor.scala 308:60]
  wire [7:0] _GEN_6622 = 8'h3 < length_2 ? _GEN_6462 : _GEN_6302; // @[executor.scala 308:60]
  wire [7:0] _GEN_6623 = 8'h3 < length_2 ? _GEN_6463 : _GEN_6303; // @[executor.scala 308:60]
  wire [7:0] _GEN_6624 = 8'h3 < length_2 ? _GEN_6464 : _GEN_6304; // @[executor.scala 308:60]
  wire [7:0] _GEN_6625 = 8'h3 < length_2 ? _GEN_6465 : _GEN_6305; // @[executor.scala 308:60]
  wire [7:0] _GEN_6626 = 8'h3 < length_2 ? _GEN_6466 : _GEN_6306; // @[executor.scala 308:60]
  wire [7:0] _GEN_6627 = 8'h3 < length_2 ? _GEN_6467 : _GEN_6307; // @[executor.scala 308:60]
  wire [7:0] _GEN_6628 = 8'h3 < length_2 ? _GEN_6468 : _GEN_6308; // @[executor.scala 308:60]
  wire [7:0] _GEN_6629 = 8'h3 < length_2 ? _GEN_6469 : _GEN_6309; // @[executor.scala 308:60]
  wire [7:0] _GEN_6630 = 8'h3 < length_2 ? _GEN_6470 : _GEN_6310; // @[executor.scala 308:60]
  wire [7:0] _GEN_6631 = 8'h3 < length_2 ? _GEN_6471 : _GEN_6311; // @[executor.scala 308:60]
  wire [7:0] _GEN_6632 = 8'h3 < length_2 ? _GEN_6472 : _GEN_6312; // @[executor.scala 308:60]
  wire [7:0] _GEN_6633 = 8'h3 < length_2 ? _GEN_6473 : _GEN_6313; // @[executor.scala 308:60]
  wire [7:0] _GEN_6634 = 8'h3 < length_2 ? _GEN_6474 : _GEN_6314; // @[executor.scala 308:60]
  wire [7:0] _GEN_6635 = 8'h3 < length_2 ? _GEN_6475 : _GEN_6315; // @[executor.scala 308:60]
  wire [7:0] _GEN_6636 = 8'h3 < length_2 ? _GEN_6476 : _GEN_6316; // @[executor.scala 308:60]
  wire [7:0] _GEN_6637 = 8'h3 < length_2 ? _GEN_6477 : _GEN_6317; // @[executor.scala 308:60]
  wire [7:0] _GEN_6638 = 8'h3 < length_2 ? _GEN_6478 : _GEN_6318; // @[executor.scala 308:60]
  wire [7:0] _GEN_6639 = 8'h3 < length_2 ? _GEN_6479 : _GEN_6319; // @[executor.scala 308:60]
  wire [7:0] _GEN_6640 = 8'h3 < length_2 ? _GEN_6480 : _GEN_6320; // @[executor.scala 308:60]
  wire [7:0] _GEN_6641 = 8'h3 < length_2 ? _GEN_6481 : _GEN_6321; // @[executor.scala 308:60]
  wire [7:0] _GEN_6642 = 8'h3 < length_2 ? _GEN_6482 : _GEN_6322; // @[executor.scala 308:60]
  wire [7:0] _GEN_6643 = 8'h3 < length_2 ? _GEN_6483 : _GEN_6323; // @[executor.scala 308:60]
  wire [7:0] _GEN_6644 = 8'h3 < length_2 ? _GEN_6484 : _GEN_6324; // @[executor.scala 308:60]
  wire [7:0] _GEN_6645 = 8'h3 < length_2 ? _GEN_6485 : _GEN_6325; // @[executor.scala 308:60]
  wire [7:0] _GEN_6646 = 8'h3 < length_2 ? _GEN_6486 : _GEN_6326; // @[executor.scala 308:60]
  wire [7:0] _GEN_6647 = 8'h3 < length_2 ? _GEN_6487 : _GEN_6327; // @[executor.scala 308:60]
  wire [7:0] _GEN_6648 = 8'h3 < length_2 ? _GEN_6488 : _GEN_6328; // @[executor.scala 308:60]
  wire [7:0] _GEN_6649 = 8'h3 < length_2 ? _GEN_6489 : _GEN_6329; // @[executor.scala 308:60]
  wire [7:0] _GEN_6650 = 8'h3 < length_2 ? _GEN_6490 : _GEN_6330; // @[executor.scala 308:60]
  wire [7:0] _GEN_6651 = 8'h3 < length_2 ? _GEN_6491 : _GEN_6331; // @[executor.scala 308:60]
  wire [7:0] _GEN_6652 = 8'h3 < length_2 ? _GEN_6492 : _GEN_6332; // @[executor.scala 308:60]
  wire [7:0] _GEN_6653 = 8'h3 < length_2 ? _GEN_6493 : _GEN_6333; // @[executor.scala 308:60]
  wire [7:0] _GEN_6654 = 8'h3 < length_2 ? _GEN_6494 : _GEN_6334; // @[executor.scala 308:60]
  wire [7:0] _GEN_6655 = 8'h3 < length_2 ? _GEN_6495 : _GEN_6335; // @[executor.scala 308:60]
  wire [7:0] _GEN_6656 = 8'h3 < length_2 ? _GEN_6496 : _GEN_6336; // @[executor.scala 308:60]
  wire [7:0] _GEN_6657 = 8'h3 < length_2 ? _GEN_6497 : _GEN_6337; // @[executor.scala 308:60]
  wire [7:0] _GEN_6658 = 8'h3 < length_2 ? _GEN_6498 : _GEN_6338; // @[executor.scala 308:60]
  wire [7:0] _GEN_6659 = 8'h3 < length_2 ? _GEN_6499 : _GEN_6339; // @[executor.scala 308:60]
  wire [7:0] _GEN_6660 = 8'h3 < length_2 ? _GEN_6500 : _GEN_6340; // @[executor.scala 308:60]
  wire [7:0] _GEN_6661 = 8'h3 < length_2 ? _GEN_6501 : _GEN_6341; // @[executor.scala 308:60]
  wire [7:0] _GEN_6662 = 8'h3 < length_2 ? _GEN_6502 : _GEN_6342; // @[executor.scala 308:60]
  wire [7:0] _GEN_6663 = 8'h3 < length_2 ? _GEN_6503 : _GEN_6343; // @[executor.scala 308:60]
  wire [7:0] _GEN_6664 = 8'h3 < length_2 ? _GEN_6504 : _GEN_6344; // @[executor.scala 308:60]
  wire [7:0] _GEN_6665 = 8'h3 < length_2 ? _GEN_6505 : _GEN_6345; // @[executor.scala 308:60]
  wire [7:0] _GEN_6666 = 8'h3 < length_2 ? _GEN_6506 : _GEN_6346; // @[executor.scala 308:60]
  wire [7:0] _GEN_6667 = 8'h3 < length_2 ? _GEN_6507 : _GEN_6347; // @[executor.scala 308:60]
  wire [7:0] _GEN_6668 = 8'h3 < length_2 ? _GEN_6508 : _GEN_6348; // @[executor.scala 308:60]
  wire [7:0] _GEN_6669 = 8'h3 < length_2 ? _GEN_6509 : _GEN_6349; // @[executor.scala 308:60]
  wire [7:0] _GEN_6670 = 8'h3 < length_2 ? _GEN_6510 : _GEN_6350; // @[executor.scala 308:60]
  wire [7:0] _GEN_6671 = 8'h3 < length_2 ? _GEN_6511 : _GEN_6351; // @[executor.scala 308:60]
  wire [7:0] _GEN_6672 = 8'h3 < length_2 ? _GEN_6512 : _GEN_6352; // @[executor.scala 308:60]
  wire [7:0] _GEN_6673 = 8'h3 < length_2 ? _GEN_6513 : _GEN_6353; // @[executor.scala 308:60]
  wire [7:0] _GEN_6674 = 8'h3 < length_2 ? _GEN_6514 : _GEN_6354; // @[executor.scala 308:60]
  wire [7:0] _GEN_6675 = 8'h3 < length_2 ? _GEN_6515 : _GEN_6355; // @[executor.scala 308:60]
  wire [7:0] _GEN_6676 = 8'h3 < length_2 ? _GEN_6516 : _GEN_6356; // @[executor.scala 308:60]
  wire [7:0] _GEN_6677 = 8'h3 < length_2 ? _GEN_6517 : _GEN_6357; // @[executor.scala 308:60]
  wire [7:0] _GEN_6678 = 8'h3 < length_2 ? _GEN_6518 : _GEN_6358; // @[executor.scala 308:60]
  wire [7:0] _GEN_6679 = 8'h3 < length_2 ? _GEN_6519 : _GEN_6359; // @[executor.scala 308:60]
  wire [7:0] _GEN_6680 = 8'h3 < length_2 ? _GEN_6520 : _GEN_6360; // @[executor.scala 308:60]
  wire [7:0] _GEN_6681 = 8'h3 < length_2 ? _GEN_6521 : _GEN_6361; // @[executor.scala 308:60]
  wire [7:0] _GEN_6682 = 8'h3 < length_2 ? _GEN_6522 : _GEN_6362; // @[executor.scala 308:60]
  wire [7:0] _GEN_6683 = 8'h3 < length_2 ? _GEN_6523 : _GEN_6363; // @[executor.scala 308:60]
  wire [7:0] _GEN_6684 = 8'h3 < length_2 ? _GEN_6524 : _GEN_6364; // @[executor.scala 308:60]
  wire [7:0] _GEN_6685 = 8'h3 < length_2 ? _GEN_6525 : _GEN_6365; // @[executor.scala 308:60]
  wire [7:0] _GEN_6686 = 8'h3 < length_2 ? _GEN_6526 : _GEN_6366; // @[executor.scala 308:60]
  wire [7:0] _GEN_6687 = 8'h3 < length_2 ? _GEN_6527 : _GEN_6367; // @[executor.scala 308:60]
  wire [7:0] _GEN_6688 = 8'h3 < length_2 ? _GEN_6528 : _GEN_6368; // @[executor.scala 308:60]
  wire [7:0] _GEN_6689 = 8'h3 < length_2 ? _GEN_6529 : _GEN_6369; // @[executor.scala 308:60]
  wire [7:0] _GEN_6690 = 8'h3 < length_2 ? _GEN_6530 : _GEN_6370; // @[executor.scala 308:60]
  wire [7:0] _GEN_6691 = 8'h3 < length_2 ? _GEN_6531 : _GEN_6371; // @[executor.scala 308:60]
  wire [7:0] _GEN_6692 = 8'h3 < length_2 ? _GEN_6532 : _GEN_6372; // @[executor.scala 308:60]
  wire [7:0] _GEN_6693 = 8'h3 < length_2 ? _GEN_6533 : _GEN_6373; // @[executor.scala 308:60]
  wire [7:0] _GEN_6694 = 8'h3 < length_2 ? _GEN_6534 : _GEN_6374; // @[executor.scala 308:60]
  wire [7:0] _GEN_6695 = 8'h3 < length_2 ? _GEN_6535 : _GEN_6375; // @[executor.scala 308:60]
  wire [7:0] _GEN_6696 = 8'h3 < length_2 ? _GEN_6536 : _GEN_6376; // @[executor.scala 308:60]
  wire [7:0] _GEN_6697 = 8'h3 < length_2 ? _GEN_6537 : _GEN_6377; // @[executor.scala 308:60]
  wire [7:0] _GEN_6698 = 8'h3 < length_2 ? _GEN_6538 : _GEN_6378; // @[executor.scala 308:60]
  wire [7:0] _GEN_6699 = 8'h3 < length_2 ? _GEN_6539 : _GEN_6379; // @[executor.scala 308:60]
  wire [7:0] _GEN_6700 = 8'h3 < length_2 ? _GEN_6540 : _GEN_6380; // @[executor.scala 308:60]
  wire [7:0] _GEN_6701 = 8'h3 < length_2 ? _GEN_6541 : _GEN_6381; // @[executor.scala 308:60]
  wire [7:0] _GEN_6702 = 8'h3 < length_2 ? _GEN_6542 : _GEN_6382; // @[executor.scala 308:60]
  wire [7:0] _GEN_6703 = 8'h3 < length_2 ? _GEN_6543 : _GEN_6383; // @[executor.scala 308:60]
  wire [7:0] _GEN_6704 = 8'h3 < length_2 ? _GEN_6544 : _GEN_6384; // @[executor.scala 308:60]
  wire [7:0] _GEN_6705 = 8'h3 < length_2 ? _GEN_6545 : _GEN_6385; // @[executor.scala 308:60]
  wire [7:0] _GEN_6706 = 8'h3 < length_2 ? _GEN_6546 : _GEN_6386; // @[executor.scala 308:60]
  wire [7:0] _GEN_6707 = 8'h3 < length_2 ? _GEN_6547 : _GEN_6387; // @[executor.scala 308:60]
  wire [7:0] _GEN_6708 = 8'h3 < length_2 ? _GEN_6548 : _GEN_6388; // @[executor.scala 308:60]
  wire [7:0] _GEN_6709 = 8'h3 < length_2 ? _GEN_6549 : _GEN_6389; // @[executor.scala 308:60]
  wire [7:0] _GEN_6710 = 8'h3 < length_2 ? _GEN_6550 : _GEN_6390; // @[executor.scala 308:60]
  wire [7:0] _GEN_6711 = 8'h3 < length_2 ? _GEN_6551 : _GEN_6391; // @[executor.scala 308:60]
  wire [7:0] _GEN_6712 = 8'h3 < length_2 ? _GEN_6552 : _GEN_6392; // @[executor.scala 308:60]
  wire [7:0] _GEN_6713 = 8'h3 < length_2 ? _GEN_6553 : _GEN_6393; // @[executor.scala 308:60]
  wire [7:0] _GEN_6714 = 8'h3 < length_2 ? _GEN_6554 : _GEN_6394; // @[executor.scala 308:60]
  wire [7:0] _GEN_6715 = 8'h3 < length_2 ? _GEN_6555 : _GEN_6395; // @[executor.scala 308:60]
  wire [7:0] _GEN_6716 = 8'h3 < length_2 ? _GEN_6556 : _GEN_6396; // @[executor.scala 308:60]
  wire [7:0] _GEN_6717 = 8'h3 < length_2 ? _GEN_6557 : _GEN_6397; // @[executor.scala 308:60]
  wire [7:0] _GEN_6718 = 8'h3 < length_2 ? _GEN_6558 : _GEN_6398; // @[executor.scala 308:60]
  wire [7:0] _GEN_6719 = 8'h3 < length_2 ? _GEN_6559 : _GEN_6399; // @[executor.scala 308:60]
  wire [7:0] _GEN_6720 = 8'h3 < length_2 ? _GEN_6560 : _GEN_6400; // @[executor.scala 308:60]
  wire [7:0] _GEN_6721 = 8'h3 < length_2 ? _GEN_6561 : _GEN_6401; // @[executor.scala 308:60]
  wire [7:0] _GEN_6722 = 8'h3 < length_2 ? _GEN_6562 : _GEN_6402; // @[executor.scala 308:60]
  wire [7:0] _GEN_6723 = 8'h3 < length_2 ? _GEN_6563 : _GEN_6403; // @[executor.scala 308:60]
  wire [7:0] field_byte_20 = field_2[31:24]; // @[executor.scala 305:57]
  wire [7:0] total_offset_20 = offset_2 + 8'h4; // @[executor.scala 307:57]
  wire [7:0] _GEN_6724 = 8'h0 == total_offset_20 ? field_byte_20 : _GEN_6564; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6725 = 8'h1 == total_offset_20 ? field_byte_20 : _GEN_6565; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6726 = 8'h2 == total_offset_20 ? field_byte_20 : _GEN_6566; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6727 = 8'h3 == total_offset_20 ? field_byte_20 : _GEN_6567; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6728 = 8'h4 == total_offset_20 ? field_byte_20 : _GEN_6568; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6729 = 8'h5 == total_offset_20 ? field_byte_20 : _GEN_6569; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6730 = 8'h6 == total_offset_20 ? field_byte_20 : _GEN_6570; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6731 = 8'h7 == total_offset_20 ? field_byte_20 : _GEN_6571; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6732 = 8'h8 == total_offset_20 ? field_byte_20 : _GEN_6572; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6733 = 8'h9 == total_offset_20 ? field_byte_20 : _GEN_6573; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6734 = 8'ha == total_offset_20 ? field_byte_20 : _GEN_6574; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6735 = 8'hb == total_offset_20 ? field_byte_20 : _GEN_6575; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6736 = 8'hc == total_offset_20 ? field_byte_20 : _GEN_6576; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6737 = 8'hd == total_offset_20 ? field_byte_20 : _GEN_6577; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6738 = 8'he == total_offset_20 ? field_byte_20 : _GEN_6578; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6739 = 8'hf == total_offset_20 ? field_byte_20 : _GEN_6579; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6740 = 8'h10 == total_offset_20 ? field_byte_20 : _GEN_6580; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6741 = 8'h11 == total_offset_20 ? field_byte_20 : _GEN_6581; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6742 = 8'h12 == total_offset_20 ? field_byte_20 : _GEN_6582; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6743 = 8'h13 == total_offset_20 ? field_byte_20 : _GEN_6583; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6744 = 8'h14 == total_offset_20 ? field_byte_20 : _GEN_6584; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6745 = 8'h15 == total_offset_20 ? field_byte_20 : _GEN_6585; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6746 = 8'h16 == total_offset_20 ? field_byte_20 : _GEN_6586; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6747 = 8'h17 == total_offset_20 ? field_byte_20 : _GEN_6587; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6748 = 8'h18 == total_offset_20 ? field_byte_20 : _GEN_6588; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6749 = 8'h19 == total_offset_20 ? field_byte_20 : _GEN_6589; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6750 = 8'h1a == total_offset_20 ? field_byte_20 : _GEN_6590; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6751 = 8'h1b == total_offset_20 ? field_byte_20 : _GEN_6591; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6752 = 8'h1c == total_offset_20 ? field_byte_20 : _GEN_6592; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6753 = 8'h1d == total_offset_20 ? field_byte_20 : _GEN_6593; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6754 = 8'h1e == total_offset_20 ? field_byte_20 : _GEN_6594; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6755 = 8'h1f == total_offset_20 ? field_byte_20 : _GEN_6595; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6756 = 8'h20 == total_offset_20 ? field_byte_20 : _GEN_6596; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6757 = 8'h21 == total_offset_20 ? field_byte_20 : _GEN_6597; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6758 = 8'h22 == total_offset_20 ? field_byte_20 : _GEN_6598; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6759 = 8'h23 == total_offset_20 ? field_byte_20 : _GEN_6599; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6760 = 8'h24 == total_offset_20 ? field_byte_20 : _GEN_6600; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6761 = 8'h25 == total_offset_20 ? field_byte_20 : _GEN_6601; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6762 = 8'h26 == total_offset_20 ? field_byte_20 : _GEN_6602; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6763 = 8'h27 == total_offset_20 ? field_byte_20 : _GEN_6603; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6764 = 8'h28 == total_offset_20 ? field_byte_20 : _GEN_6604; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6765 = 8'h29 == total_offset_20 ? field_byte_20 : _GEN_6605; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6766 = 8'h2a == total_offset_20 ? field_byte_20 : _GEN_6606; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6767 = 8'h2b == total_offset_20 ? field_byte_20 : _GEN_6607; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6768 = 8'h2c == total_offset_20 ? field_byte_20 : _GEN_6608; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6769 = 8'h2d == total_offset_20 ? field_byte_20 : _GEN_6609; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6770 = 8'h2e == total_offset_20 ? field_byte_20 : _GEN_6610; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6771 = 8'h2f == total_offset_20 ? field_byte_20 : _GEN_6611; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6772 = 8'h30 == total_offset_20 ? field_byte_20 : _GEN_6612; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6773 = 8'h31 == total_offset_20 ? field_byte_20 : _GEN_6613; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6774 = 8'h32 == total_offset_20 ? field_byte_20 : _GEN_6614; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6775 = 8'h33 == total_offset_20 ? field_byte_20 : _GEN_6615; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6776 = 8'h34 == total_offset_20 ? field_byte_20 : _GEN_6616; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6777 = 8'h35 == total_offset_20 ? field_byte_20 : _GEN_6617; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6778 = 8'h36 == total_offset_20 ? field_byte_20 : _GEN_6618; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6779 = 8'h37 == total_offset_20 ? field_byte_20 : _GEN_6619; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6780 = 8'h38 == total_offset_20 ? field_byte_20 : _GEN_6620; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6781 = 8'h39 == total_offset_20 ? field_byte_20 : _GEN_6621; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6782 = 8'h3a == total_offset_20 ? field_byte_20 : _GEN_6622; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6783 = 8'h3b == total_offset_20 ? field_byte_20 : _GEN_6623; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6784 = 8'h3c == total_offset_20 ? field_byte_20 : _GEN_6624; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6785 = 8'h3d == total_offset_20 ? field_byte_20 : _GEN_6625; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6786 = 8'h3e == total_offset_20 ? field_byte_20 : _GEN_6626; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6787 = 8'h3f == total_offset_20 ? field_byte_20 : _GEN_6627; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6788 = 8'h40 == total_offset_20 ? field_byte_20 : _GEN_6628; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6789 = 8'h41 == total_offset_20 ? field_byte_20 : _GEN_6629; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6790 = 8'h42 == total_offset_20 ? field_byte_20 : _GEN_6630; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6791 = 8'h43 == total_offset_20 ? field_byte_20 : _GEN_6631; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6792 = 8'h44 == total_offset_20 ? field_byte_20 : _GEN_6632; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6793 = 8'h45 == total_offset_20 ? field_byte_20 : _GEN_6633; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6794 = 8'h46 == total_offset_20 ? field_byte_20 : _GEN_6634; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6795 = 8'h47 == total_offset_20 ? field_byte_20 : _GEN_6635; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6796 = 8'h48 == total_offset_20 ? field_byte_20 : _GEN_6636; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6797 = 8'h49 == total_offset_20 ? field_byte_20 : _GEN_6637; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6798 = 8'h4a == total_offset_20 ? field_byte_20 : _GEN_6638; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6799 = 8'h4b == total_offset_20 ? field_byte_20 : _GEN_6639; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6800 = 8'h4c == total_offset_20 ? field_byte_20 : _GEN_6640; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6801 = 8'h4d == total_offset_20 ? field_byte_20 : _GEN_6641; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6802 = 8'h4e == total_offset_20 ? field_byte_20 : _GEN_6642; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6803 = 8'h4f == total_offset_20 ? field_byte_20 : _GEN_6643; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6804 = 8'h50 == total_offset_20 ? field_byte_20 : _GEN_6644; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6805 = 8'h51 == total_offset_20 ? field_byte_20 : _GEN_6645; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6806 = 8'h52 == total_offset_20 ? field_byte_20 : _GEN_6646; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6807 = 8'h53 == total_offset_20 ? field_byte_20 : _GEN_6647; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6808 = 8'h54 == total_offset_20 ? field_byte_20 : _GEN_6648; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6809 = 8'h55 == total_offset_20 ? field_byte_20 : _GEN_6649; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6810 = 8'h56 == total_offset_20 ? field_byte_20 : _GEN_6650; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6811 = 8'h57 == total_offset_20 ? field_byte_20 : _GEN_6651; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6812 = 8'h58 == total_offset_20 ? field_byte_20 : _GEN_6652; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6813 = 8'h59 == total_offset_20 ? field_byte_20 : _GEN_6653; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6814 = 8'h5a == total_offset_20 ? field_byte_20 : _GEN_6654; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6815 = 8'h5b == total_offset_20 ? field_byte_20 : _GEN_6655; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6816 = 8'h5c == total_offset_20 ? field_byte_20 : _GEN_6656; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6817 = 8'h5d == total_offset_20 ? field_byte_20 : _GEN_6657; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6818 = 8'h5e == total_offset_20 ? field_byte_20 : _GEN_6658; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6819 = 8'h5f == total_offset_20 ? field_byte_20 : _GEN_6659; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6820 = 8'h60 == total_offset_20 ? field_byte_20 : _GEN_6660; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6821 = 8'h61 == total_offset_20 ? field_byte_20 : _GEN_6661; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6822 = 8'h62 == total_offset_20 ? field_byte_20 : _GEN_6662; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6823 = 8'h63 == total_offset_20 ? field_byte_20 : _GEN_6663; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6824 = 8'h64 == total_offset_20 ? field_byte_20 : _GEN_6664; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6825 = 8'h65 == total_offset_20 ? field_byte_20 : _GEN_6665; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6826 = 8'h66 == total_offset_20 ? field_byte_20 : _GEN_6666; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6827 = 8'h67 == total_offset_20 ? field_byte_20 : _GEN_6667; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6828 = 8'h68 == total_offset_20 ? field_byte_20 : _GEN_6668; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6829 = 8'h69 == total_offset_20 ? field_byte_20 : _GEN_6669; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6830 = 8'h6a == total_offset_20 ? field_byte_20 : _GEN_6670; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6831 = 8'h6b == total_offset_20 ? field_byte_20 : _GEN_6671; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6832 = 8'h6c == total_offset_20 ? field_byte_20 : _GEN_6672; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6833 = 8'h6d == total_offset_20 ? field_byte_20 : _GEN_6673; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6834 = 8'h6e == total_offset_20 ? field_byte_20 : _GEN_6674; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6835 = 8'h6f == total_offset_20 ? field_byte_20 : _GEN_6675; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6836 = 8'h70 == total_offset_20 ? field_byte_20 : _GEN_6676; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6837 = 8'h71 == total_offset_20 ? field_byte_20 : _GEN_6677; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6838 = 8'h72 == total_offset_20 ? field_byte_20 : _GEN_6678; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6839 = 8'h73 == total_offset_20 ? field_byte_20 : _GEN_6679; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6840 = 8'h74 == total_offset_20 ? field_byte_20 : _GEN_6680; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6841 = 8'h75 == total_offset_20 ? field_byte_20 : _GEN_6681; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6842 = 8'h76 == total_offset_20 ? field_byte_20 : _GEN_6682; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6843 = 8'h77 == total_offset_20 ? field_byte_20 : _GEN_6683; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6844 = 8'h78 == total_offset_20 ? field_byte_20 : _GEN_6684; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6845 = 8'h79 == total_offset_20 ? field_byte_20 : _GEN_6685; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6846 = 8'h7a == total_offset_20 ? field_byte_20 : _GEN_6686; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6847 = 8'h7b == total_offset_20 ? field_byte_20 : _GEN_6687; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6848 = 8'h7c == total_offset_20 ? field_byte_20 : _GEN_6688; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6849 = 8'h7d == total_offset_20 ? field_byte_20 : _GEN_6689; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6850 = 8'h7e == total_offset_20 ? field_byte_20 : _GEN_6690; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6851 = 8'h7f == total_offset_20 ? field_byte_20 : _GEN_6691; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6852 = 8'h80 == total_offset_20 ? field_byte_20 : _GEN_6692; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6853 = 8'h81 == total_offset_20 ? field_byte_20 : _GEN_6693; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6854 = 8'h82 == total_offset_20 ? field_byte_20 : _GEN_6694; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6855 = 8'h83 == total_offset_20 ? field_byte_20 : _GEN_6695; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6856 = 8'h84 == total_offset_20 ? field_byte_20 : _GEN_6696; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6857 = 8'h85 == total_offset_20 ? field_byte_20 : _GEN_6697; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6858 = 8'h86 == total_offset_20 ? field_byte_20 : _GEN_6698; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6859 = 8'h87 == total_offset_20 ? field_byte_20 : _GEN_6699; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6860 = 8'h88 == total_offset_20 ? field_byte_20 : _GEN_6700; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6861 = 8'h89 == total_offset_20 ? field_byte_20 : _GEN_6701; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6862 = 8'h8a == total_offset_20 ? field_byte_20 : _GEN_6702; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6863 = 8'h8b == total_offset_20 ? field_byte_20 : _GEN_6703; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6864 = 8'h8c == total_offset_20 ? field_byte_20 : _GEN_6704; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6865 = 8'h8d == total_offset_20 ? field_byte_20 : _GEN_6705; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6866 = 8'h8e == total_offset_20 ? field_byte_20 : _GEN_6706; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6867 = 8'h8f == total_offset_20 ? field_byte_20 : _GEN_6707; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6868 = 8'h90 == total_offset_20 ? field_byte_20 : _GEN_6708; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6869 = 8'h91 == total_offset_20 ? field_byte_20 : _GEN_6709; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6870 = 8'h92 == total_offset_20 ? field_byte_20 : _GEN_6710; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6871 = 8'h93 == total_offset_20 ? field_byte_20 : _GEN_6711; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6872 = 8'h94 == total_offset_20 ? field_byte_20 : _GEN_6712; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6873 = 8'h95 == total_offset_20 ? field_byte_20 : _GEN_6713; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6874 = 8'h96 == total_offset_20 ? field_byte_20 : _GEN_6714; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6875 = 8'h97 == total_offset_20 ? field_byte_20 : _GEN_6715; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6876 = 8'h98 == total_offset_20 ? field_byte_20 : _GEN_6716; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6877 = 8'h99 == total_offset_20 ? field_byte_20 : _GEN_6717; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6878 = 8'h9a == total_offset_20 ? field_byte_20 : _GEN_6718; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6879 = 8'h9b == total_offset_20 ? field_byte_20 : _GEN_6719; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6880 = 8'h9c == total_offset_20 ? field_byte_20 : _GEN_6720; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6881 = 8'h9d == total_offset_20 ? field_byte_20 : _GEN_6721; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6882 = 8'h9e == total_offset_20 ? field_byte_20 : _GEN_6722; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6883 = 8'h9f == total_offset_20 ? field_byte_20 : _GEN_6723; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_6884 = 8'h4 < length_2 ? _GEN_6724 : _GEN_6564; // @[executor.scala 308:60]
  wire [7:0] _GEN_6885 = 8'h4 < length_2 ? _GEN_6725 : _GEN_6565; // @[executor.scala 308:60]
  wire [7:0] _GEN_6886 = 8'h4 < length_2 ? _GEN_6726 : _GEN_6566; // @[executor.scala 308:60]
  wire [7:0] _GEN_6887 = 8'h4 < length_2 ? _GEN_6727 : _GEN_6567; // @[executor.scala 308:60]
  wire [7:0] _GEN_6888 = 8'h4 < length_2 ? _GEN_6728 : _GEN_6568; // @[executor.scala 308:60]
  wire [7:0] _GEN_6889 = 8'h4 < length_2 ? _GEN_6729 : _GEN_6569; // @[executor.scala 308:60]
  wire [7:0] _GEN_6890 = 8'h4 < length_2 ? _GEN_6730 : _GEN_6570; // @[executor.scala 308:60]
  wire [7:0] _GEN_6891 = 8'h4 < length_2 ? _GEN_6731 : _GEN_6571; // @[executor.scala 308:60]
  wire [7:0] _GEN_6892 = 8'h4 < length_2 ? _GEN_6732 : _GEN_6572; // @[executor.scala 308:60]
  wire [7:0] _GEN_6893 = 8'h4 < length_2 ? _GEN_6733 : _GEN_6573; // @[executor.scala 308:60]
  wire [7:0] _GEN_6894 = 8'h4 < length_2 ? _GEN_6734 : _GEN_6574; // @[executor.scala 308:60]
  wire [7:0] _GEN_6895 = 8'h4 < length_2 ? _GEN_6735 : _GEN_6575; // @[executor.scala 308:60]
  wire [7:0] _GEN_6896 = 8'h4 < length_2 ? _GEN_6736 : _GEN_6576; // @[executor.scala 308:60]
  wire [7:0] _GEN_6897 = 8'h4 < length_2 ? _GEN_6737 : _GEN_6577; // @[executor.scala 308:60]
  wire [7:0] _GEN_6898 = 8'h4 < length_2 ? _GEN_6738 : _GEN_6578; // @[executor.scala 308:60]
  wire [7:0] _GEN_6899 = 8'h4 < length_2 ? _GEN_6739 : _GEN_6579; // @[executor.scala 308:60]
  wire [7:0] _GEN_6900 = 8'h4 < length_2 ? _GEN_6740 : _GEN_6580; // @[executor.scala 308:60]
  wire [7:0] _GEN_6901 = 8'h4 < length_2 ? _GEN_6741 : _GEN_6581; // @[executor.scala 308:60]
  wire [7:0] _GEN_6902 = 8'h4 < length_2 ? _GEN_6742 : _GEN_6582; // @[executor.scala 308:60]
  wire [7:0] _GEN_6903 = 8'h4 < length_2 ? _GEN_6743 : _GEN_6583; // @[executor.scala 308:60]
  wire [7:0] _GEN_6904 = 8'h4 < length_2 ? _GEN_6744 : _GEN_6584; // @[executor.scala 308:60]
  wire [7:0] _GEN_6905 = 8'h4 < length_2 ? _GEN_6745 : _GEN_6585; // @[executor.scala 308:60]
  wire [7:0] _GEN_6906 = 8'h4 < length_2 ? _GEN_6746 : _GEN_6586; // @[executor.scala 308:60]
  wire [7:0] _GEN_6907 = 8'h4 < length_2 ? _GEN_6747 : _GEN_6587; // @[executor.scala 308:60]
  wire [7:0] _GEN_6908 = 8'h4 < length_2 ? _GEN_6748 : _GEN_6588; // @[executor.scala 308:60]
  wire [7:0] _GEN_6909 = 8'h4 < length_2 ? _GEN_6749 : _GEN_6589; // @[executor.scala 308:60]
  wire [7:0] _GEN_6910 = 8'h4 < length_2 ? _GEN_6750 : _GEN_6590; // @[executor.scala 308:60]
  wire [7:0] _GEN_6911 = 8'h4 < length_2 ? _GEN_6751 : _GEN_6591; // @[executor.scala 308:60]
  wire [7:0] _GEN_6912 = 8'h4 < length_2 ? _GEN_6752 : _GEN_6592; // @[executor.scala 308:60]
  wire [7:0] _GEN_6913 = 8'h4 < length_2 ? _GEN_6753 : _GEN_6593; // @[executor.scala 308:60]
  wire [7:0] _GEN_6914 = 8'h4 < length_2 ? _GEN_6754 : _GEN_6594; // @[executor.scala 308:60]
  wire [7:0] _GEN_6915 = 8'h4 < length_2 ? _GEN_6755 : _GEN_6595; // @[executor.scala 308:60]
  wire [7:0] _GEN_6916 = 8'h4 < length_2 ? _GEN_6756 : _GEN_6596; // @[executor.scala 308:60]
  wire [7:0] _GEN_6917 = 8'h4 < length_2 ? _GEN_6757 : _GEN_6597; // @[executor.scala 308:60]
  wire [7:0] _GEN_6918 = 8'h4 < length_2 ? _GEN_6758 : _GEN_6598; // @[executor.scala 308:60]
  wire [7:0] _GEN_6919 = 8'h4 < length_2 ? _GEN_6759 : _GEN_6599; // @[executor.scala 308:60]
  wire [7:0] _GEN_6920 = 8'h4 < length_2 ? _GEN_6760 : _GEN_6600; // @[executor.scala 308:60]
  wire [7:0] _GEN_6921 = 8'h4 < length_2 ? _GEN_6761 : _GEN_6601; // @[executor.scala 308:60]
  wire [7:0] _GEN_6922 = 8'h4 < length_2 ? _GEN_6762 : _GEN_6602; // @[executor.scala 308:60]
  wire [7:0] _GEN_6923 = 8'h4 < length_2 ? _GEN_6763 : _GEN_6603; // @[executor.scala 308:60]
  wire [7:0] _GEN_6924 = 8'h4 < length_2 ? _GEN_6764 : _GEN_6604; // @[executor.scala 308:60]
  wire [7:0] _GEN_6925 = 8'h4 < length_2 ? _GEN_6765 : _GEN_6605; // @[executor.scala 308:60]
  wire [7:0] _GEN_6926 = 8'h4 < length_2 ? _GEN_6766 : _GEN_6606; // @[executor.scala 308:60]
  wire [7:0] _GEN_6927 = 8'h4 < length_2 ? _GEN_6767 : _GEN_6607; // @[executor.scala 308:60]
  wire [7:0] _GEN_6928 = 8'h4 < length_2 ? _GEN_6768 : _GEN_6608; // @[executor.scala 308:60]
  wire [7:0] _GEN_6929 = 8'h4 < length_2 ? _GEN_6769 : _GEN_6609; // @[executor.scala 308:60]
  wire [7:0] _GEN_6930 = 8'h4 < length_2 ? _GEN_6770 : _GEN_6610; // @[executor.scala 308:60]
  wire [7:0] _GEN_6931 = 8'h4 < length_2 ? _GEN_6771 : _GEN_6611; // @[executor.scala 308:60]
  wire [7:0] _GEN_6932 = 8'h4 < length_2 ? _GEN_6772 : _GEN_6612; // @[executor.scala 308:60]
  wire [7:0] _GEN_6933 = 8'h4 < length_2 ? _GEN_6773 : _GEN_6613; // @[executor.scala 308:60]
  wire [7:0] _GEN_6934 = 8'h4 < length_2 ? _GEN_6774 : _GEN_6614; // @[executor.scala 308:60]
  wire [7:0] _GEN_6935 = 8'h4 < length_2 ? _GEN_6775 : _GEN_6615; // @[executor.scala 308:60]
  wire [7:0] _GEN_6936 = 8'h4 < length_2 ? _GEN_6776 : _GEN_6616; // @[executor.scala 308:60]
  wire [7:0] _GEN_6937 = 8'h4 < length_2 ? _GEN_6777 : _GEN_6617; // @[executor.scala 308:60]
  wire [7:0] _GEN_6938 = 8'h4 < length_2 ? _GEN_6778 : _GEN_6618; // @[executor.scala 308:60]
  wire [7:0] _GEN_6939 = 8'h4 < length_2 ? _GEN_6779 : _GEN_6619; // @[executor.scala 308:60]
  wire [7:0] _GEN_6940 = 8'h4 < length_2 ? _GEN_6780 : _GEN_6620; // @[executor.scala 308:60]
  wire [7:0] _GEN_6941 = 8'h4 < length_2 ? _GEN_6781 : _GEN_6621; // @[executor.scala 308:60]
  wire [7:0] _GEN_6942 = 8'h4 < length_2 ? _GEN_6782 : _GEN_6622; // @[executor.scala 308:60]
  wire [7:0] _GEN_6943 = 8'h4 < length_2 ? _GEN_6783 : _GEN_6623; // @[executor.scala 308:60]
  wire [7:0] _GEN_6944 = 8'h4 < length_2 ? _GEN_6784 : _GEN_6624; // @[executor.scala 308:60]
  wire [7:0] _GEN_6945 = 8'h4 < length_2 ? _GEN_6785 : _GEN_6625; // @[executor.scala 308:60]
  wire [7:0] _GEN_6946 = 8'h4 < length_2 ? _GEN_6786 : _GEN_6626; // @[executor.scala 308:60]
  wire [7:0] _GEN_6947 = 8'h4 < length_2 ? _GEN_6787 : _GEN_6627; // @[executor.scala 308:60]
  wire [7:0] _GEN_6948 = 8'h4 < length_2 ? _GEN_6788 : _GEN_6628; // @[executor.scala 308:60]
  wire [7:0] _GEN_6949 = 8'h4 < length_2 ? _GEN_6789 : _GEN_6629; // @[executor.scala 308:60]
  wire [7:0] _GEN_6950 = 8'h4 < length_2 ? _GEN_6790 : _GEN_6630; // @[executor.scala 308:60]
  wire [7:0] _GEN_6951 = 8'h4 < length_2 ? _GEN_6791 : _GEN_6631; // @[executor.scala 308:60]
  wire [7:0] _GEN_6952 = 8'h4 < length_2 ? _GEN_6792 : _GEN_6632; // @[executor.scala 308:60]
  wire [7:0] _GEN_6953 = 8'h4 < length_2 ? _GEN_6793 : _GEN_6633; // @[executor.scala 308:60]
  wire [7:0] _GEN_6954 = 8'h4 < length_2 ? _GEN_6794 : _GEN_6634; // @[executor.scala 308:60]
  wire [7:0] _GEN_6955 = 8'h4 < length_2 ? _GEN_6795 : _GEN_6635; // @[executor.scala 308:60]
  wire [7:0] _GEN_6956 = 8'h4 < length_2 ? _GEN_6796 : _GEN_6636; // @[executor.scala 308:60]
  wire [7:0] _GEN_6957 = 8'h4 < length_2 ? _GEN_6797 : _GEN_6637; // @[executor.scala 308:60]
  wire [7:0] _GEN_6958 = 8'h4 < length_2 ? _GEN_6798 : _GEN_6638; // @[executor.scala 308:60]
  wire [7:0] _GEN_6959 = 8'h4 < length_2 ? _GEN_6799 : _GEN_6639; // @[executor.scala 308:60]
  wire [7:0] _GEN_6960 = 8'h4 < length_2 ? _GEN_6800 : _GEN_6640; // @[executor.scala 308:60]
  wire [7:0] _GEN_6961 = 8'h4 < length_2 ? _GEN_6801 : _GEN_6641; // @[executor.scala 308:60]
  wire [7:0] _GEN_6962 = 8'h4 < length_2 ? _GEN_6802 : _GEN_6642; // @[executor.scala 308:60]
  wire [7:0] _GEN_6963 = 8'h4 < length_2 ? _GEN_6803 : _GEN_6643; // @[executor.scala 308:60]
  wire [7:0] _GEN_6964 = 8'h4 < length_2 ? _GEN_6804 : _GEN_6644; // @[executor.scala 308:60]
  wire [7:0] _GEN_6965 = 8'h4 < length_2 ? _GEN_6805 : _GEN_6645; // @[executor.scala 308:60]
  wire [7:0] _GEN_6966 = 8'h4 < length_2 ? _GEN_6806 : _GEN_6646; // @[executor.scala 308:60]
  wire [7:0] _GEN_6967 = 8'h4 < length_2 ? _GEN_6807 : _GEN_6647; // @[executor.scala 308:60]
  wire [7:0] _GEN_6968 = 8'h4 < length_2 ? _GEN_6808 : _GEN_6648; // @[executor.scala 308:60]
  wire [7:0] _GEN_6969 = 8'h4 < length_2 ? _GEN_6809 : _GEN_6649; // @[executor.scala 308:60]
  wire [7:0] _GEN_6970 = 8'h4 < length_2 ? _GEN_6810 : _GEN_6650; // @[executor.scala 308:60]
  wire [7:0] _GEN_6971 = 8'h4 < length_2 ? _GEN_6811 : _GEN_6651; // @[executor.scala 308:60]
  wire [7:0] _GEN_6972 = 8'h4 < length_2 ? _GEN_6812 : _GEN_6652; // @[executor.scala 308:60]
  wire [7:0] _GEN_6973 = 8'h4 < length_2 ? _GEN_6813 : _GEN_6653; // @[executor.scala 308:60]
  wire [7:0] _GEN_6974 = 8'h4 < length_2 ? _GEN_6814 : _GEN_6654; // @[executor.scala 308:60]
  wire [7:0] _GEN_6975 = 8'h4 < length_2 ? _GEN_6815 : _GEN_6655; // @[executor.scala 308:60]
  wire [7:0] _GEN_6976 = 8'h4 < length_2 ? _GEN_6816 : _GEN_6656; // @[executor.scala 308:60]
  wire [7:0] _GEN_6977 = 8'h4 < length_2 ? _GEN_6817 : _GEN_6657; // @[executor.scala 308:60]
  wire [7:0] _GEN_6978 = 8'h4 < length_2 ? _GEN_6818 : _GEN_6658; // @[executor.scala 308:60]
  wire [7:0] _GEN_6979 = 8'h4 < length_2 ? _GEN_6819 : _GEN_6659; // @[executor.scala 308:60]
  wire [7:0] _GEN_6980 = 8'h4 < length_2 ? _GEN_6820 : _GEN_6660; // @[executor.scala 308:60]
  wire [7:0] _GEN_6981 = 8'h4 < length_2 ? _GEN_6821 : _GEN_6661; // @[executor.scala 308:60]
  wire [7:0] _GEN_6982 = 8'h4 < length_2 ? _GEN_6822 : _GEN_6662; // @[executor.scala 308:60]
  wire [7:0] _GEN_6983 = 8'h4 < length_2 ? _GEN_6823 : _GEN_6663; // @[executor.scala 308:60]
  wire [7:0] _GEN_6984 = 8'h4 < length_2 ? _GEN_6824 : _GEN_6664; // @[executor.scala 308:60]
  wire [7:0] _GEN_6985 = 8'h4 < length_2 ? _GEN_6825 : _GEN_6665; // @[executor.scala 308:60]
  wire [7:0] _GEN_6986 = 8'h4 < length_2 ? _GEN_6826 : _GEN_6666; // @[executor.scala 308:60]
  wire [7:0] _GEN_6987 = 8'h4 < length_2 ? _GEN_6827 : _GEN_6667; // @[executor.scala 308:60]
  wire [7:0] _GEN_6988 = 8'h4 < length_2 ? _GEN_6828 : _GEN_6668; // @[executor.scala 308:60]
  wire [7:0] _GEN_6989 = 8'h4 < length_2 ? _GEN_6829 : _GEN_6669; // @[executor.scala 308:60]
  wire [7:0] _GEN_6990 = 8'h4 < length_2 ? _GEN_6830 : _GEN_6670; // @[executor.scala 308:60]
  wire [7:0] _GEN_6991 = 8'h4 < length_2 ? _GEN_6831 : _GEN_6671; // @[executor.scala 308:60]
  wire [7:0] _GEN_6992 = 8'h4 < length_2 ? _GEN_6832 : _GEN_6672; // @[executor.scala 308:60]
  wire [7:0] _GEN_6993 = 8'h4 < length_2 ? _GEN_6833 : _GEN_6673; // @[executor.scala 308:60]
  wire [7:0] _GEN_6994 = 8'h4 < length_2 ? _GEN_6834 : _GEN_6674; // @[executor.scala 308:60]
  wire [7:0] _GEN_6995 = 8'h4 < length_2 ? _GEN_6835 : _GEN_6675; // @[executor.scala 308:60]
  wire [7:0] _GEN_6996 = 8'h4 < length_2 ? _GEN_6836 : _GEN_6676; // @[executor.scala 308:60]
  wire [7:0] _GEN_6997 = 8'h4 < length_2 ? _GEN_6837 : _GEN_6677; // @[executor.scala 308:60]
  wire [7:0] _GEN_6998 = 8'h4 < length_2 ? _GEN_6838 : _GEN_6678; // @[executor.scala 308:60]
  wire [7:0] _GEN_6999 = 8'h4 < length_2 ? _GEN_6839 : _GEN_6679; // @[executor.scala 308:60]
  wire [7:0] _GEN_7000 = 8'h4 < length_2 ? _GEN_6840 : _GEN_6680; // @[executor.scala 308:60]
  wire [7:0] _GEN_7001 = 8'h4 < length_2 ? _GEN_6841 : _GEN_6681; // @[executor.scala 308:60]
  wire [7:0] _GEN_7002 = 8'h4 < length_2 ? _GEN_6842 : _GEN_6682; // @[executor.scala 308:60]
  wire [7:0] _GEN_7003 = 8'h4 < length_2 ? _GEN_6843 : _GEN_6683; // @[executor.scala 308:60]
  wire [7:0] _GEN_7004 = 8'h4 < length_2 ? _GEN_6844 : _GEN_6684; // @[executor.scala 308:60]
  wire [7:0] _GEN_7005 = 8'h4 < length_2 ? _GEN_6845 : _GEN_6685; // @[executor.scala 308:60]
  wire [7:0] _GEN_7006 = 8'h4 < length_2 ? _GEN_6846 : _GEN_6686; // @[executor.scala 308:60]
  wire [7:0] _GEN_7007 = 8'h4 < length_2 ? _GEN_6847 : _GEN_6687; // @[executor.scala 308:60]
  wire [7:0] _GEN_7008 = 8'h4 < length_2 ? _GEN_6848 : _GEN_6688; // @[executor.scala 308:60]
  wire [7:0] _GEN_7009 = 8'h4 < length_2 ? _GEN_6849 : _GEN_6689; // @[executor.scala 308:60]
  wire [7:0] _GEN_7010 = 8'h4 < length_2 ? _GEN_6850 : _GEN_6690; // @[executor.scala 308:60]
  wire [7:0] _GEN_7011 = 8'h4 < length_2 ? _GEN_6851 : _GEN_6691; // @[executor.scala 308:60]
  wire [7:0] _GEN_7012 = 8'h4 < length_2 ? _GEN_6852 : _GEN_6692; // @[executor.scala 308:60]
  wire [7:0] _GEN_7013 = 8'h4 < length_2 ? _GEN_6853 : _GEN_6693; // @[executor.scala 308:60]
  wire [7:0] _GEN_7014 = 8'h4 < length_2 ? _GEN_6854 : _GEN_6694; // @[executor.scala 308:60]
  wire [7:0] _GEN_7015 = 8'h4 < length_2 ? _GEN_6855 : _GEN_6695; // @[executor.scala 308:60]
  wire [7:0] _GEN_7016 = 8'h4 < length_2 ? _GEN_6856 : _GEN_6696; // @[executor.scala 308:60]
  wire [7:0] _GEN_7017 = 8'h4 < length_2 ? _GEN_6857 : _GEN_6697; // @[executor.scala 308:60]
  wire [7:0] _GEN_7018 = 8'h4 < length_2 ? _GEN_6858 : _GEN_6698; // @[executor.scala 308:60]
  wire [7:0] _GEN_7019 = 8'h4 < length_2 ? _GEN_6859 : _GEN_6699; // @[executor.scala 308:60]
  wire [7:0] _GEN_7020 = 8'h4 < length_2 ? _GEN_6860 : _GEN_6700; // @[executor.scala 308:60]
  wire [7:0] _GEN_7021 = 8'h4 < length_2 ? _GEN_6861 : _GEN_6701; // @[executor.scala 308:60]
  wire [7:0] _GEN_7022 = 8'h4 < length_2 ? _GEN_6862 : _GEN_6702; // @[executor.scala 308:60]
  wire [7:0] _GEN_7023 = 8'h4 < length_2 ? _GEN_6863 : _GEN_6703; // @[executor.scala 308:60]
  wire [7:0] _GEN_7024 = 8'h4 < length_2 ? _GEN_6864 : _GEN_6704; // @[executor.scala 308:60]
  wire [7:0] _GEN_7025 = 8'h4 < length_2 ? _GEN_6865 : _GEN_6705; // @[executor.scala 308:60]
  wire [7:0] _GEN_7026 = 8'h4 < length_2 ? _GEN_6866 : _GEN_6706; // @[executor.scala 308:60]
  wire [7:0] _GEN_7027 = 8'h4 < length_2 ? _GEN_6867 : _GEN_6707; // @[executor.scala 308:60]
  wire [7:0] _GEN_7028 = 8'h4 < length_2 ? _GEN_6868 : _GEN_6708; // @[executor.scala 308:60]
  wire [7:0] _GEN_7029 = 8'h4 < length_2 ? _GEN_6869 : _GEN_6709; // @[executor.scala 308:60]
  wire [7:0] _GEN_7030 = 8'h4 < length_2 ? _GEN_6870 : _GEN_6710; // @[executor.scala 308:60]
  wire [7:0] _GEN_7031 = 8'h4 < length_2 ? _GEN_6871 : _GEN_6711; // @[executor.scala 308:60]
  wire [7:0] _GEN_7032 = 8'h4 < length_2 ? _GEN_6872 : _GEN_6712; // @[executor.scala 308:60]
  wire [7:0] _GEN_7033 = 8'h4 < length_2 ? _GEN_6873 : _GEN_6713; // @[executor.scala 308:60]
  wire [7:0] _GEN_7034 = 8'h4 < length_2 ? _GEN_6874 : _GEN_6714; // @[executor.scala 308:60]
  wire [7:0] _GEN_7035 = 8'h4 < length_2 ? _GEN_6875 : _GEN_6715; // @[executor.scala 308:60]
  wire [7:0] _GEN_7036 = 8'h4 < length_2 ? _GEN_6876 : _GEN_6716; // @[executor.scala 308:60]
  wire [7:0] _GEN_7037 = 8'h4 < length_2 ? _GEN_6877 : _GEN_6717; // @[executor.scala 308:60]
  wire [7:0] _GEN_7038 = 8'h4 < length_2 ? _GEN_6878 : _GEN_6718; // @[executor.scala 308:60]
  wire [7:0] _GEN_7039 = 8'h4 < length_2 ? _GEN_6879 : _GEN_6719; // @[executor.scala 308:60]
  wire [7:0] _GEN_7040 = 8'h4 < length_2 ? _GEN_6880 : _GEN_6720; // @[executor.scala 308:60]
  wire [7:0] _GEN_7041 = 8'h4 < length_2 ? _GEN_6881 : _GEN_6721; // @[executor.scala 308:60]
  wire [7:0] _GEN_7042 = 8'h4 < length_2 ? _GEN_6882 : _GEN_6722; // @[executor.scala 308:60]
  wire [7:0] _GEN_7043 = 8'h4 < length_2 ? _GEN_6883 : _GEN_6723; // @[executor.scala 308:60]
  wire [7:0] field_byte_21 = field_2[23:16]; // @[executor.scala 305:57]
  wire [7:0] total_offset_21 = offset_2 + 8'h5; // @[executor.scala 307:57]
  wire [7:0] _GEN_7044 = 8'h0 == total_offset_21 ? field_byte_21 : _GEN_6884; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7045 = 8'h1 == total_offset_21 ? field_byte_21 : _GEN_6885; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7046 = 8'h2 == total_offset_21 ? field_byte_21 : _GEN_6886; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7047 = 8'h3 == total_offset_21 ? field_byte_21 : _GEN_6887; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7048 = 8'h4 == total_offset_21 ? field_byte_21 : _GEN_6888; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7049 = 8'h5 == total_offset_21 ? field_byte_21 : _GEN_6889; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7050 = 8'h6 == total_offset_21 ? field_byte_21 : _GEN_6890; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7051 = 8'h7 == total_offset_21 ? field_byte_21 : _GEN_6891; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7052 = 8'h8 == total_offset_21 ? field_byte_21 : _GEN_6892; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7053 = 8'h9 == total_offset_21 ? field_byte_21 : _GEN_6893; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7054 = 8'ha == total_offset_21 ? field_byte_21 : _GEN_6894; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7055 = 8'hb == total_offset_21 ? field_byte_21 : _GEN_6895; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7056 = 8'hc == total_offset_21 ? field_byte_21 : _GEN_6896; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7057 = 8'hd == total_offset_21 ? field_byte_21 : _GEN_6897; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7058 = 8'he == total_offset_21 ? field_byte_21 : _GEN_6898; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7059 = 8'hf == total_offset_21 ? field_byte_21 : _GEN_6899; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7060 = 8'h10 == total_offset_21 ? field_byte_21 : _GEN_6900; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7061 = 8'h11 == total_offset_21 ? field_byte_21 : _GEN_6901; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7062 = 8'h12 == total_offset_21 ? field_byte_21 : _GEN_6902; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7063 = 8'h13 == total_offset_21 ? field_byte_21 : _GEN_6903; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7064 = 8'h14 == total_offset_21 ? field_byte_21 : _GEN_6904; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7065 = 8'h15 == total_offset_21 ? field_byte_21 : _GEN_6905; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7066 = 8'h16 == total_offset_21 ? field_byte_21 : _GEN_6906; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7067 = 8'h17 == total_offset_21 ? field_byte_21 : _GEN_6907; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7068 = 8'h18 == total_offset_21 ? field_byte_21 : _GEN_6908; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7069 = 8'h19 == total_offset_21 ? field_byte_21 : _GEN_6909; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7070 = 8'h1a == total_offset_21 ? field_byte_21 : _GEN_6910; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7071 = 8'h1b == total_offset_21 ? field_byte_21 : _GEN_6911; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7072 = 8'h1c == total_offset_21 ? field_byte_21 : _GEN_6912; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7073 = 8'h1d == total_offset_21 ? field_byte_21 : _GEN_6913; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7074 = 8'h1e == total_offset_21 ? field_byte_21 : _GEN_6914; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7075 = 8'h1f == total_offset_21 ? field_byte_21 : _GEN_6915; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7076 = 8'h20 == total_offset_21 ? field_byte_21 : _GEN_6916; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7077 = 8'h21 == total_offset_21 ? field_byte_21 : _GEN_6917; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7078 = 8'h22 == total_offset_21 ? field_byte_21 : _GEN_6918; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7079 = 8'h23 == total_offset_21 ? field_byte_21 : _GEN_6919; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7080 = 8'h24 == total_offset_21 ? field_byte_21 : _GEN_6920; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7081 = 8'h25 == total_offset_21 ? field_byte_21 : _GEN_6921; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7082 = 8'h26 == total_offset_21 ? field_byte_21 : _GEN_6922; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7083 = 8'h27 == total_offset_21 ? field_byte_21 : _GEN_6923; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7084 = 8'h28 == total_offset_21 ? field_byte_21 : _GEN_6924; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7085 = 8'h29 == total_offset_21 ? field_byte_21 : _GEN_6925; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7086 = 8'h2a == total_offset_21 ? field_byte_21 : _GEN_6926; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7087 = 8'h2b == total_offset_21 ? field_byte_21 : _GEN_6927; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7088 = 8'h2c == total_offset_21 ? field_byte_21 : _GEN_6928; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7089 = 8'h2d == total_offset_21 ? field_byte_21 : _GEN_6929; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7090 = 8'h2e == total_offset_21 ? field_byte_21 : _GEN_6930; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7091 = 8'h2f == total_offset_21 ? field_byte_21 : _GEN_6931; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7092 = 8'h30 == total_offset_21 ? field_byte_21 : _GEN_6932; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7093 = 8'h31 == total_offset_21 ? field_byte_21 : _GEN_6933; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7094 = 8'h32 == total_offset_21 ? field_byte_21 : _GEN_6934; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7095 = 8'h33 == total_offset_21 ? field_byte_21 : _GEN_6935; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7096 = 8'h34 == total_offset_21 ? field_byte_21 : _GEN_6936; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7097 = 8'h35 == total_offset_21 ? field_byte_21 : _GEN_6937; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7098 = 8'h36 == total_offset_21 ? field_byte_21 : _GEN_6938; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7099 = 8'h37 == total_offset_21 ? field_byte_21 : _GEN_6939; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7100 = 8'h38 == total_offset_21 ? field_byte_21 : _GEN_6940; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7101 = 8'h39 == total_offset_21 ? field_byte_21 : _GEN_6941; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7102 = 8'h3a == total_offset_21 ? field_byte_21 : _GEN_6942; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7103 = 8'h3b == total_offset_21 ? field_byte_21 : _GEN_6943; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7104 = 8'h3c == total_offset_21 ? field_byte_21 : _GEN_6944; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7105 = 8'h3d == total_offset_21 ? field_byte_21 : _GEN_6945; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7106 = 8'h3e == total_offset_21 ? field_byte_21 : _GEN_6946; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7107 = 8'h3f == total_offset_21 ? field_byte_21 : _GEN_6947; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7108 = 8'h40 == total_offset_21 ? field_byte_21 : _GEN_6948; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7109 = 8'h41 == total_offset_21 ? field_byte_21 : _GEN_6949; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7110 = 8'h42 == total_offset_21 ? field_byte_21 : _GEN_6950; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7111 = 8'h43 == total_offset_21 ? field_byte_21 : _GEN_6951; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7112 = 8'h44 == total_offset_21 ? field_byte_21 : _GEN_6952; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7113 = 8'h45 == total_offset_21 ? field_byte_21 : _GEN_6953; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7114 = 8'h46 == total_offset_21 ? field_byte_21 : _GEN_6954; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7115 = 8'h47 == total_offset_21 ? field_byte_21 : _GEN_6955; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7116 = 8'h48 == total_offset_21 ? field_byte_21 : _GEN_6956; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7117 = 8'h49 == total_offset_21 ? field_byte_21 : _GEN_6957; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7118 = 8'h4a == total_offset_21 ? field_byte_21 : _GEN_6958; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7119 = 8'h4b == total_offset_21 ? field_byte_21 : _GEN_6959; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7120 = 8'h4c == total_offset_21 ? field_byte_21 : _GEN_6960; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7121 = 8'h4d == total_offset_21 ? field_byte_21 : _GEN_6961; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7122 = 8'h4e == total_offset_21 ? field_byte_21 : _GEN_6962; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7123 = 8'h4f == total_offset_21 ? field_byte_21 : _GEN_6963; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7124 = 8'h50 == total_offset_21 ? field_byte_21 : _GEN_6964; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7125 = 8'h51 == total_offset_21 ? field_byte_21 : _GEN_6965; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7126 = 8'h52 == total_offset_21 ? field_byte_21 : _GEN_6966; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7127 = 8'h53 == total_offset_21 ? field_byte_21 : _GEN_6967; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7128 = 8'h54 == total_offset_21 ? field_byte_21 : _GEN_6968; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7129 = 8'h55 == total_offset_21 ? field_byte_21 : _GEN_6969; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7130 = 8'h56 == total_offset_21 ? field_byte_21 : _GEN_6970; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7131 = 8'h57 == total_offset_21 ? field_byte_21 : _GEN_6971; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7132 = 8'h58 == total_offset_21 ? field_byte_21 : _GEN_6972; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7133 = 8'h59 == total_offset_21 ? field_byte_21 : _GEN_6973; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7134 = 8'h5a == total_offset_21 ? field_byte_21 : _GEN_6974; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7135 = 8'h5b == total_offset_21 ? field_byte_21 : _GEN_6975; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7136 = 8'h5c == total_offset_21 ? field_byte_21 : _GEN_6976; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7137 = 8'h5d == total_offset_21 ? field_byte_21 : _GEN_6977; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7138 = 8'h5e == total_offset_21 ? field_byte_21 : _GEN_6978; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7139 = 8'h5f == total_offset_21 ? field_byte_21 : _GEN_6979; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7140 = 8'h60 == total_offset_21 ? field_byte_21 : _GEN_6980; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7141 = 8'h61 == total_offset_21 ? field_byte_21 : _GEN_6981; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7142 = 8'h62 == total_offset_21 ? field_byte_21 : _GEN_6982; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7143 = 8'h63 == total_offset_21 ? field_byte_21 : _GEN_6983; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7144 = 8'h64 == total_offset_21 ? field_byte_21 : _GEN_6984; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7145 = 8'h65 == total_offset_21 ? field_byte_21 : _GEN_6985; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7146 = 8'h66 == total_offset_21 ? field_byte_21 : _GEN_6986; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7147 = 8'h67 == total_offset_21 ? field_byte_21 : _GEN_6987; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7148 = 8'h68 == total_offset_21 ? field_byte_21 : _GEN_6988; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7149 = 8'h69 == total_offset_21 ? field_byte_21 : _GEN_6989; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7150 = 8'h6a == total_offset_21 ? field_byte_21 : _GEN_6990; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7151 = 8'h6b == total_offset_21 ? field_byte_21 : _GEN_6991; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7152 = 8'h6c == total_offset_21 ? field_byte_21 : _GEN_6992; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7153 = 8'h6d == total_offset_21 ? field_byte_21 : _GEN_6993; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7154 = 8'h6e == total_offset_21 ? field_byte_21 : _GEN_6994; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7155 = 8'h6f == total_offset_21 ? field_byte_21 : _GEN_6995; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7156 = 8'h70 == total_offset_21 ? field_byte_21 : _GEN_6996; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7157 = 8'h71 == total_offset_21 ? field_byte_21 : _GEN_6997; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7158 = 8'h72 == total_offset_21 ? field_byte_21 : _GEN_6998; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7159 = 8'h73 == total_offset_21 ? field_byte_21 : _GEN_6999; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7160 = 8'h74 == total_offset_21 ? field_byte_21 : _GEN_7000; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7161 = 8'h75 == total_offset_21 ? field_byte_21 : _GEN_7001; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7162 = 8'h76 == total_offset_21 ? field_byte_21 : _GEN_7002; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7163 = 8'h77 == total_offset_21 ? field_byte_21 : _GEN_7003; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7164 = 8'h78 == total_offset_21 ? field_byte_21 : _GEN_7004; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7165 = 8'h79 == total_offset_21 ? field_byte_21 : _GEN_7005; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7166 = 8'h7a == total_offset_21 ? field_byte_21 : _GEN_7006; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7167 = 8'h7b == total_offset_21 ? field_byte_21 : _GEN_7007; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7168 = 8'h7c == total_offset_21 ? field_byte_21 : _GEN_7008; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7169 = 8'h7d == total_offset_21 ? field_byte_21 : _GEN_7009; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7170 = 8'h7e == total_offset_21 ? field_byte_21 : _GEN_7010; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7171 = 8'h7f == total_offset_21 ? field_byte_21 : _GEN_7011; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7172 = 8'h80 == total_offset_21 ? field_byte_21 : _GEN_7012; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7173 = 8'h81 == total_offset_21 ? field_byte_21 : _GEN_7013; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7174 = 8'h82 == total_offset_21 ? field_byte_21 : _GEN_7014; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7175 = 8'h83 == total_offset_21 ? field_byte_21 : _GEN_7015; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7176 = 8'h84 == total_offset_21 ? field_byte_21 : _GEN_7016; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7177 = 8'h85 == total_offset_21 ? field_byte_21 : _GEN_7017; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7178 = 8'h86 == total_offset_21 ? field_byte_21 : _GEN_7018; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7179 = 8'h87 == total_offset_21 ? field_byte_21 : _GEN_7019; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7180 = 8'h88 == total_offset_21 ? field_byte_21 : _GEN_7020; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7181 = 8'h89 == total_offset_21 ? field_byte_21 : _GEN_7021; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7182 = 8'h8a == total_offset_21 ? field_byte_21 : _GEN_7022; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7183 = 8'h8b == total_offset_21 ? field_byte_21 : _GEN_7023; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7184 = 8'h8c == total_offset_21 ? field_byte_21 : _GEN_7024; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7185 = 8'h8d == total_offset_21 ? field_byte_21 : _GEN_7025; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7186 = 8'h8e == total_offset_21 ? field_byte_21 : _GEN_7026; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7187 = 8'h8f == total_offset_21 ? field_byte_21 : _GEN_7027; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7188 = 8'h90 == total_offset_21 ? field_byte_21 : _GEN_7028; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7189 = 8'h91 == total_offset_21 ? field_byte_21 : _GEN_7029; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7190 = 8'h92 == total_offset_21 ? field_byte_21 : _GEN_7030; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7191 = 8'h93 == total_offset_21 ? field_byte_21 : _GEN_7031; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7192 = 8'h94 == total_offset_21 ? field_byte_21 : _GEN_7032; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7193 = 8'h95 == total_offset_21 ? field_byte_21 : _GEN_7033; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7194 = 8'h96 == total_offset_21 ? field_byte_21 : _GEN_7034; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7195 = 8'h97 == total_offset_21 ? field_byte_21 : _GEN_7035; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7196 = 8'h98 == total_offset_21 ? field_byte_21 : _GEN_7036; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7197 = 8'h99 == total_offset_21 ? field_byte_21 : _GEN_7037; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7198 = 8'h9a == total_offset_21 ? field_byte_21 : _GEN_7038; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7199 = 8'h9b == total_offset_21 ? field_byte_21 : _GEN_7039; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7200 = 8'h9c == total_offset_21 ? field_byte_21 : _GEN_7040; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7201 = 8'h9d == total_offset_21 ? field_byte_21 : _GEN_7041; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7202 = 8'h9e == total_offset_21 ? field_byte_21 : _GEN_7042; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7203 = 8'h9f == total_offset_21 ? field_byte_21 : _GEN_7043; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7204 = 8'h5 < length_2 ? _GEN_7044 : _GEN_6884; // @[executor.scala 308:60]
  wire [7:0] _GEN_7205 = 8'h5 < length_2 ? _GEN_7045 : _GEN_6885; // @[executor.scala 308:60]
  wire [7:0] _GEN_7206 = 8'h5 < length_2 ? _GEN_7046 : _GEN_6886; // @[executor.scala 308:60]
  wire [7:0] _GEN_7207 = 8'h5 < length_2 ? _GEN_7047 : _GEN_6887; // @[executor.scala 308:60]
  wire [7:0] _GEN_7208 = 8'h5 < length_2 ? _GEN_7048 : _GEN_6888; // @[executor.scala 308:60]
  wire [7:0] _GEN_7209 = 8'h5 < length_2 ? _GEN_7049 : _GEN_6889; // @[executor.scala 308:60]
  wire [7:0] _GEN_7210 = 8'h5 < length_2 ? _GEN_7050 : _GEN_6890; // @[executor.scala 308:60]
  wire [7:0] _GEN_7211 = 8'h5 < length_2 ? _GEN_7051 : _GEN_6891; // @[executor.scala 308:60]
  wire [7:0] _GEN_7212 = 8'h5 < length_2 ? _GEN_7052 : _GEN_6892; // @[executor.scala 308:60]
  wire [7:0] _GEN_7213 = 8'h5 < length_2 ? _GEN_7053 : _GEN_6893; // @[executor.scala 308:60]
  wire [7:0] _GEN_7214 = 8'h5 < length_2 ? _GEN_7054 : _GEN_6894; // @[executor.scala 308:60]
  wire [7:0] _GEN_7215 = 8'h5 < length_2 ? _GEN_7055 : _GEN_6895; // @[executor.scala 308:60]
  wire [7:0] _GEN_7216 = 8'h5 < length_2 ? _GEN_7056 : _GEN_6896; // @[executor.scala 308:60]
  wire [7:0] _GEN_7217 = 8'h5 < length_2 ? _GEN_7057 : _GEN_6897; // @[executor.scala 308:60]
  wire [7:0] _GEN_7218 = 8'h5 < length_2 ? _GEN_7058 : _GEN_6898; // @[executor.scala 308:60]
  wire [7:0] _GEN_7219 = 8'h5 < length_2 ? _GEN_7059 : _GEN_6899; // @[executor.scala 308:60]
  wire [7:0] _GEN_7220 = 8'h5 < length_2 ? _GEN_7060 : _GEN_6900; // @[executor.scala 308:60]
  wire [7:0] _GEN_7221 = 8'h5 < length_2 ? _GEN_7061 : _GEN_6901; // @[executor.scala 308:60]
  wire [7:0] _GEN_7222 = 8'h5 < length_2 ? _GEN_7062 : _GEN_6902; // @[executor.scala 308:60]
  wire [7:0] _GEN_7223 = 8'h5 < length_2 ? _GEN_7063 : _GEN_6903; // @[executor.scala 308:60]
  wire [7:0] _GEN_7224 = 8'h5 < length_2 ? _GEN_7064 : _GEN_6904; // @[executor.scala 308:60]
  wire [7:0] _GEN_7225 = 8'h5 < length_2 ? _GEN_7065 : _GEN_6905; // @[executor.scala 308:60]
  wire [7:0] _GEN_7226 = 8'h5 < length_2 ? _GEN_7066 : _GEN_6906; // @[executor.scala 308:60]
  wire [7:0] _GEN_7227 = 8'h5 < length_2 ? _GEN_7067 : _GEN_6907; // @[executor.scala 308:60]
  wire [7:0] _GEN_7228 = 8'h5 < length_2 ? _GEN_7068 : _GEN_6908; // @[executor.scala 308:60]
  wire [7:0] _GEN_7229 = 8'h5 < length_2 ? _GEN_7069 : _GEN_6909; // @[executor.scala 308:60]
  wire [7:0] _GEN_7230 = 8'h5 < length_2 ? _GEN_7070 : _GEN_6910; // @[executor.scala 308:60]
  wire [7:0] _GEN_7231 = 8'h5 < length_2 ? _GEN_7071 : _GEN_6911; // @[executor.scala 308:60]
  wire [7:0] _GEN_7232 = 8'h5 < length_2 ? _GEN_7072 : _GEN_6912; // @[executor.scala 308:60]
  wire [7:0] _GEN_7233 = 8'h5 < length_2 ? _GEN_7073 : _GEN_6913; // @[executor.scala 308:60]
  wire [7:0] _GEN_7234 = 8'h5 < length_2 ? _GEN_7074 : _GEN_6914; // @[executor.scala 308:60]
  wire [7:0] _GEN_7235 = 8'h5 < length_2 ? _GEN_7075 : _GEN_6915; // @[executor.scala 308:60]
  wire [7:0] _GEN_7236 = 8'h5 < length_2 ? _GEN_7076 : _GEN_6916; // @[executor.scala 308:60]
  wire [7:0] _GEN_7237 = 8'h5 < length_2 ? _GEN_7077 : _GEN_6917; // @[executor.scala 308:60]
  wire [7:0] _GEN_7238 = 8'h5 < length_2 ? _GEN_7078 : _GEN_6918; // @[executor.scala 308:60]
  wire [7:0] _GEN_7239 = 8'h5 < length_2 ? _GEN_7079 : _GEN_6919; // @[executor.scala 308:60]
  wire [7:0] _GEN_7240 = 8'h5 < length_2 ? _GEN_7080 : _GEN_6920; // @[executor.scala 308:60]
  wire [7:0] _GEN_7241 = 8'h5 < length_2 ? _GEN_7081 : _GEN_6921; // @[executor.scala 308:60]
  wire [7:0] _GEN_7242 = 8'h5 < length_2 ? _GEN_7082 : _GEN_6922; // @[executor.scala 308:60]
  wire [7:0] _GEN_7243 = 8'h5 < length_2 ? _GEN_7083 : _GEN_6923; // @[executor.scala 308:60]
  wire [7:0] _GEN_7244 = 8'h5 < length_2 ? _GEN_7084 : _GEN_6924; // @[executor.scala 308:60]
  wire [7:0] _GEN_7245 = 8'h5 < length_2 ? _GEN_7085 : _GEN_6925; // @[executor.scala 308:60]
  wire [7:0] _GEN_7246 = 8'h5 < length_2 ? _GEN_7086 : _GEN_6926; // @[executor.scala 308:60]
  wire [7:0] _GEN_7247 = 8'h5 < length_2 ? _GEN_7087 : _GEN_6927; // @[executor.scala 308:60]
  wire [7:0] _GEN_7248 = 8'h5 < length_2 ? _GEN_7088 : _GEN_6928; // @[executor.scala 308:60]
  wire [7:0] _GEN_7249 = 8'h5 < length_2 ? _GEN_7089 : _GEN_6929; // @[executor.scala 308:60]
  wire [7:0] _GEN_7250 = 8'h5 < length_2 ? _GEN_7090 : _GEN_6930; // @[executor.scala 308:60]
  wire [7:0] _GEN_7251 = 8'h5 < length_2 ? _GEN_7091 : _GEN_6931; // @[executor.scala 308:60]
  wire [7:0] _GEN_7252 = 8'h5 < length_2 ? _GEN_7092 : _GEN_6932; // @[executor.scala 308:60]
  wire [7:0] _GEN_7253 = 8'h5 < length_2 ? _GEN_7093 : _GEN_6933; // @[executor.scala 308:60]
  wire [7:0] _GEN_7254 = 8'h5 < length_2 ? _GEN_7094 : _GEN_6934; // @[executor.scala 308:60]
  wire [7:0] _GEN_7255 = 8'h5 < length_2 ? _GEN_7095 : _GEN_6935; // @[executor.scala 308:60]
  wire [7:0] _GEN_7256 = 8'h5 < length_2 ? _GEN_7096 : _GEN_6936; // @[executor.scala 308:60]
  wire [7:0] _GEN_7257 = 8'h5 < length_2 ? _GEN_7097 : _GEN_6937; // @[executor.scala 308:60]
  wire [7:0] _GEN_7258 = 8'h5 < length_2 ? _GEN_7098 : _GEN_6938; // @[executor.scala 308:60]
  wire [7:0] _GEN_7259 = 8'h5 < length_2 ? _GEN_7099 : _GEN_6939; // @[executor.scala 308:60]
  wire [7:0] _GEN_7260 = 8'h5 < length_2 ? _GEN_7100 : _GEN_6940; // @[executor.scala 308:60]
  wire [7:0] _GEN_7261 = 8'h5 < length_2 ? _GEN_7101 : _GEN_6941; // @[executor.scala 308:60]
  wire [7:0] _GEN_7262 = 8'h5 < length_2 ? _GEN_7102 : _GEN_6942; // @[executor.scala 308:60]
  wire [7:0] _GEN_7263 = 8'h5 < length_2 ? _GEN_7103 : _GEN_6943; // @[executor.scala 308:60]
  wire [7:0] _GEN_7264 = 8'h5 < length_2 ? _GEN_7104 : _GEN_6944; // @[executor.scala 308:60]
  wire [7:0] _GEN_7265 = 8'h5 < length_2 ? _GEN_7105 : _GEN_6945; // @[executor.scala 308:60]
  wire [7:0] _GEN_7266 = 8'h5 < length_2 ? _GEN_7106 : _GEN_6946; // @[executor.scala 308:60]
  wire [7:0] _GEN_7267 = 8'h5 < length_2 ? _GEN_7107 : _GEN_6947; // @[executor.scala 308:60]
  wire [7:0] _GEN_7268 = 8'h5 < length_2 ? _GEN_7108 : _GEN_6948; // @[executor.scala 308:60]
  wire [7:0] _GEN_7269 = 8'h5 < length_2 ? _GEN_7109 : _GEN_6949; // @[executor.scala 308:60]
  wire [7:0] _GEN_7270 = 8'h5 < length_2 ? _GEN_7110 : _GEN_6950; // @[executor.scala 308:60]
  wire [7:0] _GEN_7271 = 8'h5 < length_2 ? _GEN_7111 : _GEN_6951; // @[executor.scala 308:60]
  wire [7:0] _GEN_7272 = 8'h5 < length_2 ? _GEN_7112 : _GEN_6952; // @[executor.scala 308:60]
  wire [7:0] _GEN_7273 = 8'h5 < length_2 ? _GEN_7113 : _GEN_6953; // @[executor.scala 308:60]
  wire [7:0] _GEN_7274 = 8'h5 < length_2 ? _GEN_7114 : _GEN_6954; // @[executor.scala 308:60]
  wire [7:0] _GEN_7275 = 8'h5 < length_2 ? _GEN_7115 : _GEN_6955; // @[executor.scala 308:60]
  wire [7:0] _GEN_7276 = 8'h5 < length_2 ? _GEN_7116 : _GEN_6956; // @[executor.scala 308:60]
  wire [7:0] _GEN_7277 = 8'h5 < length_2 ? _GEN_7117 : _GEN_6957; // @[executor.scala 308:60]
  wire [7:0] _GEN_7278 = 8'h5 < length_2 ? _GEN_7118 : _GEN_6958; // @[executor.scala 308:60]
  wire [7:0] _GEN_7279 = 8'h5 < length_2 ? _GEN_7119 : _GEN_6959; // @[executor.scala 308:60]
  wire [7:0] _GEN_7280 = 8'h5 < length_2 ? _GEN_7120 : _GEN_6960; // @[executor.scala 308:60]
  wire [7:0] _GEN_7281 = 8'h5 < length_2 ? _GEN_7121 : _GEN_6961; // @[executor.scala 308:60]
  wire [7:0] _GEN_7282 = 8'h5 < length_2 ? _GEN_7122 : _GEN_6962; // @[executor.scala 308:60]
  wire [7:0] _GEN_7283 = 8'h5 < length_2 ? _GEN_7123 : _GEN_6963; // @[executor.scala 308:60]
  wire [7:0] _GEN_7284 = 8'h5 < length_2 ? _GEN_7124 : _GEN_6964; // @[executor.scala 308:60]
  wire [7:0] _GEN_7285 = 8'h5 < length_2 ? _GEN_7125 : _GEN_6965; // @[executor.scala 308:60]
  wire [7:0] _GEN_7286 = 8'h5 < length_2 ? _GEN_7126 : _GEN_6966; // @[executor.scala 308:60]
  wire [7:0] _GEN_7287 = 8'h5 < length_2 ? _GEN_7127 : _GEN_6967; // @[executor.scala 308:60]
  wire [7:0] _GEN_7288 = 8'h5 < length_2 ? _GEN_7128 : _GEN_6968; // @[executor.scala 308:60]
  wire [7:0] _GEN_7289 = 8'h5 < length_2 ? _GEN_7129 : _GEN_6969; // @[executor.scala 308:60]
  wire [7:0] _GEN_7290 = 8'h5 < length_2 ? _GEN_7130 : _GEN_6970; // @[executor.scala 308:60]
  wire [7:0] _GEN_7291 = 8'h5 < length_2 ? _GEN_7131 : _GEN_6971; // @[executor.scala 308:60]
  wire [7:0] _GEN_7292 = 8'h5 < length_2 ? _GEN_7132 : _GEN_6972; // @[executor.scala 308:60]
  wire [7:0] _GEN_7293 = 8'h5 < length_2 ? _GEN_7133 : _GEN_6973; // @[executor.scala 308:60]
  wire [7:0] _GEN_7294 = 8'h5 < length_2 ? _GEN_7134 : _GEN_6974; // @[executor.scala 308:60]
  wire [7:0] _GEN_7295 = 8'h5 < length_2 ? _GEN_7135 : _GEN_6975; // @[executor.scala 308:60]
  wire [7:0] _GEN_7296 = 8'h5 < length_2 ? _GEN_7136 : _GEN_6976; // @[executor.scala 308:60]
  wire [7:0] _GEN_7297 = 8'h5 < length_2 ? _GEN_7137 : _GEN_6977; // @[executor.scala 308:60]
  wire [7:0] _GEN_7298 = 8'h5 < length_2 ? _GEN_7138 : _GEN_6978; // @[executor.scala 308:60]
  wire [7:0] _GEN_7299 = 8'h5 < length_2 ? _GEN_7139 : _GEN_6979; // @[executor.scala 308:60]
  wire [7:0] _GEN_7300 = 8'h5 < length_2 ? _GEN_7140 : _GEN_6980; // @[executor.scala 308:60]
  wire [7:0] _GEN_7301 = 8'h5 < length_2 ? _GEN_7141 : _GEN_6981; // @[executor.scala 308:60]
  wire [7:0] _GEN_7302 = 8'h5 < length_2 ? _GEN_7142 : _GEN_6982; // @[executor.scala 308:60]
  wire [7:0] _GEN_7303 = 8'h5 < length_2 ? _GEN_7143 : _GEN_6983; // @[executor.scala 308:60]
  wire [7:0] _GEN_7304 = 8'h5 < length_2 ? _GEN_7144 : _GEN_6984; // @[executor.scala 308:60]
  wire [7:0] _GEN_7305 = 8'h5 < length_2 ? _GEN_7145 : _GEN_6985; // @[executor.scala 308:60]
  wire [7:0] _GEN_7306 = 8'h5 < length_2 ? _GEN_7146 : _GEN_6986; // @[executor.scala 308:60]
  wire [7:0] _GEN_7307 = 8'h5 < length_2 ? _GEN_7147 : _GEN_6987; // @[executor.scala 308:60]
  wire [7:0] _GEN_7308 = 8'h5 < length_2 ? _GEN_7148 : _GEN_6988; // @[executor.scala 308:60]
  wire [7:0] _GEN_7309 = 8'h5 < length_2 ? _GEN_7149 : _GEN_6989; // @[executor.scala 308:60]
  wire [7:0] _GEN_7310 = 8'h5 < length_2 ? _GEN_7150 : _GEN_6990; // @[executor.scala 308:60]
  wire [7:0] _GEN_7311 = 8'h5 < length_2 ? _GEN_7151 : _GEN_6991; // @[executor.scala 308:60]
  wire [7:0] _GEN_7312 = 8'h5 < length_2 ? _GEN_7152 : _GEN_6992; // @[executor.scala 308:60]
  wire [7:0] _GEN_7313 = 8'h5 < length_2 ? _GEN_7153 : _GEN_6993; // @[executor.scala 308:60]
  wire [7:0] _GEN_7314 = 8'h5 < length_2 ? _GEN_7154 : _GEN_6994; // @[executor.scala 308:60]
  wire [7:0] _GEN_7315 = 8'h5 < length_2 ? _GEN_7155 : _GEN_6995; // @[executor.scala 308:60]
  wire [7:0] _GEN_7316 = 8'h5 < length_2 ? _GEN_7156 : _GEN_6996; // @[executor.scala 308:60]
  wire [7:0] _GEN_7317 = 8'h5 < length_2 ? _GEN_7157 : _GEN_6997; // @[executor.scala 308:60]
  wire [7:0] _GEN_7318 = 8'h5 < length_2 ? _GEN_7158 : _GEN_6998; // @[executor.scala 308:60]
  wire [7:0] _GEN_7319 = 8'h5 < length_2 ? _GEN_7159 : _GEN_6999; // @[executor.scala 308:60]
  wire [7:0] _GEN_7320 = 8'h5 < length_2 ? _GEN_7160 : _GEN_7000; // @[executor.scala 308:60]
  wire [7:0] _GEN_7321 = 8'h5 < length_2 ? _GEN_7161 : _GEN_7001; // @[executor.scala 308:60]
  wire [7:0] _GEN_7322 = 8'h5 < length_2 ? _GEN_7162 : _GEN_7002; // @[executor.scala 308:60]
  wire [7:0] _GEN_7323 = 8'h5 < length_2 ? _GEN_7163 : _GEN_7003; // @[executor.scala 308:60]
  wire [7:0] _GEN_7324 = 8'h5 < length_2 ? _GEN_7164 : _GEN_7004; // @[executor.scala 308:60]
  wire [7:0] _GEN_7325 = 8'h5 < length_2 ? _GEN_7165 : _GEN_7005; // @[executor.scala 308:60]
  wire [7:0] _GEN_7326 = 8'h5 < length_2 ? _GEN_7166 : _GEN_7006; // @[executor.scala 308:60]
  wire [7:0] _GEN_7327 = 8'h5 < length_2 ? _GEN_7167 : _GEN_7007; // @[executor.scala 308:60]
  wire [7:0] _GEN_7328 = 8'h5 < length_2 ? _GEN_7168 : _GEN_7008; // @[executor.scala 308:60]
  wire [7:0] _GEN_7329 = 8'h5 < length_2 ? _GEN_7169 : _GEN_7009; // @[executor.scala 308:60]
  wire [7:0] _GEN_7330 = 8'h5 < length_2 ? _GEN_7170 : _GEN_7010; // @[executor.scala 308:60]
  wire [7:0] _GEN_7331 = 8'h5 < length_2 ? _GEN_7171 : _GEN_7011; // @[executor.scala 308:60]
  wire [7:0] _GEN_7332 = 8'h5 < length_2 ? _GEN_7172 : _GEN_7012; // @[executor.scala 308:60]
  wire [7:0] _GEN_7333 = 8'h5 < length_2 ? _GEN_7173 : _GEN_7013; // @[executor.scala 308:60]
  wire [7:0] _GEN_7334 = 8'h5 < length_2 ? _GEN_7174 : _GEN_7014; // @[executor.scala 308:60]
  wire [7:0] _GEN_7335 = 8'h5 < length_2 ? _GEN_7175 : _GEN_7015; // @[executor.scala 308:60]
  wire [7:0] _GEN_7336 = 8'h5 < length_2 ? _GEN_7176 : _GEN_7016; // @[executor.scala 308:60]
  wire [7:0] _GEN_7337 = 8'h5 < length_2 ? _GEN_7177 : _GEN_7017; // @[executor.scala 308:60]
  wire [7:0] _GEN_7338 = 8'h5 < length_2 ? _GEN_7178 : _GEN_7018; // @[executor.scala 308:60]
  wire [7:0] _GEN_7339 = 8'h5 < length_2 ? _GEN_7179 : _GEN_7019; // @[executor.scala 308:60]
  wire [7:0] _GEN_7340 = 8'h5 < length_2 ? _GEN_7180 : _GEN_7020; // @[executor.scala 308:60]
  wire [7:0] _GEN_7341 = 8'h5 < length_2 ? _GEN_7181 : _GEN_7021; // @[executor.scala 308:60]
  wire [7:0] _GEN_7342 = 8'h5 < length_2 ? _GEN_7182 : _GEN_7022; // @[executor.scala 308:60]
  wire [7:0] _GEN_7343 = 8'h5 < length_2 ? _GEN_7183 : _GEN_7023; // @[executor.scala 308:60]
  wire [7:0] _GEN_7344 = 8'h5 < length_2 ? _GEN_7184 : _GEN_7024; // @[executor.scala 308:60]
  wire [7:0] _GEN_7345 = 8'h5 < length_2 ? _GEN_7185 : _GEN_7025; // @[executor.scala 308:60]
  wire [7:0] _GEN_7346 = 8'h5 < length_2 ? _GEN_7186 : _GEN_7026; // @[executor.scala 308:60]
  wire [7:0] _GEN_7347 = 8'h5 < length_2 ? _GEN_7187 : _GEN_7027; // @[executor.scala 308:60]
  wire [7:0] _GEN_7348 = 8'h5 < length_2 ? _GEN_7188 : _GEN_7028; // @[executor.scala 308:60]
  wire [7:0] _GEN_7349 = 8'h5 < length_2 ? _GEN_7189 : _GEN_7029; // @[executor.scala 308:60]
  wire [7:0] _GEN_7350 = 8'h5 < length_2 ? _GEN_7190 : _GEN_7030; // @[executor.scala 308:60]
  wire [7:0] _GEN_7351 = 8'h5 < length_2 ? _GEN_7191 : _GEN_7031; // @[executor.scala 308:60]
  wire [7:0] _GEN_7352 = 8'h5 < length_2 ? _GEN_7192 : _GEN_7032; // @[executor.scala 308:60]
  wire [7:0] _GEN_7353 = 8'h5 < length_2 ? _GEN_7193 : _GEN_7033; // @[executor.scala 308:60]
  wire [7:0] _GEN_7354 = 8'h5 < length_2 ? _GEN_7194 : _GEN_7034; // @[executor.scala 308:60]
  wire [7:0] _GEN_7355 = 8'h5 < length_2 ? _GEN_7195 : _GEN_7035; // @[executor.scala 308:60]
  wire [7:0] _GEN_7356 = 8'h5 < length_2 ? _GEN_7196 : _GEN_7036; // @[executor.scala 308:60]
  wire [7:0] _GEN_7357 = 8'h5 < length_2 ? _GEN_7197 : _GEN_7037; // @[executor.scala 308:60]
  wire [7:0] _GEN_7358 = 8'h5 < length_2 ? _GEN_7198 : _GEN_7038; // @[executor.scala 308:60]
  wire [7:0] _GEN_7359 = 8'h5 < length_2 ? _GEN_7199 : _GEN_7039; // @[executor.scala 308:60]
  wire [7:0] _GEN_7360 = 8'h5 < length_2 ? _GEN_7200 : _GEN_7040; // @[executor.scala 308:60]
  wire [7:0] _GEN_7361 = 8'h5 < length_2 ? _GEN_7201 : _GEN_7041; // @[executor.scala 308:60]
  wire [7:0] _GEN_7362 = 8'h5 < length_2 ? _GEN_7202 : _GEN_7042; // @[executor.scala 308:60]
  wire [7:0] _GEN_7363 = 8'h5 < length_2 ? _GEN_7203 : _GEN_7043; // @[executor.scala 308:60]
  wire [7:0] field_byte_22 = field_2[15:8]; // @[executor.scala 305:57]
  wire [7:0] total_offset_22 = offset_2 + 8'h6; // @[executor.scala 307:57]
  wire [7:0] _GEN_7364 = 8'h0 == total_offset_22 ? field_byte_22 : _GEN_7204; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7365 = 8'h1 == total_offset_22 ? field_byte_22 : _GEN_7205; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7366 = 8'h2 == total_offset_22 ? field_byte_22 : _GEN_7206; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7367 = 8'h3 == total_offset_22 ? field_byte_22 : _GEN_7207; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7368 = 8'h4 == total_offset_22 ? field_byte_22 : _GEN_7208; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7369 = 8'h5 == total_offset_22 ? field_byte_22 : _GEN_7209; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7370 = 8'h6 == total_offset_22 ? field_byte_22 : _GEN_7210; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7371 = 8'h7 == total_offset_22 ? field_byte_22 : _GEN_7211; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7372 = 8'h8 == total_offset_22 ? field_byte_22 : _GEN_7212; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7373 = 8'h9 == total_offset_22 ? field_byte_22 : _GEN_7213; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7374 = 8'ha == total_offset_22 ? field_byte_22 : _GEN_7214; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7375 = 8'hb == total_offset_22 ? field_byte_22 : _GEN_7215; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7376 = 8'hc == total_offset_22 ? field_byte_22 : _GEN_7216; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7377 = 8'hd == total_offset_22 ? field_byte_22 : _GEN_7217; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7378 = 8'he == total_offset_22 ? field_byte_22 : _GEN_7218; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7379 = 8'hf == total_offset_22 ? field_byte_22 : _GEN_7219; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7380 = 8'h10 == total_offset_22 ? field_byte_22 : _GEN_7220; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7381 = 8'h11 == total_offset_22 ? field_byte_22 : _GEN_7221; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7382 = 8'h12 == total_offset_22 ? field_byte_22 : _GEN_7222; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7383 = 8'h13 == total_offset_22 ? field_byte_22 : _GEN_7223; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7384 = 8'h14 == total_offset_22 ? field_byte_22 : _GEN_7224; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7385 = 8'h15 == total_offset_22 ? field_byte_22 : _GEN_7225; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7386 = 8'h16 == total_offset_22 ? field_byte_22 : _GEN_7226; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7387 = 8'h17 == total_offset_22 ? field_byte_22 : _GEN_7227; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7388 = 8'h18 == total_offset_22 ? field_byte_22 : _GEN_7228; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7389 = 8'h19 == total_offset_22 ? field_byte_22 : _GEN_7229; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7390 = 8'h1a == total_offset_22 ? field_byte_22 : _GEN_7230; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7391 = 8'h1b == total_offset_22 ? field_byte_22 : _GEN_7231; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7392 = 8'h1c == total_offset_22 ? field_byte_22 : _GEN_7232; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7393 = 8'h1d == total_offset_22 ? field_byte_22 : _GEN_7233; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7394 = 8'h1e == total_offset_22 ? field_byte_22 : _GEN_7234; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7395 = 8'h1f == total_offset_22 ? field_byte_22 : _GEN_7235; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7396 = 8'h20 == total_offset_22 ? field_byte_22 : _GEN_7236; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7397 = 8'h21 == total_offset_22 ? field_byte_22 : _GEN_7237; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7398 = 8'h22 == total_offset_22 ? field_byte_22 : _GEN_7238; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7399 = 8'h23 == total_offset_22 ? field_byte_22 : _GEN_7239; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7400 = 8'h24 == total_offset_22 ? field_byte_22 : _GEN_7240; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7401 = 8'h25 == total_offset_22 ? field_byte_22 : _GEN_7241; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7402 = 8'h26 == total_offset_22 ? field_byte_22 : _GEN_7242; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7403 = 8'h27 == total_offset_22 ? field_byte_22 : _GEN_7243; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7404 = 8'h28 == total_offset_22 ? field_byte_22 : _GEN_7244; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7405 = 8'h29 == total_offset_22 ? field_byte_22 : _GEN_7245; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7406 = 8'h2a == total_offset_22 ? field_byte_22 : _GEN_7246; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7407 = 8'h2b == total_offset_22 ? field_byte_22 : _GEN_7247; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7408 = 8'h2c == total_offset_22 ? field_byte_22 : _GEN_7248; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7409 = 8'h2d == total_offset_22 ? field_byte_22 : _GEN_7249; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7410 = 8'h2e == total_offset_22 ? field_byte_22 : _GEN_7250; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7411 = 8'h2f == total_offset_22 ? field_byte_22 : _GEN_7251; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7412 = 8'h30 == total_offset_22 ? field_byte_22 : _GEN_7252; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7413 = 8'h31 == total_offset_22 ? field_byte_22 : _GEN_7253; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7414 = 8'h32 == total_offset_22 ? field_byte_22 : _GEN_7254; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7415 = 8'h33 == total_offset_22 ? field_byte_22 : _GEN_7255; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7416 = 8'h34 == total_offset_22 ? field_byte_22 : _GEN_7256; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7417 = 8'h35 == total_offset_22 ? field_byte_22 : _GEN_7257; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7418 = 8'h36 == total_offset_22 ? field_byte_22 : _GEN_7258; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7419 = 8'h37 == total_offset_22 ? field_byte_22 : _GEN_7259; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7420 = 8'h38 == total_offset_22 ? field_byte_22 : _GEN_7260; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7421 = 8'h39 == total_offset_22 ? field_byte_22 : _GEN_7261; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7422 = 8'h3a == total_offset_22 ? field_byte_22 : _GEN_7262; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7423 = 8'h3b == total_offset_22 ? field_byte_22 : _GEN_7263; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7424 = 8'h3c == total_offset_22 ? field_byte_22 : _GEN_7264; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7425 = 8'h3d == total_offset_22 ? field_byte_22 : _GEN_7265; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7426 = 8'h3e == total_offset_22 ? field_byte_22 : _GEN_7266; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7427 = 8'h3f == total_offset_22 ? field_byte_22 : _GEN_7267; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7428 = 8'h40 == total_offset_22 ? field_byte_22 : _GEN_7268; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7429 = 8'h41 == total_offset_22 ? field_byte_22 : _GEN_7269; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7430 = 8'h42 == total_offset_22 ? field_byte_22 : _GEN_7270; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7431 = 8'h43 == total_offset_22 ? field_byte_22 : _GEN_7271; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7432 = 8'h44 == total_offset_22 ? field_byte_22 : _GEN_7272; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7433 = 8'h45 == total_offset_22 ? field_byte_22 : _GEN_7273; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7434 = 8'h46 == total_offset_22 ? field_byte_22 : _GEN_7274; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7435 = 8'h47 == total_offset_22 ? field_byte_22 : _GEN_7275; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7436 = 8'h48 == total_offset_22 ? field_byte_22 : _GEN_7276; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7437 = 8'h49 == total_offset_22 ? field_byte_22 : _GEN_7277; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7438 = 8'h4a == total_offset_22 ? field_byte_22 : _GEN_7278; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7439 = 8'h4b == total_offset_22 ? field_byte_22 : _GEN_7279; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7440 = 8'h4c == total_offset_22 ? field_byte_22 : _GEN_7280; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7441 = 8'h4d == total_offset_22 ? field_byte_22 : _GEN_7281; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7442 = 8'h4e == total_offset_22 ? field_byte_22 : _GEN_7282; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7443 = 8'h4f == total_offset_22 ? field_byte_22 : _GEN_7283; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7444 = 8'h50 == total_offset_22 ? field_byte_22 : _GEN_7284; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7445 = 8'h51 == total_offset_22 ? field_byte_22 : _GEN_7285; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7446 = 8'h52 == total_offset_22 ? field_byte_22 : _GEN_7286; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7447 = 8'h53 == total_offset_22 ? field_byte_22 : _GEN_7287; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7448 = 8'h54 == total_offset_22 ? field_byte_22 : _GEN_7288; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7449 = 8'h55 == total_offset_22 ? field_byte_22 : _GEN_7289; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7450 = 8'h56 == total_offset_22 ? field_byte_22 : _GEN_7290; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7451 = 8'h57 == total_offset_22 ? field_byte_22 : _GEN_7291; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7452 = 8'h58 == total_offset_22 ? field_byte_22 : _GEN_7292; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7453 = 8'h59 == total_offset_22 ? field_byte_22 : _GEN_7293; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7454 = 8'h5a == total_offset_22 ? field_byte_22 : _GEN_7294; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7455 = 8'h5b == total_offset_22 ? field_byte_22 : _GEN_7295; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7456 = 8'h5c == total_offset_22 ? field_byte_22 : _GEN_7296; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7457 = 8'h5d == total_offset_22 ? field_byte_22 : _GEN_7297; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7458 = 8'h5e == total_offset_22 ? field_byte_22 : _GEN_7298; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7459 = 8'h5f == total_offset_22 ? field_byte_22 : _GEN_7299; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7460 = 8'h60 == total_offset_22 ? field_byte_22 : _GEN_7300; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7461 = 8'h61 == total_offset_22 ? field_byte_22 : _GEN_7301; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7462 = 8'h62 == total_offset_22 ? field_byte_22 : _GEN_7302; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7463 = 8'h63 == total_offset_22 ? field_byte_22 : _GEN_7303; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7464 = 8'h64 == total_offset_22 ? field_byte_22 : _GEN_7304; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7465 = 8'h65 == total_offset_22 ? field_byte_22 : _GEN_7305; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7466 = 8'h66 == total_offset_22 ? field_byte_22 : _GEN_7306; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7467 = 8'h67 == total_offset_22 ? field_byte_22 : _GEN_7307; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7468 = 8'h68 == total_offset_22 ? field_byte_22 : _GEN_7308; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7469 = 8'h69 == total_offset_22 ? field_byte_22 : _GEN_7309; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7470 = 8'h6a == total_offset_22 ? field_byte_22 : _GEN_7310; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7471 = 8'h6b == total_offset_22 ? field_byte_22 : _GEN_7311; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7472 = 8'h6c == total_offset_22 ? field_byte_22 : _GEN_7312; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7473 = 8'h6d == total_offset_22 ? field_byte_22 : _GEN_7313; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7474 = 8'h6e == total_offset_22 ? field_byte_22 : _GEN_7314; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7475 = 8'h6f == total_offset_22 ? field_byte_22 : _GEN_7315; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7476 = 8'h70 == total_offset_22 ? field_byte_22 : _GEN_7316; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7477 = 8'h71 == total_offset_22 ? field_byte_22 : _GEN_7317; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7478 = 8'h72 == total_offset_22 ? field_byte_22 : _GEN_7318; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7479 = 8'h73 == total_offset_22 ? field_byte_22 : _GEN_7319; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7480 = 8'h74 == total_offset_22 ? field_byte_22 : _GEN_7320; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7481 = 8'h75 == total_offset_22 ? field_byte_22 : _GEN_7321; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7482 = 8'h76 == total_offset_22 ? field_byte_22 : _GEN_7322; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7483 = 8'h77 == total_offset_22 ? field_byte_22 : _GEN_7323; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7484 = 8'h78 == total_offset_22 ? field_byte_22 : _GEN_7324; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7485 = 8'h79 == total_offset_22 ? field_byte_22 : _GEN_7325; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7486 = 8'h7a == total_offset_22 ? field_byte_22 : _GEN_7326; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7487 = 8'h7b == total_offset_22 ? field_byte_22 : _GEN_7327; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7488 = 8'h7c == total_offset_22 ? field_byte_22 : _GEN_7328; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7489 = 8'h7d == total_offset_22 ? field_byte_22 : _GEN_7329; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7490 = 8'h7e == total_offset_22 ? field_byte_22 : _GEN_7330; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7491 = 8'h7f == total_offset_22 ? field_byte_22 : _GEN_7331; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7492 = 8'h80 == total_offset_22 ? field_byte_22 : _GEN_7332; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7493 = 8'h81 == total_offset_22 ? field_byte_22 : _GEN_7333; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7494 = 8'h82 == total_offset_22 ? field_byte_22 : _GEN_7334; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7495 = 8'h83 == total_offset_22 ? field_byte_22 : _GEN_7335; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7496 = 8'h84 == total_offset_22 ? field_byte_22 : _GEN_7336; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7497 = 8'h85 == total_offset_22 ? field_byte_22 : _GEN_7337; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7498 = 8'h86 == total_offset_22 ? field_byte_22 : _GEN_7338; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7499 = 8'h87 == total_offset_22 ? field_byte_22 : _GEN_7339; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7500 = 8'h88 == total_offset_22 ? field_byte_22 : _GEN_7340; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7501 = 8'h89 == total_offset_22 ? field_byte_22 : _GEN_7341; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7502 = 8'h8a == total_offset_22 ? field_byte_22 : _GEN_7342; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7503 = 8'h8b == total_offset_22 ? field_byte_22 : _GEN_7343; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7504 = 8'h8c == total_offset_22 ? field_byte_22 : _GEN_7344; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7505 = 8'h8d == total_offset_22 ? field_byte_22 : _GEN_7345; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7506 = 8'h8e == total_offset_22 ? field_byte_22 : _GEN_7346; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7507 = 8'h8f == total_offset_22 ? field_byte_22 : _GEN_7347; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7508 = 8'h90 == total_offset_22 ? field_byte_22 : _GEN_7348; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7509 = 8'h91 == total_offset_22 ? field_byte_22 : _GEN_7349; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7510 = 8'h92 == total_offset_22 ? field_byte_22 : _GEN_7350; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7511 = 8'h93 == total_offset_22 ? field_byte_22 : _GEN_7351; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7512 = 8'h94 == total_offset_22 ? field_byte_22 : _GEN_7352; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7513 = 8'h95 == total_offset_22 ? field_byte_22 : _GEN_7353; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7514 = 8'h96 == total_offset_22 ? field_byte_22 : _GEN_7354; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7515 = 8'h97 == total_offset_22 ? field_byte_22 : _GEN_7355; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7516 = 8'h98 == total_offset_22 ? field_byte_22 : _GEN_7356; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7517 = 8'h99 == total_offset_22 ? field_byte_22 : _GEN_7357; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7518 = 8'h9a == total_offset_22 ? field_byte_22 : _GEN_7358; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7519 = 8'h9b == total_offset_22 ? field_byte_22 : _GEN_7359; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7520 = 8'h9c == total_offset_22 ? field_byte_22 : _GEN_7360; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7521 = 8'h9d == total_offset_22 ? field_byte_22 : _GEN_7361; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7522 = 8'h9e == total_offset_22 ? field_byte_22 : _GEN_7362; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7523 = 8'h9f == total_offset_22 ? field_byte_22 : _GEN_7363; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7524 = 8'h6 < length_2 ? _GEN_7364 : _GEN_7204; // @[executor.scala 308:60]
  wire [7:0] _GEN_7525 = 8'h6 < length_2 ? _GEN_7365 : _GEN_7205; // @[executor.scala 308:60]
  wire [7:0] _GEN_7526 = 8'h6 < length_2 ? _GEN_7366 : _GEN_7206; // @[executor.scala 308:60]
  wire [7:0] _GEN_7527 = 8'h6 < length_2 ? _GEN_7367 : _GEN_7207; // @[executor.scala 308:60]
  wire [7:0] _GEN_7528 = 8'h6 < length_2 ? _GEN_7368 : _GEN_7208; // @[executor.scala 308:60]
  wire [7:0] _GEN_7529 = 8'h6 < length_2 ? _GEN_7369 : _GEN_7209; // @[executor.scala 308:60]
  wire [7:0] _GEN_7530 = 8'h6 < length_2 ? _GEN_7370 : _GEN_7210; // @[executor.scala 308:60]
  wire [7:0] _GEN_7531 = 8'h6 < length_2 ? _GEN_7371 : _GEN_7211; // @[executor.scala 308:60]
  wire [7:0] _GEN_7532 = 8'h6 < length_2 ? _GEN_7372 : _GEN_7212; // @[executor.scala 308:60]
  wire [7:0] _GEN_7533 = 8'h6 < length_2 ? _GEN_7373 : _GEN_7213; // @[executor.scala 308:60]
  wire [7:0] _GEN_7534 = 8'h6 < length_2 ? _GEN_7374 : _GEN_7214; // @[executor.scala 308:60]
  wire [7:0] _GEN_7535 = 8'h6 < length_2 ? _GEN_7375 : _GEN_7215; // @[executor.scala 308:60]
  wire [7:0] _GEN_7536 = 8'h6 < length_2 ? _GEN_7376 : _GEN_7216; // @[executor.scala 308:60]
  wire [7:0] _GEN_7537 = 8'h6 < length_2 ? _GEN_7377 : _GEN_7217; // @[executor.scala 308:60]
  wire [7:0] _GEN_7538 = 8'h6 < length_2 ? _GEN_7378 : _GEN_7218; // @[executor.scala 308:60]
  wire [7:0] _GEN_7539 = 8'h6 < length_2 ? _GEN_7379 : _GEN_7219; // @[executor.scala 308:60]
  wire [7:0] _GEN_7540 = 8'h6 < length_2 ? _GEN_7380 : _GEN_7220; // @[executor.scala 308:60]
  wire [7:0] _GEN_7541 = 8'h6 < length_2 ? _GEN_7381 : _GEN_7221; // @[executor.scala 308:60]
  wire [7:0] _GEN_7542 = 8'h6 < length_2 ? _GEN_7382 : _GEN_7222; // @[executor.scala 308:60]
  wire [7:0] _GEN_7543 = 8'h6 < length_2 ? _GEN_7383 : _GEN_7223; // @[executor.scala 308:60]
  wire [7:0] _GEN_7544 = 8'h6 < length_2 ? _GEN_7384 : _GEN_7224; // @[executor.scala 308:60]
  wire [7:0] _GEN_7545 = 8'h6 < length_2 ? _GEN_7385 : _GEN_7225; // @[executor.scala 308:60]
  wire [7:0] _GEN_7546 = 8'h6 < length_2 ? _GEN_7386 : _GEN_7226; // @[executor.scala 308:60]
  wire [7:0] _GEN_7547 = 8'h6 < length_2 ? _GEN_7387 : _GEN_7227; // @[executor.scala 308:60]
  wire [7:0] _GEN_7548 = 8'h6 < length_2 ? _GEN_7388 : _GEN_7228; // @[executor.scala 308:60]
  wire [7:0] _GEN_7549 = 8'h6 < length_2 ? _GEN_7389 : _GEN_7229; // @[executor.scala 308:60]
  wire [7:0] _GEN_7550 = 8'h6 < length_2 ? _GEN_7390 : _GEN_7230; // @[executor.scala 308:60]
  wire [7:0] _GEN_7551 = 8'h6 < length_2 ? _GEN_7391 : _GEN_7231; // @[executor.scala 308:60]
  wire [7:0] _GEN_7552 = 8'h6 < length_2 ? _GEN_7392 : _GEN_7232; // @[executor.scala 308:60]
  wire [7:0] _GEN_7553 = 8'h6 < length_2 ? _GEN_7393 : _GEN_7233; // @[executor.scala 308:60]
  wire [7:0] _GEN_7554 = 8'h6 < length_2 ? _GEN_7394 : _GEN_7234; // @[executor.scala 308:60]
  wire [7:0] _GEN_7555 = 8'h6 < length_2 ? _GEN_7395 : _GEN_7235; // @[executor.scala 308:60]
  wire [7:0] _GEN_7556 = 8'h6 < length_2 ? _GEN_7396 : _GEN_7236; // @[executor.scala 308:60]
  wire [7:0] _GEN_7557 = 8'h6 < length_2 ? _GEN_7397 : _GEN_7237; // @[executor.scala 308:60]
  wire [7:0] _GEN_7558 = 8'h6 < length_2 ? _GEN_7398 : _GEN_7238; // @[executor.scala 308:60]
  wire [7:0] _GEN_7559 = 8'h6 < length_2 ? _GEN_7399 : _GEN_7239; // @[executor.scala 308:60]
  wire [7:0] _GEN_7560 = 8'h6 < length_2 ? _GEN_7400 : _GEN_7240; // @[executor.scala 308:60]
  wire [7:0] _GEN_7561 = 8'h6 < length_2 ? _GEN_7401 : _GEN_7241; // @[executor.scala 308:60]
  wire [7:0] _GEN_7562 = 8'h6 < length_2 ? _GEN_7402 : _GEN_7242; // @[executor.scala 308:60]
  wire [7:0] _GEN_7563 = 8'h6 < length_2 ? _GEN_7403 : _GEN_7243; // @[executor.scala 308:60]
  wire [7:0] _GEN_7564 = 8'h6 < length_2 ? _GEN_7404 : _GEN_7244; // @[executor.scala 308:60]
  wire [7:0] _GEN_7565 = 8'h6 < length_2 ? _GEN_7405 : _GEN_7245; // @[executor.scala 308:60]
  wire [7:0] _GEN_7566 = 8'h6 < length_2 ? _GEN_7406 : _GEN_7246; // @[executor.scala 308:60]
  wire [7:0] _GEN_7567 = 8'h6 < length_2 ? _GEN_7407 : _GEN_7247; // @[executor.scala 308:60]
  wire [7:0] _GEN_7568 = 8'h6 < length_2 ? _GEN_7408 : _GEN_7248; // @[executor.scala 308:60]
  wire [7:0] _GEN_7569 = 8'h6 < length_2 ? _GEN_7409 : _GEN_7249; // @[executor.scala 308:60]
  wire [7:0] _GEN_7570 = 8'h6 < length_2 ? _GEN_7410 : _GEN_7250; // @[executor.scala 308:60]
  wire [7:0] _GEN_7571 = 8'h6 < length_2 ? _GEN_7411 : _GEN_7251; // @[executor.scala 308:60]
  wire [7:0] _GEN_7572 = 8'h6 < length_2 ? _GEN_7412 : _GEN_7252; // @[executor.scala 308:60]
  wire [7:0] _GEN_7573 = 8'h6 < length_2 ? _GEN_7413 : _GEN_7253; // @[executor.scala 308:60]
  wire [7:0] _GEN_7574 = 8'h6 < length_2 ? _GEN_7414 : _GEN_7254; // @[executor.scala 308:60]
  wire [7:0] _GEN_7575 = 8'h6 < length_2 ? _GEN_7415 : _GEN_7255; // @[executor.scala 308:60]
  wire [7:0] _GEN_7576 = 8'h6 < length_2 ? _GEN_7416 : _GEN_7256; // @[executor.scala 308:60]
  wire [7:0] _GEN_7577 = 8'h6 < length_2 ? _GEN_7417 : _GEN_7257; // @[executor.scala 308:60]
  wire [7:0] _GEN_7578 = 8'h6 < length_2 ? _GEN_7418 : _GEN_7258; // @[executor.scala 308:60]
  wire [7:0] _GEN_7579 = 8'h6 < length_2 ? _GEN_7419 : _GEN_7259; // @[executor.scala 308:60]
  wire [7:0] _GEN_7580 = 8'h6 < length_2 ? _GEN_7420 : _GEN_7260; // @[executor.scala 308:60]
  wire [7:0] _GEN_7581 = 8'h6 < length_2 ? _GEN_7421 : _GEN_7261; // @[executor.scala 308:60]
  wire [7:0] _GEN_7582 = 8'h6 < length_2 ? _GEN_7422 : _GEN_7262; // @[executor.scala 308:60]
  wire [7:0] _GEN_7583 = 8'h6 < length_2 ? _GEN_7423 : _GEN_7263; // @[executor.scala 308:60]
  wire [7:0] _GEN_7584 = 8'h6 < length_2 ? _GEN_7424 : _GEN_7264; // @[executor.scala 308:60]
  wire [7:0] _GEN_7585 = 8'h6 < length_2 ? _GEN_7425 : _GEN_7265; // @[executor.scala 308:60]
  wire [7:0] _GEN_7586 = 8'h6 < length_2 ? _GEN_7426 : _GEN_7266; // @[executor.scala 308:60]
  wire [7:0] _GEN_7587 = 8'h6 < length_2 ? _GEN_7427 : _GEN_7267; // @[executor.scala 308:60]
  wire [7:0] _GEN_7588 = 8'h6 < length_2 ? _GEN_7428 : _GEN_7268; // @[executor.scala 308:60]
  wire [7:0] _GEN_7589 = 8'h6 < length_2 ? _GEN_7429 : _GEN_7269; // @[executor.scala 308:60]
  wire [7:0] _GEN_7590 = 8'h6 < length_2 ? _GEN_7430 : _GEN_7270; // @[executor.scala 308:60]
  wire [7:0] _GEN_7591 = 8'h6 < length_2 ? _GEN_7431 : _GEN_7271; // @[executor.scala 308:60]
  wire [7:0] _GEN_7592 = 8'h6 < length_2 ? _GEN_7432 : _GEN_7272; // @[executor.scala 308:60]
  wire [7:0] _GEN_7593 = 8'h6 < length_2 ? _GEN_7433 : _GEN_7273; // @[executor.scala 308:60]
  wire [7:0] _GEN_7594 = 8'h6 < length_2 ? _GEN_7434 : _GEN_7274; // @[executor.scala 308:60]
  wire [7:0] _GEN_7595 = 8'h6 < length_2 ? _GEN_7435 : _GEN_7275; // @[executor.scala 308:60]
  wire [7:0] _GEN_7596 = 8'h6 < length_2 ? _GEN_7436 : _GEN_7276; // @[executor.scala 308:60]
  wire [7:0] _GEN_7597 = 8'h6 < length_2 ? _GEN_7437 : _GEN_7277; // @[executor.scala 308:60]
  wire [7:0] _GEN_7598 = 8'h6 < length_2 ? _GEN_7438 : _GEN_7278; // @[executor.scala 308:60]
  wire [7:0] _GEN_7599 = 8'h6 < length_2 ? _GEN_7439 : _GEN_7279; // @[executor.scala 308:60]
  wire [7:0] _GEN_7600 = 8'h6 < length_2 ? _GEN_7440 : _GEN_7280; // @[executor.scala 308:60]
  wire [7:0] _GEN_7601 = 8'h6 < length_2 ? _GEN_7441 : _GEN_7281; // @[executor.scala 308:60]
  wire [7:0] _GEN_7602 = 8'h6 < length_2 ? _GEN_7442 : _GEN_7282; // @[executor.scala 308:60]
  wire [7:0] _GEN_7603 = 8'h6 < length_2 ? _GEN_7443 : _GEN_7283; // @[executor.scala 308:60]
  wire [7:0] _GEN_7604 = 8'h6 < length_2 ? _GEN_7444 : _GEN_7284; // @[executor.scala 308:60]
  wire [7:0] _GEN_7605 = 8'h6 < length_2 ? _GEN_7445 : _GEN_7285; // @[executor.scala 308:60]
  wire [7:0] _GEN_7606 = 8'h6 < length_2 ? _GEN_7446 : _GEN_7286; // @[executor.scala 308:60]
  wire [7:0] _GEN_7607 = 8'h6 < length_2 ? _GEN_7447 : _GEN_7287; // @[executor.scala 308:60]
  wire [7:0] _GEN_7608 = 8'h6 < length_2 ? _GEN_7448 : _GEN_7288; // @[executor.scala 308:60]
  wire [7:0] _GEN_7609 = 8'h6 < length_2 ? _GEN_7449 : _GEN_7289; // @[executor.scala 308:60]
  wire [7:0] _GEN_7610 = 8'h6 < length_2 ? _GEN_7450 : _GEN_7290; // @[executor.scala 308:60]
  wire [7:0] _GEN_7611 = 8'h6 < length_2 ? _GEN_7451 : _GEN_7291; // @[executor.scala 308:60]
  wire [7:0] _GEN_7612 = 8'h6 < length_2 ? _GEN_7452 : _GEN_7292; // @[executor.scala 308:60]
  wire [7:0] _GEN_7613 = 8'h6 < length_2 ? _GEN_7453 : _GEN_7293; // @[executor.scala 308:60]
  wire [7:0] _GEN_7614 = 8'h6 < length_2 ? _GEN_7454 : _GEN_7294; // @[executor.scala 308:60]
  wire [7:0] _GEN_7615 = 8'h6 < length_2 ? _GEN_7455 : _GEN_7295; // @[executor.scala 308:60]
  wire [7:0] _GEN_7616 = 8'h6 < length_2 ? _GEN_7456 : _GEN_7296; // @[executor.scala 308:60]
  wire [7:0] _GEN_7617 = 8'h6 < length_2 ? _GEN_7457 : _GEN_7297; // @[executor.scala 308:60]
  wire [7:0] _GEN_7618 = 8'h6 < length_2 ? _GEN_7458 : _GEN_7298; // @[executor.scala 308:60]
  wire [7:0] _GEN_7619 = 8'h6 < length_2 ? _GEN_7459 : _GEN_7299; // @[executor.scala 308:60]
  wire [7:0] _GEN_7620 = 8'h6 < length_2 ? _GEN_7460 : _GEN_7300; // @[executor.scala 308:60]
  wire [7:0] _GEN_7621 = 8'h6 < length_2 ? _GEN_7461 : _GEN_7301; // @[executor.scala 308:60]
  wire [7:0] _GEN_7622 = 8'h6 < length_2 ? _GEN_7462 : _GEN_7302; // @[executor.scala 308:60]
  wire [7:0] _GEN_7623 = 8'h6 < length_2 ? _GEN_7463 : _GEN_7303; // @[executor.scala 308:60]
  wire [7:0] _GEN_7624 = 8'h6 < length_2 ? _GEN_7464 : _GEN_7304; // @[executor.scala 308:60]
  wire [7:0] _GEN_7625 = 8'h6 < length_2 ? _GEN_7465 : _GEN_7305; // @[executor.scala 308:60]
  wire [7:0] _GEN_7626 = 8'h6 < length_2 ? _GEN_7466 : _GEN_7306; // @[executor.scala 308:60]
  wire [7:0] _GEN_7627 = 8'h6 < length_2 ? _GEN_7467 : _GEN_7307; // @[executor.scala 308:60]
  wire [7:0] _GEN_7628 = 8'h6 < length_2 ? _GEN_7468 : _GEN_7308; // @[executor.scala 308:60]
  wire [7:0] _GEN_7629 = 8'h6 < length_2 ? _GEN_7469 : _GEN_7309; // @[executor.scala 308:60]
  wire [7:0] _GEN_7630 = 8'h6 < length_2 ? _GEN_7470 : _GEN_7310; // @[executor.scala 308:60]
  wire [7:0] _GEN_7631 = 8'h6 < length_2 ? _GEN_7471 : _GEN_7311; // @[executor.scala 308:60]
  wire [7:0] _GEN_7632 = 8'h6 < length_2 ? _GEN_7472 : _GEN_7312; // @[executor.scala 308:60]
  wire [7:0] _GEN_7633 = 8'h6 < length_2 ? _GEN_7473 : _GEN_7313; // @[executor.scala 308:60]
  wire [7:0] _GEN_7634 = 8'h6 < length_2 ? _GEN_7474 : _GEN_7314; // @[executor.scala 308:60]
  wire [7:0] _GEN_7635 = 8'h6 < length_2 ? _GEN_7475 : _GEN_7315; // @[executor.scala 308:60]
  wire [7:0] _GEN_7636 = 8'h6 < length_2 ? _GEN_7476 : _GEN_7316; // @[executor.scala 308:60]
  wire [7:0] _GEN_7637 = 8'h6 < length_2 ? _GEN_7477 : _GEN_7317; // @[executor.scala 308:60]
  wire [7:0] _GEN_7638 = 8'h6 < length_2 ? _GEN_7478 : _GEN_7318; // @[executor.scala 308:60]
  wire [7:0] _GEN_7639 = 8'h6 < length_2 ? _GEN_7479 : _GEN_7319; // @[executor.scala 308:60]
  wire [7:0] _GEN_7640 = 8'h6 < length_2 ? _GEN_7480 : _GEN_7320; // @[executor.scala 308:60]
  wire [7:0] _GEN_7641 = 8'h6 < length_2 ? _GEN_7481 : _GEN_7321; // @[executor.scala 308:60]
  wire [7:0] _GEN_7642 = 8'h6 < length_2 ? _GEN_7482 : _GEN_7322; // @[executor.scala 308:60]
  wire [7:0] _GEN_7643 = 8'h6 < length_2 ? _GEN_7483 : _GEN_7323; // @[executor.scala 308:60]
  wire [7:0] _GEN_7644 = 8'h6 < length_2 ? _GEN_7484 : _GEN_7324; // @[executor.scala 308:60]
  wire [7:0] _GEN_7645 = 8'h6 < length_2 ? _GEN_7485 : _GEN_7325; // @[executor.scala 308:60]
  wire [7:0] _GEN_7646 = 8'h6 < length_2 ? _GEN_7486 : _GEN_7326; // @[executor.scala 308:60]
  wire [7:0] _GEN_7647 = 8'h6 < length_2 ? _GEN_7487 : _GEN_7327; // @[executor.scala 308:60]
  wire [7:0] _GEN_7648 = 8'h6 < length_2 ? _GEN_7488 : _GEN_7328; // @[executor.scala 308:60]
  wire [7:0] _GEN_7649 = 8'h6 < length_2 ? _GEN_7489 : _GEN_7329; // @[executor.scala 308:60]
  wire [7:0] _GEN_7650 = 8'h6 < length_2 ? _GEN_7490 : _GEN_7330; // @[executor.scala 308:60]
  wire [7:0] _GEN_7651 = 8'h6 < length_2 ? _GEN_7491 : _GEN_7331; // @[executor.scala 308:60]
  wire [7:0] _GEN_7652 = 8'h6 < length_2 ? _GEN_7492 : _GEN_7332; // @[executor.scala 308:60]
  wire [7:0] _GEN_7653 = 8'h6 < length_2 ? _GEN_7493 : _GEN_7333; // @[executor.scala 308:60]
  wire [7:0] _GEN_7654 = 8'h6 < length_2 ? _GEN_7494 : _GEN_7334; // @[executor.scala 308:60]
  wire [7:0] _GEN_7655 = 8'h6 < length_2 ? _GEN_7495 : _GEN_7335; // @[executor.scala 308:60]
  wire [7:0] _GEN_7656 = 8'h6 < length_2 ? _GEN_7496 : _GEN_7336; // @[executor.scala 308:60]
  wire [7:0] _GEN_7657 = 8'h6 < length_2 ? _GEN_7497 : _GEN_7337; // @[executor.scala 308:60]
  wire [7:0] _GEN_7658 = 8'h6 < length_2 ? _GEN_7498 : _GEN_7338; // @[executor.scala 308:60]
  wire [7:0] _GEN_7659 = 8'h6 < length_2 ? _GEN_7499 : _GEN_7339; // @[executor.scala 308:60]
  wire [7:0] _GEN_7660 = 8'h6 < length_2 ? _GEN_7500 : _GEN_7340; // @[executor.scala 308:60]
  wire [7:0] _GEN_7661 = 8'h6 < length_2 ? _GEN_7501 : _GEN_7341; // @[executor.scala 308:60]
  wire [7:0] _GEN_7662 = 8'h6 < length_2 ? _GEN_7502 : _GEN_7342; // @[executor.scala 308:60]
  wire [7:0] _GEN_7663 = 8'h6 < length_2 ? _GEN_7503 : _GEN_7343; // @[executor.scala 308:60]
  wire [7:0] _GEN_7664 = 8'h6 < length_2 ? _GEN_7504 : _GEN_7344; // @[executor.scala 308:60]
  wire [7:0] _GEN_7665 = 8'h6 < length_2 ? _GEN_7505 : _GEN_7345; // @[executor.scala 308:60]
  wire [7:0] _GEN_7666 = 8'h6 < length_2 ? _GEN_7506 : _GEN_7346; // @[executor.scala 308:60]
  wire [7:0] _GEN_7667 = 8'h6 < length_2 ? _GEN_7507 : _GEN_7347; // @[executor.scala 308:60]
  wire [7:0] _GEN_7668 = 8'h6 < length_2 ? _GEN_7508 : _GEN_7348; // @[executor.scala 308:60]
  wire [7:0] _GEN_7669 = 8'h6 < length_2 ? _GEN_7509 : _GEN_7349; // @[executor.scala 308:60]
  wire [7:0] _GEN_7670 = 8'h6 < length_2 ? _GEN_7510 : _GEN_7350; // @[executor.scala 308:60]
  wire [7:0] _GEN_7671 = 8'h6 < length_2 ? _GEN_7511 : _GEN_7351; // @[executor.scala 308:60]
  wire [7:0] _GEN_7672 = 8'h6 < length_2 ? _GEN_7512 : _GEN_7352; // @[executor.scala 308:60]
  wire [7:0] _GEN_7673 = 8'h6 < length_2 ? _GEN_7513 : _GEN_7353; // @[executor.scala 308:60]
  wire [7:0] _GEN_7674 = 8'h6 < length_2 ? _GEN_7514 : _GEN_7354; // @[executor.scala 308:60]
  wire [7:0] _GEN_7675 = 8'h6 < length_2 ? _GEN_7515 : _GEN_7355; // @[executor.scala 308:60]
  wire [7:0] _GEN_7676 = 8'h6 < length_2 ? _GEN_7516 : _GEN_7356; // @[executor.scala 308:60]
  wire [7:0] _GEN_7677 = 8'h6 < length_2 ? _GEN_7517 : _GEN_7357; // @[executor.scala 308:60]
  wire [7:0] _GEN_7678 = 8'h6 < length_2 ? _GEN_7518 : _GEN_7358; // @[executor.scala 308:60]
  wire [7:0] _GEN_7679 = 8'h6 < length_2 ? _GEN_7519 : _GEN_7359; // @[executor.scala 308:60]
  wire [7:0] _GEN_7680 = 8'h6 < length_2 ? _GEN_7520 : _GEN_7360; // @[executor.scala 308:60]
  wire [7:0] _GEN_7681 = 8'h6 < length_2 ? _GEN_7521 : _GEN_7361; // @[executor.scala 308:60]
  wire [7:0] _GEN_7682 = 8'h6 < length_2 ? _GEN_7522 : _GEN_7362; // @[executor.scala 308:60]
  wire [7:0] _GEN_7683 = 8'h6 < length_2 ? _GEN_7523 : _GEN_7363; // @[executor.scala 308:60]
  wire [7:0] field_byte_23 = field_2[7:0]; // @[executor.scala 305:57]
  wire [7:0] total_offset_23 = offset_2 + 8'h7; // @[executor.scala 307:57]
  wire [7:0] _GEN_7684 = 8'h0 == total_offset_23 ? field_byte_23 : _GEN_7524; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7685 = 8'h1 == total_offset_23 ? field_byte_23 : _GEN_7525; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7686 = 8'h2 == total_offset_23 ? field_byte_23 : _GEN_7526; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7687 = 8'h3 == total_offset_23 ? field_byte_23 : _GEN_7527; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7688 = 8'h4 == total_offset_23 ? field_byte_23 : _GEN_7528; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7689 = 8'h5 == total_offset_23 ? field_byte_23 : _GEN_7529; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7690 = 8'h6 == total_offset_23 ? field_byte_23 : _GEN_7530; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7691 = 8'h7 == total_offset_23 ? field_byte_23 : _GEN_7531; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7692 = 8'h8 == total_offset_23 ? field_byte_23 : _GEN_7532; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7693 = 8'h9 == total_offset_23 ? field_byte_23 : _GEN_7533; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7694 = 8'ha == total_offset_23 ? field_byte_23 : _GEN_7534; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7695 = 8'hb == total_offset_23 ? field_byte_23 : _GEN_7535; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7696 = 8'hc == total_offset_23 ? field_byte_23 : _GEN_7536; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7697 = 8'hd == total_offset_23 ? field_byte_23 : _GEN_7537; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7698 = 8'he == total_offset_23 ? field_byte_23 : _GEN_7538; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7699 = 8'hf == total_offset_23 ? field_byte_23 : _GEN_7539; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7700 = 8'h10 == total_offset_23 ? field_byte_23 : _GEN_7540; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7701 = 8'h11 == total_offset_23 ? field_byte_23 : _GEN_7541; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7702 = 8'h12 == total_offset_23 ? field_byte_23 : _GEN_7542; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7703 = 8'h13 == total_offset_23 ? field_byte_23 : _GEN_7543; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7704 = 8'h14 == total_offset_23 ? field_byte_23 : _GEN_7544; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7705 = 8'h15 == total_offset_23 ? field_byte_23 : _GEN_7545; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7706 = 8'h16 == total_offset_23 ? field_byte_23 : _GEN_7546; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7707 = 8'h17 == total_offset_23 ? field_byte_23 : _GEN_7547; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7708 = 8'h18 == total_offset_23 ? field_byte_23 : _GEN_7548; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7709 = 8'h19 == total_offset_23 ? field_byte_23 : _GEN_7549; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7710 = 8'h1a == total_offset_23 ? field_byte_23 : _GEN_7550; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7711 = 8'h1b == total_offset_23 ? field_byte_23 : _GEN_7551; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7712 = 8'h1c == total_offset_23 ? field_byte_23 : _GEN_7552; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7713 = 8'h1d == total_offset_23 ? field_byte_23 : _GEN_7553; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7714 = 8'h1e == total_offset_23 ? field_byte_23 : _GEN_7554; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7715 = 8'h1f == total_offset_23 ? field_byte_23 : _GEN_7555; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7716 = 8'h20 == total_offset_23 ? field_byte_23 : _GEN_7556; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7717 = 8'h21 == total_offset_23 ? field_byte_23 : _GEN_7557; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7718 = 8'h22 == total_offset_23 ? field_byte_23 : _GEN_7558; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7719 = 8'h23 == total_offset_23 ? field_byte_23 : _GEN_7559; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7720 = 8'h24 == total_offset_23 ? field_byte_23 : _GEN_7560; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7721 = 8'h25 == total_offset_23 ? field_byte_23 : _GEN_7561; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7722 = 8'h26 == total_offset_23 ? field_byte_23 : _GEN_7562; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7723 = 8'h27 == total_offset_23 ? field_byte_23 : _GEN_7563; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7724 = 8'h28 == total_offset_23 ? field_byte_23 : _GEN_7564; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7725 = 8'h29 == total_offset_23 ? field_byte_23 : _GEN_7565; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7726 = 8'h2a == total_offset_23 ? field_byte_23 : _GEN_7566; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7727 = 8'h2b == total_offset_23 ? field_byte_23 : _GEN_7567; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7728 = 8'h2c == total_offset_23 ? field_byte_23 : _GEN_7568; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7729 = 8'h2d == total_offset_23 ? field_byte_23 : _GEN_7569; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7730 = 8'h2e == total_offset_23 ? field_byte_23 : _GEN_7570; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7731 = 8'h2f == total_offset_23 ? field_byte_23 : _GEN_7571; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7732 = 8'h30 == total_offset_23 ? field_byte_23 : _GEN_7572; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7733 = 8'h31 == total_offset_23 ? field_byte_23 : _GEN_7573; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7734 = 8'h32 == total_offset_23 ? field_byte_23 : _GEN_7574; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7735 = 8'h33 == total_offset_23 ? field_byte_23 : _GEN_7575; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7736 = 8'h34 == total_offset_23 ? field_byte_23 : _GEN_7576; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7737 = 8'h35 == total_offset_23 ? field_byte_23 : _GEN_7577; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7738 = 8'h36 == total_offset_23 ? field_byte_23 : _GEN_7578; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7739 = 8'h37 == total_offset_23 ? field_byte_23 : _GEN_7579; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7740 = 8'h38 == total_offset_23 ? field_byte_23 : _GEN_7580; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7741 = 8'h39 == total_offset_23 ? field_byte_23 : _GEN_7581; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7742 = 8'h3a == total_offset_23 ? field_byte_23 : _GEN_7582; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7743 = 8'h3b == total_offset_23 ? field_byte_23 : _GEN_7583; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7744 = 8'h3c == total_offset_23 ? field_byte_23 : _GEN_7584; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7745 = 8'h3d == total_offset_23 ? field_byte_23 : _GEN_7585; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7746 = 8'h3e == total_offset_23 ? field_byte_23 : _GEN_7586; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7747 = 8'h3f == total_offset_23 ? field_byte_23 : _GEN_7587; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7748 = 8'h40 == total_offset_23 ? field_byte_23 : _GEN_7588; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7749 = 8'h41 == total_offset_23 ? field_byte_23 : _GEN_7589; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7750 = 8'h42 == total_offset_23 ? field_byte_23 : _GEN_7590; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7751 = 8'h43 == total_offset_23 ? field_byte_23 : _GEN_7591; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7752 = 8'h44 == total_offset_23 ? field_byte_23 : _GEN_7592; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7753 = 8'h45 == total_offset_23 ? field_byte_23 : _GEN_7593; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7754 = 8'h46 == total_offset_23 ? field_byte_23 : _GEN_7594; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7755 = 8'h47 == total_offset_23 ? field_byte_23 : _GEN_7595; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7756 = 8'h48 == total_offset_23 ? field_byte_23 : _GEN_7596; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7757 = 8'h49 == total_offset_23 ? field_byte_23 : _GEN_7597; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7758 = 8'h4a == total_offset_23 ? field_byte_23 : _GEN_7598; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7759 = 8'h4b == total_offset_23 ? field_byte_23 : _GEN_7599; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7760 = 8'h4c == total_offset_23 ? field_byte_23 : _GEN_7600; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7761 = 8'h4d == total_offset_23 ? field_byte_23 : _GEN_7601; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7762 = 8'h4e == total_offset_23 ? field_byte_23 : _GEN_7602; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7763 = 8'h4f == total_offset_23 ? field_byte_23 : _GEN_7603; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7764 = 8'h50 == total_offset_23 ? field_byte_23 : _GEN_7604; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7765 = 8'h51 == total_offset_23 ? field_byte_23 : _GEN_7605; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7766 = 8'h52 == total_offset_23 ? field_byte_23 : _GEN_7606; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7767 = 8'h53 == total_offset_23 ? field_byte_23 : _GEN_7607; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7768 = 8'h54 == total_offset_23 ? field_byte_23 : _GEN_7608; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7769 = 8'h55 == total_offset_23 ? field_byte_23 : _GEN_7609; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7770 = 8'h56 == total_offset_23 ? field_byte_23 : _GEN_7610; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7771 = 8'h57 == total_offset_23 ? field_byte_23 : _GEN_7611; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7772 = 8'h58 == total_offset_23 ? field_byte_23 : _GEN_7612; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7773 = 8'h59 == total_offset_23 ? field_byte_23 : _GEN_7613; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7774 = 8'h5a == total_offset_23 ? field_byte_23 : _GEN_7614; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7775 = 8'h5b == total_offset_23 ? field_byte_23 : _GEN_7615; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7776 = 8'h5c == total_offset_23 ? field_byte_23 : _GEN_7616; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7777 = 8'h5d == total_offset_23 ? field_byte_23 : _GEN_7617; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7778 = 8'h5e == total_offset_23 ? field_byte_23 : _GEN_7618; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7779 = 8'h5f == total_offset_23 ? field_byte_23 : _GEN_7619; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7780 = 8'h60 == total_offset_23 ? field_byte_23 : _GEN_7620; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7781 = 8'h61 == total_offset_23 ? field_byte_23 : _GEN_7621; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7782 = 8'h62 == total_offset_23 ? field_byte_23 : _GEN_7622; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7783 = 8'h63 == total_offset_23 ? field_byte_23 : _GEN_7623; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7784 = 8'h64 == total_offset_23 ? field_byte_23 : _GEN_7624; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7785 = 8'h65 == total_offset_23 ? field_byte_23 : _GEN_7625; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7786 = 8'h66 == total_offset_23 ? field_byte_23 : _GEN_7626; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7787 = 8'h67 == total_offset_23 ? field_byte_23 : _GEN_7627; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7788 = 8'h68 == total_offset_23 ? field_byte_23 : _GEN_7628; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7789 = 8'h69 == total_offset_23 ? field_byte_23 : _GEN_7629; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7790 = 8'h6a == total_offset_23 ? field_byte_23 : _GEN_7630; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7791 = 8'h6b == total_offset_23 ? field_byte_23 : _GEN_7631; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7792 = 8'h6c == total_offset_23 ? field_byte_23 : _GEN_7632; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7793 = 8'h6d == total_offset_23 ? field_byte_23 : _GEN_7633; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7794 = 8'h6e == total_offset_23 ? field_byte_23 : _GEN_7634; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7795 = 8'h6f == total_offset_23 ? field_byte_23 : _GEN_7635; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7796 = 8'h70 == total_offset_23 ? field_byte_23 : _GEN_7636; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7797 = 8'h71 == total_offset_23 ? field_byte_23 : _GEN_7637; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7798 = 8'h72 == total_offset_23 ? field_byte_23 : _GEN_7638; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7799 = 8'h73 == total_offset_23 ? field_byte_23 : _GEN_7639; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7800 = 8'h74 == total_offset_23 ? field_byte_23 : _GEN_7640; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7801 = 8'h75 == total_offset_23 ? field_byte_23 : _GEN_7641; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7802 = 8'h76 == total_offset_23 ? field_byte_23 : _GEN_7642; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7803 = 8'h77 == total_offset_23 ? field_byte_23 : _GEN_7643; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7804 = 8'h78 == total_offset_23 ? field_byte_23 : _GEN_7644; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7805 = 8'h79 == total_offset_23 ? field_byte_23 : _GEN_7645; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7806 = 8'h7a == total_offset_23 ? field_byte_23 : _GEN_7646; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7807 = 8'h7b == total_offset_23 ? field_byte_23 : _GEN_7647; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7808 = 8'h7c == total_offset_23 ? field_byte_23 : _GEN_7648; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7809 = 8'h7d == total_offset_23 ? field_byte_23 : _GEN_7649; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7810 = 8'h7e == total_offset_23 ? field_byte_23 : _GEN_7650; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7811 = 8'h7f == total_offset_23 ? field_byte_23 : _GEN_7651; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7812 = 8'h80 == total_offset_23 ? field_byte_23 : _GEN_7652; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7813 = 8'h81 == total_offset_23 ? field_byte_23 : _GEN_7653; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7814 = 8'h82 == total_offset_23 ? field_byte_23 : _GEN_7654; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7815 = 8'h83 == total_offset_23 ? field_byte_23 : _GEN_7655; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7816 = 8'h84 == total_offset_23 ? field_byte_23 : _GEN_7656; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7817 = 8'h85 == total_offset_23 ? field_byte_23 : _GEN_7657; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7818 = 8'h86 == total_offset_23 ? field_byte_23 : _GEN_7658; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7819 = 8'h87 == total_offset_23 ? field_byte_23 : _GEN_7659; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7820 = 8'h88 == total_offset_23 ? field_byte_23 : _GEN_7660; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7821 = 8'h89 == total_offset_23 ? field_byte_23 : _GEN_7661; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7822 = 8'h8a == total_offset_23 ? field_byte_23 : _GEN_7662; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7823 = 8'h8b == total_offset_23 ? field_byte_23 : _GEN_7663; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7824 = 8'h8c == total_offset_23 ? field_byte_23 : _GEN_7664; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7825 = 8'h8d == total_offset_23 ? field_byte_23 : _GEN_7665; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7826 = 8'h8e == total_offset_23 ? field_byte_23 : _GEN_7666; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7827 = 8'h8f == total_offset_23 ? field_byte_23 : _GEN_7667; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7828 = 8'h90 == total_offset_23 ? field_byte_23 : _GEN_7668; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7829 = 8'h91 == total_offset_23 ? field_byte_23 : _GEN_7669; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7830 = 8'h92 == total_offset_23 ? field_byte_23 : _GEN_7670; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7831 = 8'h93 == total_offset_23 ? field_byte_23 : _GEN_7671; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7832 = 8'h94 == total_offset_23 ? field_byte_23 : _GEN_7672; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7833 = 8'h95 == total_offset_23 ? field_byte_23 : _GEN_7673; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7834 = 8'h96 == total_offset_23 ? field_byte_23 : _GEN_7674; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7835 = 8'h97 == total_offset_23 ? field_byte_23 : _GEN_7675; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7836 = 8'h98 == total_offset_23 ? field_byte_23 : _GEN_7676; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7837 = 8'h99 == total_offset_23 ? field_byte_23 : _GEN_7677; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7838 = 8'h9a == total_offset_23 ? field_byte_23 : _GEN_7678; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7839 = 8'h9b == total_offset_23 ? field_byte_23 : _GEN_7679; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7840 = 8'h9c == total_offset_23 ? field_byte_23 : _GEN_7680; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7841 = 8'h9d == total_offset_23 ? field_byte_23 : _GEN_7681; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7842 = 8'h9e == total_offset_23 ? field_byte_23 : _GEN_7682; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7843 = 8'h9f == total_offset_23 ? field_byte_23 : _GEN_7683; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_7844 = 8'h7 < length_2 ? _GEN_7684 : _GEN_7524; // @[executor.scala 308:60]
  wire [7:0] _GEN_7845 = 8'h7 < length_2 ? _GEN_7685 : _GEN_7525; // @[executor.scala 308:60]
  wire [7:0] _GEN_7846 = 8'h7 < length_2 ? _GEN_7686 : _GEN_7526; // @[executor.scala 308:60]
  wire [7:0] _GEN_7847 = 8'h7 < length_2 ? _GEN_7687 : _GEN_7527; // @[executor.scala 308:60]
  wire [7:0] _GEN_7848 = 8'h7 < length_2 ? _GEN_7688 : _GEN_7528; // @[executor.scala 308:60]
  wire [7:0] _GEN_7849 = 8'h7 < length_2 ? _GEN_7689 : _GEN_7529; // @[executor.scala 308:60]
  wire [7:0] _GEN_7850 = 8'h7 < length_2 ? _GEN_7690 : _GEN_7530; // @[executor.scala 308:60]
  wire [7:0] _GEN_7851 = 8'h7 < length_2 ? _GEN_7691 : _GEN_7531; // @[executor.scala 308:60]
  wire [7:0] _GEN_7852 = 8'h7 < length_2 ? _GEN_7692 : _GEN_7532; // @[executor.scala 308:60]
  wire [7:0] _GEN_7853 = 8'h7 < length_2 ? _GEN_7693 : _GEN_7533; // @[executor.scala 308:60]
  wire [7:0] _GEN_7854 = 8'h7 < length_2 ? _GEN_7694 : _GEN_7534; // @[executor.scala 308:60]
  wire [7:0] _GEN_7855 = 8'h7 < length_2 ? _GEN_7695 : _GEN_7535; // @[executor.scala 308:60]
  wire [7:0] _GEN_7856 = 8'h7 < length_2 ? _GEN_7696 : _GEN_7536; // @[executor.scala 308:60]
  wire [7:0] _GEN_7857 = 8'h7 < length_2 ? _GEN_7697 : _GEN_7537; // @[executor.scala 308:60]
  wire [7:0] _GEN_7858 = 8'h7 < length_2 ? _GEN_7698 : _GEN_7538; // @[executor.scala 308:60]
  wire [7:0] _GEN_7859 = 8'h7 < length_2 ? _GEN_7699 : _GEN_7539; // @[executor.scala 308:60]
  wire [7:0] _GEN_7860 = 8'h7 < length_2 ? _GEN_7700 : _GEN_7540; // @[executor.scala 308:60]
  wire [7:0] _GEN_7861 = 8'h7 < length_2 ? _GEN_7701 : _GEN_7541; // @[executor.scala 308:60]
  wire [7:0] _GEN_7862 = 8'h7 < length_2 ? _GEN_7702 : _GEN_7542; // @[executor.scala 308:60]
  wire [7:0] _GEN_7863 = 8'h7 < length_2 ? _GEN_7703 : _GEN_7543; // @[executor.scala 308:60]
  wire [7:0] _GEN_7864 = 8'h7 < length_2 ? _GEN_7704 : _GEN_7544; // @[executor.scala 308:60]
  wire [7:0] _GEN_7865 = 8'h7 < length_2 ? _GEN_7705 : _GEN_7545; // @[executor.scala 308:60]
  wire [7:0] _GEN_7866 = 8'h7 < length_2 ? _GEN_7706 : _GEN_7546; // @[executor.scala 308:60]
  wire [7:0] _GEN_7867 = 8'h7 < length_2 ? _GEN_7707 : _GEN_7547; // @[executor.scala 308:60]
  wire [7:0] _GEN_7868 = 8'h7 < length_2 ? _GEN_7708 : _GEN_7548; // @[executor.scala 308:60]
  wire [7:0] _GEN_7869 = 8'h7 < length_2 ? _GEN_7709 : _GEN_7549; // @[executor.scala 308:60]
  wire [7:0] _GEN_7870 = 8'h7 < length_2 ? _GEN_7710 : _GEN_7550; // @[executor.scala 308:60]
  wire [7:0] _GEN_7871 = 8'h7 < length_2 ? _GEN_7711 : _GEN_7551; // @[executor.scala 308:60]
  wire [7:0] _GEN_7872 = 8'h7 < length_2 ? _GEN_7712 : _GEN_7552; // @[executor.scala 308:60]
  wire [7:0] _GEN_7873 = 8'h7 < length_2 ? _GEN_7713 : _GEN_7553; // @[executor.scala 308:60]
  wire [7:0] _GEN_7874 = 8'h7 < length_2 ? _GEN_7714 : _GEN_7554; // @[executor.scala 308:60]
  wire [7:0] _GEN_7875 = 8'h7 < length_2 ? _GEN_7715 : _GEN_7555; // @[executor.scala 308:60]
  wire [7:0] _GEN_7876 = 8'h7 < length_2 ? _GEN_7716 : _GEN_7556; // @[executor.scala 308:60]
  wire [7:0] _GEN_7877 = 8'h7 < length_2 ? _GEN_7717 : _GEN_7557; // @[executor.scala 308:60]
  wire [7:0] _GEN_7878 = 8'h7 < length_2 ? _GEN_7718 : _GEN_7558; // @[executor.scala 308:60]
  wire [7:0] _GEN_7879 = 8'h7 < length_2 ? _GEN_7719 : _GEN_7559; // @[executor.scala 308:60]
  wire [7:0] _GEN_7880 = 8'h7 < length_2 ? _GEN_7720 : _GEN_7560; // @[executor.scala 308:60]
  wire [7:0] _GEN_7881 = 8'h7 < length_2 ? _GEN_7721 : _GEN_7561; // @[executor.scala 308:60]
  wire [7:0] _GEN_7882 = 8'h7 < length_2 ? _GEN_7722 : _GEN_7562; // @[executor.scala 308:60]
  wire [7:0] _GEN_7883 = 8'h7 < length_2 ? _GEN_7723 : _GEN_7563; // @[executor.scala 308:60]
  wire [7:0] _GEN_7884 = 8'h7 < length_2 ? _GEN_7724 : _GEN_7564; // @[executor.scala 308:60]
  wire [7:0] _GEN_7885 = 8'h7 < length_2 ? _GEN_7725 : _GEN_7565; // @[executor.scala 308:60]
  wire [7:0] _GEN_7886 = 8'h7 < length_2 ? _GEN_7726 : _GEN_7566; // @[executor.scala 308:60]
  wire [7:0] _GEN_7887 = 8'h7 < length_2 ? _GEN_7727 : _GEN_7567; // @[executor.scala 308:60]
  wire [7:0] _GEN_7888 = 8'h7 < length_2 ? _GEN_7728 : _GEN_7568; // @[executor.scala 308:60]
  wire [7:0] _GEN_7889 = 8'h7 < length_2 ? _GEN_7729 : _GEN_7569; // @[executor.scala 308:60]
  wire [7:0] _GEN_7890 = 8'h7 < length_2 ? _GEN_7730 : _GEN_7570; // @[executor.scala 308:60]
  wire [7:0] _GEN_7891 = 8'h7 < length_2 ? _GEN_7731 : _GEN_7571; // @[executor.scala 308:60]
  wire [7:0] _GEN_7892 = 8'h7 < length_2 ? _GEN_7732 : _GEN_7572; // @[executor.scala 308:60]
  wire [7:0] _GEN_7893 = 8'h7 < length_2 ? _GEN_7733 : _GEN_7573; // @[executor.scala 308:60]
  wire [7:0] _GEN_7894 = 8'h7 < length_2 ? _GEN_7734 : _GEN_7574; // @[executor.scala 308:60]
  wire [7:0] _GEN_7895 = 8'h7 < length_2 ? _GEN_7735 : _GEN_7575; // @[executor.scala 308:60]
  wire [7:0] _GEN_7896 = 8'h7 < length_2 ? _GEN_7736 : _GEN_7576; // @[executor.scala 308:60]
  wire [7:0] _GEN_7897 = 8'h7 < length_2 ? _GEN_7737 : _GEN_7577; // @[executor.scala 308:60]
  wire [7:0] _GEN_7898 = 8'h7 < length_2 ? _GEN_7738 : _GEN_7578; // @[executor.scala 308:60]
  wire [7:0] _GEN_7899 = 8'h7 < length_2 ? _GEN_7739 : _GEN_7579; // @[executor.scala 308:60]
  wire [7:0] _GEN_7900 = 8'h7 < length_2 ? _GEN_7740 : _GEN_7580; // @[executor.scala 308:60]
  wire [7:0] _GEN_7901 = 8'h7 < length_2 ? _GEN_7741 : _GEN_7581; // @[executor.scala 308:60]
  wire [7:0] _GEN_7902 = 8'h7 < length_2 ? _GEN_7742 : _GEN_7582; // @[executor.scala 308:60]
  wire [7:0] _GEN_7903 = 8'h7 < length_2 ? _GEN_7743 : _GEN_7583; // @[executor.scala 308:60]
  wire [7:0] _GEN_7904 = 8'h7 < length_2 ? _GEN_7744 : _GEN_7584; // @[executor.scala 308:60]
  wire [7:0] _GEN_7905 = 8'h7 < length_2 ? _GEN_7745 : _GEN_7585; // @[executor.scala 308:60]
  wire [7:0] _GEN_7906 = 8'h7 < length_2 ? _GEN_7746 : _GEN_7586; // @[executor.scala 308:60]
  wire [7:0] _GEN_7907 = 8'h7 < length_2 ? _GEN_7747 : _GEN_7587; // @[executor.scala 308:60]
  wire [7:0] _GEN_7908 = 8'h7 < length_2 ? _GEN_7748 : _GEN_7588; // @[executor.scala 308:60]
  wire [7:0] _GEN_7909 = 8'h7 < length_2 ? _GEN_7749 : _GEN_7589; // @[executor.scala 308:60]
  wire [7:0] _GEN_7910 = 8'h7 < length_2 ? _GEN_7750 : _GEN_7590; // @[executor.scala 308:60]
  wire [7:0] _GEN_7911 = 8'h7 < length_2 ? _GEN_7751 : _GEN_7591; // @[executor.scala 308:60]
  wire [7:0] _GEN_7912 = 8'h7 < length_2 ? _GEN_7752 : _GEN_7592; // @[executor.scala 308:60]
  wire [7:0] _GEN_7913 = 8'h7 < length_2 ? _GEN_7753 : _GEN_7593; // @[executor.scala 308:60]
  wire [7:0] _GEN_7914 = 8'h7 < length_2 ? _GEN_7754 : _GEN_7594; // @[executor.scala 308:60]
  wire [7:0] _GEN_7915 = 8'h7 < length_2 ? _GEN_7755 : _GEN_7595; // @[executor.scala 308:60]
  wire [7:0] _GEN_7916 = 8'h7 < length_2 ? _GEN_7756 : _GEN_7596; // @[executor.scala 308:60]
  wire [7:0] _GEN_7917 = 8'h7 < length_2 ? _GEN_7757 : _GEN_7597; // @[executor.scala 308:60]
  wire [7:0] _GEN_7918 = 8'h7 < length_2 ? _GEN_7758 : _GEN_7598; // @[executor.scala 308:60]
  wire [7:0] _GEN_7919 = 8'h7 < length_2 ? _GEN_7759 : _GEN_7599; // @[executor.scala 308:60]
  wire [7:0] _GEN_7920 = 8'h7 < length_2 ? _GEN_7760 : _GEN_7600; // @[executor.scala 308:60]
  wire [7:0] _GEN_7921 = 8'h7 < length_2 ? _GEN_7761 : _GEN_7601; // @[executor.scala 308:60]
  wire [7:0] _GEN_7922 = 8'h7 < length_2 ? _GEN_7762 : _GEN_7602; // @[executor.scala 308:60]
  wire [7:0] _GEN_7923 = 8'h7 < length_2 ? _GEN_7763 : _GEN_7603; // @[executor.scala 308:60]
  wire [7:0] _GEN_7924 = 8'h7 < length_2 ? _GEN_7764 : _GEN_7604; // @[executor.scala 308:60]
  wire [7:0] _GEN_7925 = 8'h7 < length_2 ? _GEN_7765 : _GEN_7605; // @[executor.scala 308:60]
  wire [7:0] _GEN_7926 = 8'h7 < length_2 ? _GEN_7766 : _GEN_7606; // @[executor.scala 308:60]
  wire [7:0] _GEN_7927 = 8'h7 < length_2 ? _GEN_7767 : _GEN_7607; // @[executor.scala 308:60]
  wire [7:0] _GEN_7928 = 8'h7 < length_2 ? _GEN_7768 : _GEN_7608; // @[executor.scala 308:60]
  wire [7:0] _GEN_7929 = 8'h7 < length_2 ? _GEN_7769 : _GEN_7609; // @[executor.scala 308:60]
  wire [7:0] _GEN_7930 = 8'h7 < length_2 ? _GEN_7770 : _GEN_7610; // @[executor.scala 308:60]
  wire [7:0] _GEN_7931 = 8'h7 < length_2 ? _GEN_7771 : _GEN_7611; // @[executor.scala 308:60]
  wire [7:0] _GEN_7932 = 8'h7 < length_2 ? _GEN_7772 : _GEN_7612; // @[executor.scala 308:60]
  wire [7:0] _GEN_7933 = 8'h7 < length_2 ? _GEN_7773 : _GEN_7613; // @[executor.scala 308:60]
  wire [7:0] _GEN_7934 = 8'h7 < length_2 ? _GEN_7774 : _GEN_7614; // @[executor.scala 308:60]
  wire [7:0] _GEN_7935 = 8'h7 < length_2 ? _GEN_7775 : _GEN_7615; // @[executor.scala 308:60]
  wire [7:0] _GEN_7936 = 8'h7 < length_2 ? _GEN_7776 : _GEN_7616; // @[executor.scala 308:60]
  wire [7:0] _GEN_7937 = 8'h7 < length_2 ? _GEN_7777 : _GEN_7617; // @[executor.scala 308:60]
  wire [7:0] _GEN_7938 = 8'h7 < length_2 ? _GEN_7778 : _GEN_7618; // @[executor.scala 308:60]
  wire [7:0] _GEN_7939 = 8'h7 < length_2 ? _GEN_7779 : _GEN_7619; // @[executor.scala 308:60]
  wire [7:0] _GEN_7940 = 8'h7 < length_2 ? _GEN_7780 : _GEN_7620; // @[executor.scala 308:60]
  wire [7:0] _GEN_7941 = 8'h7 < length_2 ? _GEN_7781 : _GEN_7621; // @[executor.scala 308:60]
  wire [7:0] _GEN_7942 = 8'h7 < length_2 ? _GEN_7782 : _GEN_7622; // @[executor.scala 308:60]
  wire [7:0] _GEN_7943 = 8'h7 < length_2 ? _GEN_7783 : _GEN_7623; // @[executor.scala 308:60]
  wire [7:0] _GEN_7944 = 8'h7 < length_2 ? _GEN_7784 : _GEN_7624; // @[executor.scala 308:60]
  wire [7:0] _GEN_7945 = 8'h7 < length_2 ? _GEN_7785 : _GEN_7625; // @[executor.scala 308:60]
  wire [7:0] _GEN_7946 = 8'h7 < length_2 ? _GEN_7786 : _GEN_7626; // @[executor.scala 308:60]
  wire [7:0] _GEN_7947 = 8'h7 < length_2 ? _GEN_7787 : _GEN_7627; // @[executor.scala 308:60]
  wire [7:0] _GEN_7948 = 8'h7 < length_2 ? _GEN_7788 : _GEN_7628; // @[executor.scala 308:60]
  wire [7:0] _GEN_7949 = 8'h7 < length_2 ? _GEN_7789 : _GEN_7629; // @[executor.scala 308:60]
  wire [7:0] _GEN_7950 = 8'h7 < length_2 ? _GEN_7790 : _GEN_7630; // @[executor.scala 308:60]
  wire [7:0] _GEN_7951 = 8'h7 < length_2 ? _GEN_7791 : _GEN_7631; // @[executor.scala 308:60]
  wire [7:0] _GEN_7952 = 8'h7 < length_2 ? _GEN_7792 : _GEN_7632; // @[executor.scala 308:60]
  wire [7:0] _GEN_7953 = 8'h7 < length_2 ? _GEN_7793 : _GEN_7633; // @[executor.scala 308:60]
  wire [7:0] _GEN_7954 = 8'h7 < length_2 ? _GEN_7794 : _GEN_7634; // @[executor.scala 308:60]
  wire [7:0] _GEN_7955 = 8'h7 < length_2 ? _GEN_7795 : _GEN_7635; // @[executor.scala 308:60]
  wire [7:0] _GEN_7956 = 8'h7 < length_2 ? _GEN_7796 : _GEN_7636; // @[executor.scala 308:60]
  wire [7:0] _GEN_7957 = 8'h7 < length_2 ? _GEN_7797 : _GEN_7637; // @[executor.scala 308:60]
  wire [7:0] _GEN_7958 = 8'h7 < length_2 ? _GEN_7798 : _GEN_7638; // @[executor.scala 308:60]
  wire [7:0] _GEN_7959 = 8'h7 < length_2 ? _GEN_7799 : _GEN_7639; // @[executor.scala 308:60]
  wire [7:0] _GEN_7960 = 8'h7 < length_2 ? _GEN_7800 : _GEN_7640; // @[executor.scala 308:60]
  wire [7:0] _GEN_7961 = 8'h7 < length_2 ? _GEN_7801 : _GEN_7641; // @[executor.scala 308:60]
  wire [7:0] _GEN_7962 = 8'h7 < length_2 ? _GEN_7802 : _GEN_7642; // @[executor.scala 308:60]
  wire [7:0] _GEN_7963 = 8'h7 < length_2 ? _GEN_7803 : _GEN_7643; // @[executor.scala 308:60]
  wire [7:0] _GEN_7964 = 8'h7 < length_2 ? _GEN_7804 : _GEN_7644; // @[executor.scala 308:60]
  wire [7:0] _GEN_7965 = 8'h7 < length_2 ? _GEN_7805 : _GEN_7645; // @[executor.scala 308:60]
  wire [7:0] _GEN_7966 = 8'h7 < length_2 ? _GEN_7806 : _GEN_7646; // @[executor.scala 308:60]
  wire [7:0] _GEN_7967 = 8'h7 < length_2 ? _GEN_7807 : _GEN_7647; // @[executor.scala 308:60]
  wire [7:0] _GEN_7968 = 8'h7 < length_2 ? _GEN_7808 : _GEN_7648; // @[executor.scala 308:60]
  wire [7:0] _GEN_7969 = 8'h7 < length_2 ? _GEN_7809 : _GEN_7649; // @[executor.scala 308:60]
  wire [7:0] _GEN_7970 = 8'h7 < length_2 ? _GEN_7810 : _GEN_7650; // @[executor.scala 308:60]
  wire [7:0] _GEN_7971 = 8'h7 < length_2 ? _GEN_7811 : _GEN_7651; // @[executor.scala 308:60]
  wire [7:0] _GEN_7972 = 8'h7 < length_2 ? _GEN_7812 : _GEN_7652; // @[executor.scala 308:60]
  wire [7:0] _GEN_7973 = 8'h7 < length_2 ? _GEN_7813 : _GEN_7653; // @[executor.scala 308:60]
  wire [7:0] _GEN_7974 = 8'h7 < length_2 ? _GEN_7814 : _GEN_7654; // @[executor.scala 308:60]
  wire [7:0] _GEN_7975 = 8'h7 < length_2 ? _GEN_7815 : _GEN_7655; // @[executor.scala 308:60]
  wire [7:0] _GEN_7976 = 8'h7 < length_2 ? _GEN_7816 : _GEN_7656; // @[executor.scala 308:60]
  wire [7:0] _GEN_7977 = 8'h7 < length_2 ? _GEN_7817 : _GEN_7657; // @[executor.scala 308:60]
  wire [7:0] _GEN_7978 = 8'h7 < length_2 ? _GEN_7818 : _GEN_7658; // @[executor.scala 308:60]
  wire [7:0] _GEN_7979 = 8'h7 < length_2 ? _GEN_7819 : _GEN_7659; // @[executor.scala 308:60]
  wire [7:0] _GEN_7980 = 8'h7 < length_2 ? _GEN_7820 : _GEN_7660; // @[executor.scala 308:60]
  wire [7:0] _GEN_7981 = 8'h7 < length_2 ? _GEN_7821 : _GEN_7661; // @[executor.scala 308:60]
  wire [7:0] _GEN_7982 = 8'h7 < length_2 ? _GEN_7822 : _GEN_7662; // @[executor.scala 308:60]
  wire [7:0] _GEN_7983 = 8'h7 < length_2 ? _GEN_7823 : _GEN_7663; // @[executor.scala 308:60]
  wire [7:0] _GEN_7984 = 8'h7 < length_2 ? _GEN_7824 : _GEN_7664; // @[executor.scala 308:60]
  wire [7:0] _GEN_7985 = 8'h7 < length_2 ? _GEN_7825 : _GEN_7665; // @[executor.scala 308:60]
  wire [7:0] _GEN_7986 = 8'h7 < length_2 ? _GEN_7826 : _GEN_7666; // @[executor.scala 308:60]
  wire [7:0] _GEN_7987 = 8'h7 < length_2 ? _GEN_7827 : _GEN_7667; // @[executor.scala 308:60]
  wire [7:0] _GEN_7988 = 8'h7 < length_2 ? _GEN_7828 : _GEN_7668; // @[executor.scala 308:60]
  wire [7:0] _GEN_7989 = 8'h7 < length_2 ? _GEN_7829 : _GEN_7669; // @[executor.scala 308:60]
  wire [7:0] _GEN_7990 = 8'h7 < length_2 ? _GEN_7830 : _GEN_7670; // @[executor.scala 308:60]
  wire [7:0] _GEN_7991 = 8'h7 < length_2 ? _GEN_7831 : _GEN_7671; // @[executor.scala 308:60]
  wire [7:0] _GEN_7992 = 8'h7 < length_2 ? _GEN_7832 : _GEN_7672; // @[executor.scala 308:60]
  wire [7:0] _GEN_7993 = 8'h7 < length_2 ? _GEN_7833 : _GEN_7673; // @[executor.scala 308:60]
  wire [7:0] _GEN_7994 = 8'h7 < length_2 ? _GEN_7834 : _GEN_7674; // @[executor.scala 308:60]
  wire [7:0] _GEN_7995 = 8'h7 < length_2 ? _GEN_7835 : _GEN_7675; // @[executor.scala 308:60]
  wire [7:0] _GEN_7996 = 8'h7 < length_2 ? _GEN_7836 : _GEN_7676; // @[executor.scala 308:60]
  wire [7:0] _GEN_7997 = 8'h7 < length_2 ? _GEN_7837 : _GEN_7677; // @[executor.scala 308:60]
  wire [7:0] _GEN_7998 = 8'h7 < length_2 ? _GEN_7838 : _GEN_7678; // @[executor.scala 308:60]
  wire [7:0] _GEN_7999 = 8'h7 < length_2 ? _GEN_7839 : _GEN_7679; // @[executor.scala 308:60]
  wire [7:0] _GEN_8000 = 8'h7 < length_2 ? _GEN_7840 : _GEN_7680; // @[executor.scala 308:60]
  wire [7:0] _GEN_8001 = 8'h7 < length_2 ? _GEN_7841 : _GEN_7681; // @[executor.scala 308:60]
  wire [7:0] _GEN_8002 = 8'h7 < length_2 ? _GEN_7842 : _GEN_7682; // @[executor.scala 308:60]
  wire [7:0] _GEN_8003 = 8'h7 < length_2 ? _GEN_7843 : _GEN_7683; // @[executor.scala 308:60]
  wire [3:0] _GEN_8004 = length_2 == 8'h0 ? field_2[13:10] : _GEN_5282; // @[executor.scala 300:71 executor.scala 301:55]
  wire  _GEN_8005 = length_2 == 8'h0 ? field_2[0] : _GEN_5283; // @[executor.scala 300:71 executor.scala 302:55]
  wire [7:0] _GEN_8006 = length_2 == 8'h0 ? _GEN_5284 : _GEN_7844; // @[executor.scala 300:71]
  wire [7:0] _GEN_8007 = length_2 == 8'h0 ? _GEN_5285 : _GEN_7845; // @[executor.scala 300:71]
  wire [7:0] _GEN_8008 = length_2 == 8'h0 ? _GEN_5286 : _GEN_7846; // @[executor.scala 300:71]
  wire [7:0] _GEN_8009 = length_2 == 8'h0 ? _GEN_5287 : _GEN_7847; // @[executor.scala 300:71]
  wire [7:0] _GEN_8010 = length_2 == 8'h0 ? _GEN_5288 : _GEN_7848; // @[executor.scala 300:71]
  wire [7:0] _GEN_8011 = length_2 == 8'h0 ? _GEN_5289 : _GEN_7849; // @[executor.scala 300:71]
  wire [7:0] _GEN_8012 = length_2 == 8'h0 ? _GEN_5290 : _GEN_7850; // @[executor.scala 300:71]
  wire [7:0] _GEN_8013 = length_2 == 8'h0 ? _GEN_5291 : _GEN_7851; // @[executor.scala 300:71]
  wire [7:0] _GEN_8014 = length_2 == 8'h0 ? _GEN_5292 : _GEN_7852; // @[executor.scala 300:71]
  wire [7:0] _GEN_8015 = length_2 == 8'h0 ? _GEN_5293 : _GEN_7853; // @[executor.scala 300:71]
  wire [7:0] _GEN_8016 = length_2 == 8'h0 ? _GEN_5294 : _GEN_7854; // @[executor.scala 300:71]
  wire [7:0] _GEN_8017 = length_2 == 8'h0 ? _GEN_5295 : _GEN_7855; // @[executor.scala 300:71]
  wire [7:0] _GEN_8018 = length_2 == 8'h0 ? _GEN_5296 : _GEN_7856; // @[executor.scala 300:71]
  wire [7:0] _GEN_8019 = length_2 == 8'h0 ? _GEN_5297 : _GEN_7857; // @[executor.scala 300:71]
  wire [7:0] _GEN_8020 = length_2 == 8'h0 ? _GEN_5298 : _GEN_7858; // @[executor.scala 300:71]
  wire [7:0] _GEN_8021 = length_2 == 8'h0 ? _GEN_5299 : _GEN_7859; // @[executor.scala 300:71]
  wire [7:0] _GEN_8022 = length_2 == 8'h0 ? _GEN_5300 : _GEN_7860; // @[executor.scala 300:71]
  wire [7:0] _GEN_8023 = length_2 == 8'h0 ? _GEN_5301 : _GEN_7861; // @[executor.scala 300:71]
  wire [7:0] _GEN_8024 = length_2 == 8'h0 ? _GEN_5302 : _GEN_7862; // @[executor.scala 300:71]
  wire [7:0] _GEN_8025 = length_2 == 8'h0 ? _GEN_5303 : _GEN_7863; // @[executor.scala 300:71]
  wire [7:0] _GEN_8026 = length_2 == 8'h0 ? _GEN_5304 : _GEN_7864; // @[executor.scala 300:71]
  wire [7:0] _GEN_8027 = length_2 == 8'h0 ? _GEN_5305 : _GEN_7865; // @[executor.scala 300:71]
  wire [7:0] _GEN_8028 = length_2 == 8'h0 ? _GEN_5306 : _GEN_7866; // @[executor.scala 300:71]
  wire [7:0] _GEN_8029 = length_2 == 8'h0 ? _GEN_5307 : _GEN_7867; // @[executor.scala 300:71]
  wire [7:0] _GEN_8030 = length_2 == 8'h0 ? _GEN_5308 : _GEN_7868; // @[executor.scala 300:71]
  wire [7:0] _GEN_8031 = length_2 == 8'h0 ? _GEN_5309 : _GEN_7869; // @[executor.scala 300:71]
  wire [7:0] _GEN_8032 = length_2 == 8'h0 ? _GEN_5310 : _GEN_7870; // @[executor.scala 300:71]
  wire [7:0] _GEN_8033 = length_2 == 8'h0 ? _GEN_5311 : _GEN_7871; // @[executor.scala 300:71]
  wire [7:0] _GEN_8034 = length_2 == 8'h0 ? _GEN_5312 : _GEN_7872; // @[executor.scala 300:71]
  wire [7:0] _GEN_8035 = length_2 == 8'h0 ? _GEN_5313 : _GEN_7873; // @[executor.scala 300:71]
  wire [7:0] _GEN_8036 = length_2 == 8'h0 ? _GEN_5314 : _GEN_7874; // @[executor.scala 300:71]
  wire [7:0] _GEN_8037 = length_2 == 8'h0 ? _GEN_5315 : _GEN_7875; // @[executor.scala 300:71]
  wire [7:0] _GEN_8038 = length_2 == 8'h0 ? _GEN_5316 : _GEN_7876; // @[executor.scala 300:71]
  wire [7:0] _GEN_8039 = length_2 == 8'h0 ? _GEN_5317 : _GEN_7877; // @[executor.scala 300:71]
  wire [7:0] _GEN_8040 = length_2 == 8'h0 ? _GEN_5318 : _GEN_7878; // @[executor.scala 300:71]
  wire [7:0] _GEN_8041 = length_2 == 8'h0 ? _GEN_5319 : _GEN_7879; // @[executor.scala 300:71]
  wire [7:0] _GEN_8042 = length_2 == 8'h0 ? _GEN_5320 : _GEN_7880; // @[executor.scala 300:71]
  wire [7:0] _GEN_8043 = length_2 == 8'h0 ? _GEN_5321 : _GEN_7881; // @[executor.scala 300:71]
  wire [7:0] _GEN_8044 = length_2 == 8'h0 ? _GEN_5322 : _GEN_7882; // @[executor.scala 300:71]
  wire [7:0] _GEN_8045 = length_2 == 8'h0 ? _GEN_5323 : _GEN_7883; // @[executor.scala 300:71]
  wire [7:0] _GEN_8046 = length_2 == 8'h0 ? _GEN_5324 : _GEN_7884; // @[executor.scala 300:71]
  wire [7:0] _GEN_8047 = length_2 == 8'h0 ? _GEN_5325 : _GEN_7885; // @[executor.scala 300:71]
  wire [7:0] _GEN_8048 = length_2 == 8'h0 ? _GEN_5326 : _GEN_7886; // @[executor.scala 300:71]
  wire [7:0] _GEN_8049 = length_2 == 8'h0 ? _GEN_5327 : _GEN_7887; // @[executor.scala 300:71]
  wire [7:0] _GEN_8050 = length_2 == 8'h0 ? _GEN_5328 : _GEN_7888; // @[executor.scala 300:71]
  wire [7:0] _GEN_8051 = length_2 == 8'h0 ? _GEN_5329 : _GEN_7889; // @[executor.scala 300:71]
  wire [7:0] _GEN_8052 = length_2 == 8'h0 ? _GEN_5330 : _GEN_7890; // @[executor.scala 300:71]
  wire [7:0] _GEN_8053 = length_2 == 8'h0 ? _GEN_5331 : _GEN_7891; // @[executor.scala 300:71]
  wire [7:0] _GEN_8054 = length_2 == 8'h0 ? _GEN_5332 : _GEN_7892; // @[executor.scala 300:71]
  wire [7:0] _GEN_8055 = length_2 == 8'h0 ? _GEN_5333 : _GEN_7893; // @[executor.scala 300:71]
  wire [7:0] _GEN_8056 = length_2 == 8'h0 ? _GEN_5334 : _GEN_7894; // @[executor.scala 300:71]
  wire [7:0] _GEN_8057 = length_2 == 8'h0 ? _GEN_5335 : _GEN_7895; // @[executor.scala 300:71]
  wire [7:0] _GEN_8058 = length_2 == 8'h0 ? _GEN_5336 : _GEN_7896; // @[executor.scala 300:71]
  wire [7:0] _GEN_8059 = length_2 == 8'h0 ? _GEN_5337 : _GEN_7897; // @[executor.scala 300:71]
  wire [7:0] _GEN_8060 = length_2 == 8'h0 ? _GEN_5338 : _GEN_7898; // @[executor.scala 300:71]
  wire [7:0] _GEN_8061 = length_2 == 8'h0 ? _GEN_5339 : _GEN_7899; // @[executor.scala 300:71]
  wire [7:0] _GEN_8062 = length_2 == 8'h0 ? _GEN_5340 : _GEN_7900; // @[executor.scala 300:71]
  wire [7:0] _GEN_8063 = length_2 == 8'h0 ? _GEN_5341 : _GEN_7901; // @[executor.scala 300:71]
  wire [7:0] _GEN_8064 = length_2 == 8'h0 ? _GEN_5342 : _GEN_7902; // @[executor.scala 300:71]
  wire [7:0] _GEN_8065 = length_2 == 8'h0 ? _GEN_5343 : _GEN_7903; // @[executor.scala 300:71]
  wire [7:0] _GEN_8066 = length_2 == 8'h0 ? _GEN_5344 : _GEN_7904; // @[executor.scala 300:71]
  wire [7:0] _GEN_8067 = length_2 == 8'h0 ? _GEN_5345 : _GEN_7905; // @[executor.scala 300:71]
  wire [7:0] _GEN_8068 = length_2 == 8'h0 ? _GEN_5346 : _GEN_7906; // @[executor.scala 300:71]
  wire [7:0] _GEN_8069 = length_2 == 8'h0 ? _GEN_5347 : _GEN_7907; // @[executor.scala 300:71]
  wire [7:0] _GEN_8070 = length_2 == 8'h0 ? _GEN_5348 : _GEN_7908; // @[executor.scala 300:71]
  wire [7:0] _GEN_8071 = length_2 == 8'h0 ? _GEN_5349 : _GEN_7909; // @[executor.scala 300:71]
  wire [7:0] _GEN_8072 = length_2 == 8'h0 ? _GEN_5350 : _GEN_7910; // @[executor.scala 300:71]
  wire [7:0] _GEN_8073 = length_2 == 8'h0 ? _GEN_5351 : _GEN_7911; // @[executor.scala 300:71]
  wire [7:0] _GEN_8074 = length_2 == 8'h0 ? _GEN_5352 : _GEN_7912; // @[executor.scala 300:71]
  wire [7:0] _GEN_8075 = length_2 == 8'h0 ? _GEN_5353 : _GEN_7913; // @[executor.scala 300:71]
  wire [7:0] _GEN_8076 = length_2 == 8'h0 ? _GEN_5354 : _GEN_7914; // @[executor.scala 300:71]
  wire [7:0] _GEN_8077 = length_2 == 8'h0 ? _GEN_5355 : _GEN_7915; // @[executor.scala 300:71]
  wire [7:0] _GEN_8078 = length_2 == 8'h0 ? _GEN_5356 : _GEN_7916; // @[executor.scala 300:71]
  wire [7:0] _GEN_8079 = length_2 == 8'h0 ? _GEN_5357 : _GEN_7917; // @[executor.scala 300:71]
  wire [7:0] _GEN_8080 = length_2 == 8'h0 ? _GEN_5358 : _GEN_7918; // @[executor.scala 300:71]
  wire [7:0] _GEN_8081 = length_2 == 8'h0 ? _GEN_5359 : _GEN_7919; // @[executor.scala 300:71]
  wire [7:0] _GEN_8082 = length_2 == 8'h0 ? _GEN_5360 : _GEN_7920; // @[executor.scala 300:71]
  wire [7:0] _GEN_8083 = length_2 == 8'h0 ? _GEN_5361 : _GEN_7921; // @[executor.scala 300:71]
  wire [7:0] _GEN_8084 = length_2 == 8'h0 ? _GEN_5362 : _GEN_7922; // @[executor.scala 300:71]
  wire [7:0] _GEN_8085 = length_2 == 8'h0 ? _GEN_5363 : _GEN_7923; // @[executor.scala 300:71]
  wire [7:0] _GEN_8086 = length_2 == 8'h0 ? _GEN_5364 : _GEN_7924; // @[executor.scala 300:71]
  wire [7:0] _GEN_8087 = length_2 == 8'h0 ? _GEN_5365 : _GEN_7925; // @[executor.scala 300:71]
  wire [7:0] _GEN_8088 = length_2 == 8'h0 ? _GEN_5366 : _GEN_7926; // @[executor.scala 300:71]
  wire [7:0] _GEN_8089 = length_2 == 8'h0 ? _GEN_5367 : _GEN_7927; // @[executor.scala 300:71]
  wire [7:0] _GEN_8090 = length_2 == 8'h0 ? _GEN_5368 : _GEN_7928; // @[executor.scala 300:71]
  wire [7:0] _GEN_8091 = length_2 == 8'h0 ? _GEN_5369 : _GEN_7929; // @[executor.scala 300:71]
  wire [7:0] _GEN_8092 = length_2 == 8'h0 ? _GEN_5370 : _GEN_7930; // @[executor.scala 300:71]
  wire [7:0] _GEN_8093 = length_2 == 8'h0 ? _GEN_5371 : _GEN_7931; // @[executor.scala 300:71]
  wire [7:0] _GEN_8094 = length_2 == 8'h0 ? _GEN_5372 : _GEN_7932; // @[executor.scala 300:71]
  wire [7:0] _GEN_8095 = length_2 == 8'h0 ? _GEN_5373 : _GEN_7933; // @[executor.scala 300:71]
  wire [7:0] _GEN_8096 = length_2 == 8'h0 ? _GEN_5374 : _GEN_7934; // @[executor.scala 300:71]
  wire [7:0] _GEN_8097 = length_2 == 8'h0 ? _GEN_5375 : _GEN_7935; // @[executor.scala 300:71]
  wire [7:0] _GEN_8098 = length_2 == 8'h0 ? _GEN_5376 : _GEN_7936; // @[executor.scala 300:71]
  wire [7:0] _GEN_8099 = length_2 == 8'h0 ? _GEN_5377 : _GEN_7937; // @[executor.scala 300:71]
  wire [7:0] _GEN_8100 = length_2 == 8'h0 ? _GEN_5378 : _GEN_7938; // @[executor.scala 300:71]
  wire [7:0] _GEN_8101 = length_2 == 8'h0 ? _GEN_5379 : _GEN_7939; // @[executor.scala 300:71]
  wire [7:0] _GEN_8102 = length_2 == 8'h0 ? _GEN_5380 : _GEN_7940; // @[executor.scala 300:71]
  wire [7:0] _GEN_8103 = length_2 == 8'h0 ? _GEN_5381 : _GEN_7941; // @[executor.scala 300:71]
  wire [7:0] _GEN_8104 = length_2 == 8'h0 ? _GEN_5382 : _GEN_7942; // @[executor.scala 300:71]
  wire [7:0] _GEN_8105 = length_2 == 8'h0 ? _GEN_5383 : _GEN_7943; // @[executor.scala 300:71]
  wire [7:0] _GEN_8106 = length_2 == 8'h0 ? _GEN_5384 : _GEN_7944; // @[executor.scala 300:71]
  wire [7:0] _GEN_8107 = length_2 == 8'h0 ? _GEN_5385 : _GEN_7945; // @[executor.scala 300:71]
  wire [7:0] _GEN_8108 = length_2 == 8'h0 ? _GEN_5386 : _GEN_7946; // @[executor.scala 300:71]
  wire [7:0] _GEN_8109 = length_2 == 8'h0 ? _GEN_5387 : _GEN_7947; // @[executor.scala 300:71]
  wire [7:0] _GEN_8110 = length_2 == 8'h0 ? _GEN_5388 : _GEN_7948; // @[executor.scala 300:71]
  wire [7:0] _GEN_8111 = length_2 == 8'h0 ? _GEN_5389 : _GEN_7949; // @[executor.scala 300:71]
  wire [7:0] _GEN_8112 = length_2 == 8'h0 ? _GEN_5390 : _GEN_7950; // @[executor.scala 300:71]
  wire [7:0] _GEN_8113 = length_2 == 8'h0 ? _GEN_5391 : _GEN_7951; // @[executor.scala 300:71]
  wire [7:0] _GEN_8114 = length_2 == 8'h0 ? _GEN_5392 : _GEN_7952; // @[executor.scala 300:71]
  wire [7:0] _GEN_8115 = length_2 == 8'h0 ? _GEN_5393 : _GEN_7953; // @[executor.scala 300:71]
  wire [7:0] _GEN_8116 = length_2 == 8'h0 ? _GEN_5394 : _GEN_7954; // @[executor.scala 300:71]
  wire [7:0] _GEN_8117 = length_2 == 8'h0 ? _GEN_5395 : _GEN_7955; // @[executor.scala 300:71]
  wire [7:0] _GEN_8118 = length_2 == 8'h0 ? _GEN_5396 : _GEN_7956; // @[executor.scala 300:71]
  wire [7:0] _GEN_8119 = length_2 == 8'h0 ? _GEN_5397 : _GEN_7957; // @[executor.scala 300:71]
  wire [7:0] _GEN_8120 = length_2 == 8'h0 ? _GEN_5398 : _GEN_7958; // @[executor.scala 300:71]
  wire [7:0] _GEN_8121 = length_2 == 8'h0 ? _GEN_5399 : _GEN_7959; // @[executor.scala 300:71]
  wire [7:0] _GEN_8122 = length_2 == 8'h0 ? _GEN_5400 : _GEN_7960; // @[executor.scala 300:71]
  wire [7:0] _GEN_8123 = length_2 == 8'h0 ? _GEN_5401 : _GEN_7961; // @[executor.scala 300:71]
  wire [7:0] _GEN_8124 = length_2 == 8'h0 ? _GEN_5402 : _GEN_7962; // @[executor.scala 300:71]
  wire [7:0] _GEN_8125 = length_2 == 8'h0 ? _GEN_5403 : _GEN_7963; // @[executor.scala 300:71]
  wire [7:0] _GEN_8126 = length_2 == 8'h0 ? _GEN_5404 : _GEN_7964; // @[executor.scala 300:71]
  wire [7:0] _GEN_8127 = length_2 == 8'h0 ? _GEN_5405 : _GEN_7965; // @[executor.scala 300:71]
  wire [7:0] _GEN_8128 = length_2 == 8'h0 ? _GEN_5406 : _GEN_7966; // @[executor.scala 300:71]
  wire [7:0] _GEN_8129 = length_2 == 8'h0 ? _GEN_5407 : _GEN_7967; // @[executor.scala 300:71]
  wire [7:0] _GEN_8130 = length_2 == 8'h0 ? _GEN_5408 : _GEN_7968; // @[executor.scala 300:71]
  wire [7:0] _GEN_8131 = length_2 == 8'h0 ? _GEN_5409 : _GEN_7969; // @[executor.scala 300:71]
  wire [7:0] _GEN_8132 = length_2 == 8'h0 ? _GEN_5410 : _GEN_7970; // @[executor.scala 300:71]
  wire [7:0] _GEN_8133 = length_2 == 8'h0 ? _GEN_5411 : _GEN_7971; // @[executor.scala 300:71]
  wire [7:0] _GEN_8134 = length_2 == 8'h0 ? _GEN_5412 : _GEN_7972; // @[executor.scala 300:71]
  wire [7:0] _GEN_8135 = length_2 == 8'h0 ? _GEN_5413 : _GEN_7973; // @[executor.scala 300:71]
  wire [7:0] _GEN_8136 = length_2 == 8'h0 ? _GEN_5414 : _GEN_7974; // @[executor.scala 300:71]
  wire [7:0] _GEN_8137 = length_2 == 8'h0 ? _GEN_5415 : _GEN_7975; // @[executor.scala 300:71]
  wire [7:0] _GEN_8138 = length_2 == 8'h0 ? _GEN_5416 : _GEN_7976; // @[executor.scala 300:71]
  wire [7:0] _GEN_8139 = length_2 == 8'h0 ? _GEN_5417 : _GEN_7977; // @[executor.scala 300:71]
  wire [7:0] _GEN_8140 = length_2 == 8'h0 ? _GEN_5418 : _GEN_7978; // @[executor.scala 300:71]
  wire [7:0] _GEN_8141 = length_2 == 8'h0 ? _GEN_5419 : _GEN_7979; // @[executor.scala 300:71]
  wire [7:0] _GEN_8142 = length_2 == 8'h0 ? _GEN_5420 : _GEN_7980; // @[executor.scala 300:71]
  wire [7:0] _GEN_8143 = length_2 == 8'h0 ? _GEN_5421 : _GEN_7981; // @[executor.scala 300:71]
  wire [7:0] _GEN_8144 = length_2 == 8'h0 ? _GEN_5422 : _GEN_7982; // @[executor.scala 300:71]
  wire [7:0] _GEN_8145 = length_2 == 8'h0 ? _GEN_5423 : _GEN_7983; // @[executor.scala 300:71]
  wire [7:0] _GEN_8146 = length_2 == 8'h0 ? _GEN_5424 : _GEN_7984; // @[executor.scala 300:71]
  wire [7:0] _GEN_8147 = length_2 == 8'h0 ? _GEN_5425 : _GEN_7985; // @[executor.scala 300:71]
  wire [7:0] _GEN_8148 = length_2 == 8'h0 ? _GEN_5426 : _GEN_7986; // @[executor.scala 300:71]
  wire [7:0] _GEN_8149 = length_2 == 8'h0 ? _GEN_5427 : _GEN_7987; // @[executor.scala 300:71]
  wire [7:0] _GEN_8150 = length_2 == 8'h0 ? _GEN_5428 : _GEN_7988; // @[executor.scala 300:71]
  wire [7:0] _GEN_8151 = length_2 == 8'h0 ? _GEN_5429 : _GEN_7989; // @[executor.scala 300:71]
  wire [7:0] _GEN_8152 = length_2 == 8'h0 ? _GEN_5430 : _GEN_7990; // @[executor.scala 300:71]
  wire [7:0] _GEN_8153 = length_2 == 8'h0 ? _GEN_5431 : _GEN_7991; // @[executor.scala 300:71]
  wire [7:0] _GEN_8154 = length_2 == 8'h0 ? _GEN_5432 : _GEN_7992; // @[executor.scala 300:71]
  wire [7:0] _GEN_8155 = length_2 == 8'h0 ? _GEN_5433 : _GEN_7993; // @[executor.scala 300:71]
  wire [7:0] _GEN_8156 = length_2 == 8'h0 ? _GEN_5434 : _GEN_7994; // @[executor.scala 300:71]
  wire [7:0] _GEN_8157 = length_2 == 8'h0 ? _GEN_5435 : _GEN_7995; // @[executor.scala 300:71]
  wire [7:0] _GEN_8158 = length_2 == 8'h0 ? _GEN_5436 : _GEN_7996; // @[executor.scala 300:71]
  wire [7:0] _GEN_8159 = length_2 == 8'h0 ? _GEN_5437 : _GEN_7997; // @[executor.scala 300:71]
  wire [7:0] _GEN_8160 = length_2 == 8'h0 ? _GEN_5438 : _GEN_7998; // @[executor.scala 300:71]
  wire [7:0] _GEN_8161 = length_2 == 8'h0 ? _GEN_5439 : _GEN_7999; // @[executor.scala 300:71]
  wire [7:0] _GEN_8162 = length_2 == 8'h0 ? _GEN_5440 : _GEN_8000; // @[executor.scala 300:71]
  wire [7:0] _GEN_8163 = length_2 == 8'h0 ? _GEN_5441 : _GEN_8001; // @[executor.scala 300:71]
  wire [7:0] _GEN_8164 = length_2 == 8'h0 ? _GEN_5442 : _GEN_8002; // @[executor.scala 300:71]
  wire [7:0] _GEN_8165 = length_2 == 8'h0 ? _GEN_5443 : _GEN_8003; // @[executor.scala 300:71]
  wire [7:0] field_byte_24 = field_3[63:56]; // @[executor.scala 305:57]
  wire [8:0] _total_offset_T_24 = {{1'd0}, offset_3}; // @[executor.scala 307:57]
  wire [7:0] total_offset_24 = _total_offset_T_24[7:0]; // @[executor.scala 307:57]
  wire [7:0] _GEN_8166 = 8'h0 == total_offset_24 ? field_byte_24 : _GEN_8006; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8167 = 8'h1 == total_offset_24 ? field_byte_24 : _GEN_8007; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8168 = 8'h2 == total_offset_24 ? field_byte_24 : _GEN_8008; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8169 = 8'h3 == total_offset_24 ? field_byte_24 : _GEN_8009; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8170 = 8'h4 == total_offset_24 ? field_byte_24 : _GEN_8010; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8171 = 8'h5 == total_offset_24 ? field_byte_24 : _GEN_8011; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8172 = 8'h6 == total_offset_24 ? field_byte_24 : _GEN_8012; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8173 = 8'h7 == total_offset_24 ? field_byte_24 : _GEN_8013; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8174 = 8'h8 == total_offset_24 ? field_byte_24 : _GEN_8014; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8175 = 8'h9 == total_offset_24 ? field_byte_24 : _GEN_8015; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8176 = 8'ha == total_offset_24 ? field_byte_24 : _GEN_8016; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8177 = 8'hb == total_offset_24 ? field_byte_24 : _GEN_8017; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8178 = 8'hc == total_offset_24 ? field_byte_24 : _GEN_8018; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8179 = 8'hd == total_offset_24 ? field_byte_24 : _GEN_8019; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8180 = 8'he == total_offset_24 ? field_byte_24 : _GEN_8020; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8181 = 8'hf == total_offset_24 ? field_byte_24 : _GEN_8021; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8182 = 8'h10 == total_offset_24 ? field_byte_24 : _GEN_8022; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8183 = 8'h11 == total_offset_24 ? field_byte_24 : _GEN_8023; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8184 = 8'h12 == total_offset_24 ? field_byte_24 : _GEN_8024; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8185 = 8'h13 == total_offset_24 ? field_byte_24 : _GEN_8025; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8186 = 8'h14 == total_offset_24 ? field_byte_24 : _GEN_8026; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8187 = 8'h15 == total_offset_24 ? field_byte_24 : _GEN_8027; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8188 = 8'h16 == total_offset_24 ? field_byte_24 : _GEN_8028; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8189 = 8'h17 == total_offset_24 ? field_byte_24 : _GEN_8029; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8190 = 8'h18 == total_offset_24 ? field_byte_24 : _GEN_8030; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8191 = 8'h19 == total_offset_24 ? field_byte_24 : _GEN_8031; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8192 = 8'h1a == total_offset_24 ? field_byte_24 : _GEN_8032; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8193 = 8'h1b == total_offset_24 ? field_byte_24 : _GEN_8033; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8194 = 8'h1c == total_offset_24 ? field_byte_24 : _GEN_8034; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8195 = 8'h1d == total_offset_24 ? field_byte_24 : _GEN_8035; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8196 = 8'h1e == total_offset_24 ? field_byte_24 : _GEN_8036; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8197 = 8'h1f == total_offset_24 ? field_byte_24 : _GEN_8037; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8198 = 8'h20 == total_offset_24 ? field_byte_24 : _GEN_8038; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8199 = 8'h21 == total_offset_24 ? field_byte_24 : _GEN_8039; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8200 = 8'h22 == total_offset_24 ? field_byte_24 : _GEN_8040; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8201 = 8'h23 == total_offset_24 ? field_byte_24 : _GEN_8041; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8202 = 8'h24 == total_offset_24 ? field_byte_24 : _GEN_8042; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8203 = 8'h25 == total_offset_24 ? field_byte_24 : _GEN_8043; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8204 = 8'h26 == total_offset_24 ? field_byte_24 : _GEN_8044; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8205 = 8'h27 == total_offset_24 ? field_byte_24 : _GEN_8045; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8206 = 8'h28 == total_offset_24 ? field_byte_24 : _GEN_8046; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8207 = 8'h29 == total_offset_24 ? field_byte_24 : _GEN_8047; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8208 = 8'h2a == total_offset_24 ? field_byte_24 : _GEN_8048; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8209 = 8'h2b == total_offset_24 ? field_byte_24 : _GEN_8049; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8210 = 8'h2c == total_offset_24 ? field_byte_24 : _GEN_8050; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8211 = 8'h2d == total_offset_24 ? field_byte_24 : _GEN_8051; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8212 = 8'h2e == total_offset_24 ? field_byte_24 : _GEN_8052; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8213 = 8'h2f == total_offset_24 ? field_byte_24 : _GEN_8053; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8214 = 8'h30 == total_offset_24 ? field_byte_24 : _GEN_8054; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8215 = 8'h31 == total_offset_24 ? field_byte_24 : _GEN_8055; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8216 = 8'h32 == total_offset_24 ? field_byte_24 : _GEN_8056; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8217 = 8'h33 == total_offset_24 ? field_byte_24 : _GEN_8057; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8218 = 8'h34 == total_offset_24 ? field_byte_24 : _GEN_8058; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8219 = 8'h35 == total_offset_24 ? field_byte_24 : _GEN_8059; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8220 = 8'h36 == total_offset_24 ? field_byte_24 : _GEN_8060; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8221 = 8'h37 == total_offset_24 ? field_byte_24 : _GEN_8061; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8222 = 8'h38 == total_offset_24 ? field_byte_24 : _GEN_8062; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8223 = 8'h39 == total_offset_24 ? field_byte_24 : _GEN_8063; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8224 = 8'h3a == total_offset_24 ? field_byte_24 : _GEN_8064; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8225 = 8'h3b == total_offset_24 ? field_byte_24 : _GEN_8065; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8226 = 8'h3c == total_offset_24 ? field_byte_24 : _GEN_8066; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8227 = 8'h3d == total_offset_24 ? field_byte_24 : _GEN_8067; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8228 = 8'h3e == total_offset_24 ? field_byte_24 : _GEN_8068; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8229 = 8'h3f == total_offset_24 ? field_byte_24 : _GEN_8069; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8230 = 8'h40 == total_offset_24 ? field_byte_24 : _GEN_8070; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8231 = 8'h41 == total_offset_24 ? field_byte_24 : _GEN_8071; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8232 = 8'h42 == total_offset_24 ? field_byte_24 : _GEN_8072; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8233 = 8'h43 == total_offset_24 ? field_byte_24 : _GEN_8073; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8234 = 8'h44 == total_offset_24 ? field_byte_24 : _GEN_8074; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8235 = 8'h45 == total_offset_24 ? field_byte_24 : _GEN_8075; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8236 = 8'h46 == total_offset_24 ? field_byte_24 : _GEN_8076; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8237 = 8'h47 == total_offset_24 ? field_byte_24 : _GEN_8077; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8238 = 8'h48 == total_offset_24 ? field_byte_24 : _GEN_8078; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8239 = 8'h49 == total_offset_24 ? field_byte_24 : _GEN_8079; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8240 = 8'h4a == total_offset_24 ? field_byte_24 : _GEN_8080; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8241 = 8'h4b == total_offset_24 ? field_byte_24 : _GEN_8081; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8242 = 8'h4c == total_offset_24 ? field_byte_24 : _GEN_8082; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8243 = 8'h4d == total_offset_24 ? field_byte_24 : _GEN_8083; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8244 = 8'h4e == total_offset_24 ? field_byte_24 : _GEN_8084; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8245 = 8'h4f == total_offset_24 ? field_byte_24 : _GEN_8085; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8246 = 8'h50 == total_offset_24 ? field_byte_24 : _GEN_8086; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8247 = 8'h51 == total_offset_24 ? field_byte_24 : _GEN_8087; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8248 = 8'h52 == total_offset_24 ? field_byte_24 : _GEN_8088; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8249 = 8'h53 == total_offset_24 ? field_byte_24 : _GEN_8089; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8250 = 8'h54 == total_offset_24 ? field_byte_24 : _GEN_8090; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8251 = 8'h55 == total_offset_24 ? field_byte_24 : _GEN_8091; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8252 = 8'h56 == total_offset_24 ? field_byte_24 : _GEN_8092; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8253 = 8'h57 == total_offset_24 ? field_byte_24 : _GEN_8093; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8254 = 8'h58 == total_offset_24 ? field_byte_24 : _GEN_8094; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8255 = 8'h59 == total_offset_24 ? field_byte_24 : _GEN_8095; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8256 = 8'h5a == total_offset_24 ? field_byte_24 : _GEN_8096; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8257 = 8'h5b == total_offset_24 ? field_byte_24 : _GEN_8097; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8258 = 8'h5c == total_offset_24 ? field_byte_24 : _GEN_8098; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8259 = 8'h5d == total_offset_24 ? field_byte_24 : _GEN_8099; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8260 = 8'h5e == total_offset_24 ? field_byte_24 : _GEN_8100; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8261 = 8'h5f == total_offset_24 ? field_byte_24 : _GEN_8101; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8262 = 8'h60 == total_offset_24 ? field_byte_24 : _GEN_8102; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8263 = 8'h61 == total_offset_24 ? field_byte_24 : _GEN_8103; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8264 = 8'h62 == total_offset_24 ? field_byte_24 : _GEN_8104; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8265 = 8'h63 == total_offset_24 ? field_byte_24 : _GEN_8105; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8266 = 8'h64 == total_offset_24 ? field_byte_24 : _GEN_8106; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8267 = 8'h65 == total_offset_24 ? field_byte_24 : _GEN_8107; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8268 = 8'h66 == total_offset_24 ? field_byte_24 : _GEN_8108; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8269 = 8'h67 == total_offset_24 ? field_byte_24 : _GEN_8109; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8270 = 8'h68 == total_offset_24 ? field_byte_24 : _GEN_8110; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8271 = 8'h69 == total_offset_24 ? field_byte_24 : _GEN_8111; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8272 = 8'h6a == total_offset_24 ? field_byte_24 : _GEN_8112; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8273 = 8'h6b == total_offset_24 ? field_byte_24 : _GEN_8113; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8274 = 8'h6c == total_offset_24 ? field_byte_24 : _GEN_8114; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8275 = 8'h6d == total_offset_24 ? field_byte_24 : _GEN_8115; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8276 = 8'h6e == total_offset_24 ? field_byte_24 : _GEN_8116; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8277 = 8'h6f == total_offset_24 ? field_byte_24 : _GEN_8117; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8278 = 8'h70 == total_offset_24 ? field_byte_24 : _GEN_8118; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8279 = 8'h71 == total_offset_24 ? field_byte_24 : _GEN_8119; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8280 = 8'h72 == total_offset_24 ? field_byte_24 : _GEN_8120; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8281 = 8'h73 == total_offset_24 ? field_byte_24 : _GEN_8121; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8282 = 8'h74 == total_offset_24 ? field_byte_24 : _GEN_8122; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8283 = 8'h75 == total_offset_24 ? field_byte_24 : _GEN_8123; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8284 = 8'h76 == total_offset_24 ? field_byte_24 : _GEN_8124; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8285 = 8'h77 == total_offset_24 ? field_byte_24 : _GEN_8125; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8286 = 8'h78 == total_offset_24 ? field_byte_24 : _GEN_8126; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8287 = 8'h79 == total_offset_24 ? field_byte_24 : _GEN_8127; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8288 = 8'h7a == total_offset_24 ? field_byte_24 : _GEN_8128; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8289 = 8'h7b == total_offset_24 ? field_byte_24 : _GEN_8129; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8290 = 8'h7c == total_offset_24 ? field_byte_24 : _GEN_8130; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8291 = 8'h7d == total_offset_24 ? field_byte_24 : _GEN_8131; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8292 = 8'h7e == total_offset_24 ? field_byte_24 : _GEN_8132; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8293 = 8'h7f == total_offset_24 ? field_byte_24 : _GEN_8133; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8294 = 8'h80 == total_offset_24 ? field_byte_24 : _GEN_8134; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8295 = 8'h81 == total_offset_24 ? field_byte_24 : _GEN_8135; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8296 = 8'h82 == total_offset_24 ? field_byte_24 : _GEN_8136; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8297 = 8'h83 == total_offset_24 ? field_byte_24 : _GEN_8137; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8298 = 8'h84 == total_offset_24 ? field_byte_24 : _GEN_8138; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8299 = 8'h85 == total_offset_24 ? field_byte_24 : _GEN_8139; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8300 = 8'h86 == total_offset_24 ? field_byte_24 : _GEN_8140; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8301 = 8'h87 == total_offset_24 ? field_byte_24 : _GEN_8141; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8302 = 8'h88 == total_offset_24 ? field_byte_24 : _GEN_8142; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8303 = 8'h89 == total_offset_24 ? field_byte_24 : _GEN_8143; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8304 = 8'h8a == total_offset_24 ? field_byte_24 : _GEN_8144; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8305 = 8'h8b == total_offset_24 ? field_byte_24 : _GEN_8145; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8306 = 8'h8c == total_offset_24 ? field_byte_24 : _GEN_8146; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8307 = 8'h8d == total_offset_24 ? field_byte_24 : _GEN_8147; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8308 = 8'h8e == total_offset_24 ? field_byte_24 : _GEN_8148; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8309 = 8'h8f == total_offset_24 ? field_byte_24 : _GEN_8149; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8310 = 8'h90 == total_offset_24 ? field_byte_24 : _GEN_8150; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8311 = 8'h91 == total_offset_24 ? field_byte_24 : _GEN_8151; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8312 = 8'h92 == total_offset_24 ? field_byte_24 : _GEN_8152; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8313 = 8'h93 == total_offset_24 ? field_byte_24 : _GEN_8153; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8314 = 8'h94 == total_offset_24 ? field_byte_24 : _GEN_8154; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8315 = 8'h95 == total_offset_24 ? field_byte_24 : _GEN_8155; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8316 = 8'h96 == total_offset_24 ? field_byte_24 : _GEN_8156; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8317 = 8'h97 == total_offset_24 ? field_byte_24 : _GEN_8157; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8318 = 8'h98 == total_offset_24 ? field_byte_24 : _GEN_8158; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8319 = 8'h99 == total_offset_24 ? field_byte_24 : _GEN_8159; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8320 = 8'h9a == total_offset_24 ? field_byte_24 : _GEN_8160; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8321 = 8'h9b == total_offset_24 ? field_byte_24 : _GEN_8161; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8322 = 8'h9c == total_offset_24 ? field_byte_24 : _GEN_8162; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8323 = 8'h9d == total_offset_24 ? field_byte_24 : _GEN_8163; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8324 = 8'h9e == total_offset_24 ? field_byte_24 : _GEN_8164; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8325 = 8'h9f == total_offset_24 ? field_byte_24 : _GEN_8165; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8326 = 8'h0 < length_3 ? _GEN_8166 : _GEN_8006; // @[executor.scala 308:60]
  wire [7:0] _GEN_8327 = 8'h0 < length_3 ? _GEN_8167 : _GEN_8007; // @[executor.scala 308:60]
  wire [7:0] _GEN_8328 = 8'h0 < length_3 ? _GEN_8168 : _GEN_8008; // @[executor.scala 308:60]
  wire [7:0] _GEN_8329 = 8'h0 < length_3 ? _GEN_8169 : _GEN_8009; // @[executor.scala 308:60]
  wire [7:0] _GEN_8330 = 8'h0 < length_3 ? _GEN_8170 : _GEN_8010; // @[executor.scala 308:60]
  wire [7:0] _GEN_8331 = 8'h0 < length_3 ? _GEN_8171 : _GEN_8011; // @[executor.scala 308:60]
  wire [7:0] _GEN_8332 = 8'h0 < length_3 ? _GEN_8172 : _GEN_8012; // @[executor.scala 308:60]
  wire [7:0] _GEN_8333 = 8'h0 < length_3 ? _GEN_8173 : _GEN_8013; // @[executor.scala 308:60]
  wire [7:0] _GEN_8334 = 8'h0 < length_3 ? _GEN_8174 : _GEN_8014; // @[executor.scala 308:60]
  wire [7:0] _GEN_8335 = 8'h0 < length_3 ? _GEN_8175 : _GEN_8015; // @[executor.scala 308:60]
  wire [7:0] _GEN_8336 = 8'h0 < length_3 ? _GEN_8176 : _GEN_8016; // @[executor.scala 308:60]
  wire [7:0] _GEN_8337 = 8'h0 < length_3 ? _GEN_8177 : _GEN_8017; // @[executor.scala 308:60]
  wire [7:0] _GEN_8338 = 8'h0 < length_3 ? _GEN_8178 : _GEN_8018; // @[executor.scala 308:60]
  wire [7:0] _GEN_8339 = 8'h0 < length_3 ? _GEN_8179 : _GEN_8019; // @[executor.scala 308:60]
  wire [7:0] _GEN_8340 = 8'h0 < length_3 ? _GEN_8180 : _GEN_8020; // @[executor.scala 308:60]
  wire [7:0] _GEN_8341 = 8'h0 < length_3 ? _GEN_8181 : _GEN_8021; // @[executor.scala 308:60]
  wire [7:0] _GEN_8342 = 8'h0 < length_3 ? _GEN_8182 : _GEN_8022; // @[executor.scala 308:60]
  wire [7:0] _GEN_8343 = 8'h0 < length_3 ? _GEN_8183 : _GEN_8023; // @[executor.scala 308:60]
  wire [7:0] _GEN_8344 = 8'h0 < length_3 ? _GEN_8184 : _GEN_8024; // @[executor.scala 308:60]
  wire [7:0] _GEN_8345 = 8'h0 < length_3 ? _GEN_8185 : _GEN_8025; // @[executor.scala 308:60]
  wire [7:0] _GEN_8346 = 8'h0 < length_3 ? _GEN_8186 : _GEN_8026; // @[executor.scala 308:60]
  wire [7:0] _GEN_8347 = 8'h0 < length_3 ? _GEN_8187 : _GEN_8027; // @[executor.scala 308:60]
  wire [7:0] _GEN_8348 = 8'h0 < length_3 ? _GEN_8188 : _GEN_8028; // @[executor.scala 308:60]
  wire [7:0] _GEN_8349 = 8'h0 < length_3 ? _GEN_8189 : _GEN_8029; // @[executor.scala 308:60]
  wire [7:0] _GEN_8350 = 8'h0 < length_3 ? _GEN_8190 : _GEN_8030; // @[executor.scala 308:60]
  wire [7:0] _GEN_8351 = 8'h0 < length_3 ? _GEN_8191 : _GEN_8031; // @[executor.scala 308:60]
  wire [7:0] _GEN_8352 = 8'h0 < length_3 ? _GEN_8192 : _GEN_8032; // @[executor.scala 308:60]
  wire [7:0] _GEN_8353 = 8'h0 < length_3 ? _GEN_8193 : _GEN_8033; // @[executor.scala 308:60]
  wire [7:0] _GEN_8354 = 8'h0 < length_3 ? _GEN_8194 : _GEN_8034; // @[executor.scala 308:60]
  wire [7:0] _GEN_8355 = 8'h0 < length_3 ? _GEN_8195 : _GEN_8035; // @[executor.scala 308:60]
  wire [7:0] _GEN_8356 = 8'h0 < length_3 ? _GEN_8196 : _GEN_8036; // @[executor.scala 308:60]
  wire [7:0] _GEN_8357 = 8'h0 < length_3 ? _GEN_8197 : _GEN_8037; // @[executor.scala 308:60]
  wire [7:0] _GEN_8358 = 8'h0 < length_3 ? _GEN_8198 : _GEN_8038; // @[executor.scala 308:60]
  wire [7:0] _GEN_8359 = 8'h0 < length_3 ? _GEN_8199 : _GEN_8039; // @[executor.scala 308:60]
  wire [7:0] _GEN_8360 = 8'h0 < length_3 ? _GEN_8200 : _GEN_8040; // @[executor.scala 308:60]
  wire [7:0] _GEN_8361 = 8'h0 < length_3 ? _GEN_8201 : _GEN_8041; // @[executor.scala 308:60]
  wire [7:0] _GEN_8362 = 8'h0 < length_3 ? _GEN_8202 : _GEN_8042; // @[executor.scala 308:60]
  wire [7:0] _GEN_8363 = 8'h0 < length_3 ? _GEN_8203 : _GEN_8043; // @[executor.scala 308:60]
  wire [7:0] _GEN_8364 = 8'h0 < length_3 ? _GEN_8204 : _GEN_8044; // @[executor.scala 308:60]
  wire [7:0] _GEN_8365 = 8'h0 < length_3 ? _GEN_8205 : _GEN_8045; // @[executor.scala 308:60]
  wire [7:0] _GEN_8366 = 8'h0 < length_3 ? _GEN_8206 : _GEN_8046; // @[executor.scala 308:60]
  wire [7:0] _GEN_8367 = 8'h0 < length_3 ? _GEN_8207 : _GEN_8047; // @[executor.scala 308:60]
  wire [7:0] _GEN_8368 = 8'h0 < length_3 ? _GEN_8208 : _GEN_8048; // @[executor.scala 308:60]
  wire [7:0] _GEN_8369 = 8'h0 < length_3 ? _GEN_8209 : _GEN_8049; // @[executor.scala 308:60]
  wire [7:0] _GEN_8370 = 8'h0 < length_3 ? _GEN_8210 : _GEN_8050; // @[executor.scala 308:60]
  wire [7:0] _GEN_8371 = 8'h0 < length_3 ? _GEN_8211 : _GEN_8051; // @[executor.scala 308:60]
  wire [7:0] _GEN_8372 = 8'h0 < length_3 ? _GEN_8212 : _GEN_8052; // @[executor.scala 308:60]
  wire [7:0] _GEN_8373 = 8'h0 < length_3 ? _GEN_8213 : _GEN_8053; // @[executor.scala 308:60]
  wire [7:0] _GEN_8374 = 8'h0 < length_3 ? _GEN_8214 : _GEN_8054; // @[executor.scala 308:60]
  wire [7:0] _GEN_8375 = 8'h0 < length_3 ? _GEN_8215 : _GEN_8055; // @[executor.scala 308:60]
  wire [7:0] _GEN_8376 = 8'h0 < length_3 ? _GEN_8216 : _GEN_8056; // @[executor.scala 308:60]
  wire [7:0] _GEN_8377 = 8'h0 < length_3 ? _GEN_8217 : _GEN_8057; // @[executor.scala 308:60]
  wire [7:0] _GEN_8378 = 8'h0 < length_3 ? _GEN_8218 : _GEN_8058; // @[executor.scala 308:60]
  wire [7:0] _GEN_8379 = 8'h0 < length_3 ? _GEN_8219 : _GEN_8059; // @[executor.scala 308:60]
  wire [7:0] _GEN_8380 = 8'h0 < length_3 ? _GEN_8220 : _GEN_8060; // @[executor.scala 308:60]
  wire [7:0] _GEN_8381 = 8'h0 < length_3 ? _GEN_8221 : _GEN_8061; // @[executor.scala 308:60]
  wire [7:0] _GEN_8382 = 8'h0 < length_3 ? _GEN_8222 : _GEN_8062; // @[executor.scala 308:60]
  wire [7:0] _GEN_8383 = 8'h0 < length_3 ? _GEN_8223 : _GEN_8063; // @[executor.scala 308:60]
  wire [7:0] _GEN_8384 = 8'h0 < length_3 ? _GEN_8224 : _GEN_8064; // @[executor.scala 308:60]
  wire [7:0] _GEN_8385 = 8'h0 < length_3 ? _GEN_8225 : _GEN_8065; // @[executor.scala 308:60]
  wire [7:0] _GEN_8386 = 8'h0 < length_3 ? _GEN_8226 : _GEN_8066; // @[executor.scala 308:60]
  wire [7:0] _GEN_8387 = 8'h0 < length_3 ? _GEN_8227 : _GEN_8067; // @[executor.scala 308:60]
  wire [7:0] _GEN_8388 = 8'h0 < length_3 ? _GEN_8228 : _GEN_8068; // @[executor.scala 308:60]
  wire [7:0] _GEN_8389 = 8'h0 < length_3 ? _GEN_8229 : _GEN_8069; // @[executor.scala 308:60]
  wire [7:0] _GEN_8390 = 8'h0 < length_3 ? _GEN_8230 : _GEN_8070; // @[executor.scala 308:60]
  wire [7:0] _GEN_8391 = 8'h0 < length_3 ? _GEN_8231 : _GEN_8071; // @[executor.scala 308:60]
  wire [7:0] _GEN_8392 = 8'h0 < length_3 ? _GEN_8232 : _GEN_8072; // @[executor.scala 308:60]
  wire [7:0] _GEN_8393 = 8'h0 < length_3 ? _GEN_8233 : _GEN_8073; // @[executor.scala 308:60]
  wire [7:0] _GEN_8394 = 8'h0 < length_3 ? _GEN_8234 : _GEN_8074; // @[executor.scala 308:60]
  wire [7:0] _GEN_8395 = 8'h0 < length_3 ? _GEN_8235 : _GEN_8075; // @[executor.scala 308:60]
  wire [7:0] _GEN_8396 = 8'h0 < length_3 ? _GEN_8236 : _GEN_8076; // @[executor.scala 308:60]
  wire [7:0] _GEN_8397 = 8'h0 < length_3 ? _GEN_8237 : _GEN_8077; // @[executor.scala 308:60]
  wire [7:0] _GEN_8398 = 8'h0 < length_3 ? _GEN_8238 : _GEN_8078; // @[executor.scala 308:60]
  wire [7:0] _GEN_8399 = 8'h0 < length_3 ? _GEN_8239 : _GEN_8079; // @[executor.scala 308:60]
  wire [7:0] _GEN_8400 = 8'h0 < length_3 ? _GEN_8240 : _GEN_8080; // @[executor.scala 308:60]
  wire [7:0] _GEN_8401 = 8'h0 < length_3 ? _GEN_8241 : _GEN_8081; // @[executor.scala 308:60]
  wire [7:0] _GEN_8402 = 8'h0 < length_3 ? _GEN_8242 : _GEN_8082; // @[executor.scala 308:60]
  wire [7:0] _GEN_8403 = 8'h0 < length_3 ? _GEN_8243 : _GEN_8083; // @[executor.scala 308:60]
  wire [7:0] _GEN_8404 = 8'h0 < length_3 ? _GEN_8244 : _GEN_8084; // @[executor.scala 308:60]
  wire [7:0] _GEN_8405 = 8'h0 < length_3 ? _GEN_8245 : _GEN_8085; // @[executor.scala 308:60]
  wire [7:0] _GEN_8406 = 8'h0 < length_3 ? _GEN_8246 : _GEN_8086; // @[executor.scala 308:60]
  wire [7:0] _GEN_8407 = 8'h0 < length_3 ? _GEN_8247 : _GEN_8087; // @[executor.scala 308:60]
  wire [7:0] _GEN_8408 = 8'h0 < length_3 ? _GEN_8248 : _GEN_8088; // @[executor.scala 308:60]
  wire [7:0] _GEN_8409 = 8'h0 < length_3 ? _GEN_8249 : _GEN_8089; // @[executor.scala 308:60]
  wire [7:0] _GEN_8410 = 8'h0 < length_3 ? _GEN_8250 : _GEN_8090; // @[executor.scala 308:60]
  wire [7:0] _GEN_8411 = 8'h0 < length_3 ? _GEN_8251 : _GEN_8091; // @[executor.scala 308:60]
  wire [7:0] _GEN_8412 = 8'h0 < length_3 ? _GEN_8252 : _GEN_8092; // @[executor.scala 308:60]
  wire [7:0] _GEN_8413 = 8'h0 < length_3 ? _GEN_8253 : _GEN_8093; // @[executor.scala 308:60]
  wire [7:0] _GEN_8414 = 8'h0 < length_3 ? _GEN_8254 : _GEN_8094; // @[executor.scala 308:60]
  wire [7:0] _GEN_8415 = 8'h0 < length_3 ? _GEN_8255 : _GEN_8095; // @[executor.scala 308:60]
  wire [7:0] _GEN_8416 = 8'h0 < length_3 ? _GEN_8256 : _GEN_8096; // @[executor.scala 308:60]
  wire [7:0] _GEN_8417 = 8'h0 < length_3 ? _GEN_8257 : _GEN_8097; // @[executor.scala 308:60]
  wire [7:0] _GEN_8418 = 8'h0 < length_3 ? _GEN_8258 : _GEN_8098; // @[executor.scala 308:60]
  wire [7:0] _GEN_8419 = 8'h0 < length_3 ? _GEN_8259 : _GEN_8099; // @[executor.scala 308:60]
  wire [7:0] _GEN_8420 = 8'h0 < length_3 ? _GEN_8260 : _GEN_8100; // @[executor.scala 308:60]
  wire [7:0] _GEN_8421 = 8'h0 < length_3 ? _GEN_8261 : _GEN_8101; // @[executor.scala 308:60]
  wire [7:0] _GEN_8422 = 8'h0 < length_3 ? _GEN_8262 : _GEN_8102; // @[executor.scala 308:60]
  wire [7:0] _GEN_8423 = 8'h0 < length_3 ? _GEN_8263 : _GEN_8103; // @[executor.scala 308:60]
  wire [7:0] _GEN_8424 = 8'h0 < length_3 ? _GEN_8264 : _GEN_8104; // @[executor.scala 308:60]
  wire [7:0] _GEN_8425 = 8'h0 < length_3 ? _GEN_8265 : _GEN_8105; // @[executor.scala 308:60]
  wire [7:0] _GEN_8426 = 8'h0 < length_3 ? _GEN_8266 : _GEN_8106; // @[executor.scala 308:60]
  wire [7:0] _GEN_8427 = 8'h0 < length_3 ? _GEN_8267 : _GEN_8107; // @[executor.scala 308:60]
  wire [7:0] _GEN_8428 = 8'h0 < length_3 ? _GEN_8268 : _GEN_8108; // @[executor.scala 308:60]
  wire [7:0] _GEN_8429 = 8'h0 < length_3 ? _GEN_8269 : _GEN_8109; // @[executor.scala 308:60]
  wire [7:0] _GEN_8430 = 8'h0 < length_3 ? _GEN_8270 : _GEN_8110; // @[executor.scala 308:60]
  wire [7:0] _GEN_8431 = 8'h0 < length_3 ? _GEN_8271 : _GEN_8111; // @[executor.scala 308:60]
  wire [7:0] _GEN_8432 = 8'h0 < length_3 ? _GEN_8272 : _GEN_8112; // @[executor.scala 308:60]
  wire [7:0] _GEN_8433 = 8'h0 < length_3 ? _GEN_8273 : _GEN_8113; // @[executor.scala 308:60]
  wire [7:0] _GEN_8434 = 8'h0 < length_3 ? _GEN_8274 : _GEN_8114; // @[executor.scala 308:60]
  wire [7:0] _GEN_8435 = 8'h0 < length_3 ? _GEN_8275 : _GEN_8115; // @[executor.scala 308:60]
  wire [7:0] _GEN_8436 = 8'h0 < length_3 ? _GEN_8276 : _GEN_8116; // @[executor.scala 308:60]
  wire [7:0] _GEN_8437 = 8'h0 < length_3 ? _GEN_8277 : _GEN_8117; // @[executor.scala 308:60]
  wire [7:0] _GEN_8438 = 8'h0 < length_3 ? _GEN_8278 : _GEN_8118; // @[executor.scala 308:60]
  wire [7:0] _GEN_8439 = 8'h0 < length_3 ? _GEN_8279 : _GEN_8119; // @[executor.scala 308:60]
  wire [7:0] _GEN_8440 = 8'h0 < length_3 ? _GEN_8280 : _GEN_8120; // @[executor.scala 308:60]
  wire [7:0] _GEN_8441 = 8'h0 < length_3 ? _GEN_8281 : _GEN_8121; // @[executor.scala 308:60]
  wire [7:0] _GEN_8442 = 8'h0 < length_3 ? _GEN_8282 : _GEN_8122; // @[executor.scala 308:60]
  wire [7:0] _GEN_8443 = 8'h0 < length_3 ? _GEN_8283 : _GEN_8123; // @[executor.scala 308:60]
  wire [7:0] _GEN_8444 = 8'h0 < length_3 ? _GEN_8284 : _GEN_8124; // @[executor.scala 308:60]
  wire [7:0] _GEN_8445 = 8'h0 < length_3 ? _GEN_8285 : _GEN_8125; // @[executor.scala 308:60]
  wire [7:0] _GEN_8446 = 8'h0 < length_3 ? _GEN_8286 : _GEN_8126; // @[executor.scala 308:60]
  wire [7:0] _GEN_8447 = 8'h0 < length_3 ? _GEN_8287 : _GEN_8127; // @[executor.scala 308:60]
  wire [7:0] _GEN_8448 = 8'h0 < length_3 ? _GEN_8288 : _GEN_8128; // @[executor.scala 308:60]
  wire [7:0] _GEN_8449 = 8'h0 < length_3 ? _GEN_8289 : _GEN_8129; // @[executor.scala 308:60]
  wire [7:0] _GEN_8450 = 8'h0 < length_3 ? _GEN_8290 : _GEN_8130; // @[executor.scala 308:60]
  wire [7:0] _GEN_8451 = 8'h0 < length_3 ? _GEN_8291 : _GEN_8131; // @[executor.scala 308:60]
  wire [7:0] _GEN_8452 = 8'h0 < length_3 ? _GEN_8292 : _GEN_8132; // @[executor.scala 308:60]
  wire [7:0] _GEN_8453 = 8'h0 < length_3 ? _GEN_8293 : _GEN_8133; // @[executor.scala 308:60]
  wire [7:0] _GEN_8454 = 8'h0 < length_3 ? _GEN_8294 : _GEN_8134; // @[executor.scala 308:60]
  wire [7:0] _GEN_8455 = 8'h0 < length_3 ? _GEN_8295 : _GEN_8135; // @[executor.scala 308:60]
  wire [7:0] _GEN_8456 = 8'h0 < length_3 ? _GEN_8296 : _GEN_8136; // @[executor.scala 308:60]
  wire [7:0] _GEN_8457 = 8'h0 < length_3 ? _GEN_8297 : _GEN_8137; // @[executor.scala 308:60]
  wire [7:0] _GEN_8458 = 8'h0 < length_3 ? _GEN_8298 : _GEN_8138; // @[executor.scala 308:60]
  wire [7:0] _GEN_8459 = 8'h0 < length_3 ? _GEN_8299 : _GEN_8139; // @[executor.scala 308:60]
  wire [7:0] _GEN_8460 = 8'h0 < length_3 ? _GEN_8300 : _GEN_8140; // @[executor.scala 308:60]
  wire [7:0] _GEN_8461 = 8'h0 < length_3 ? _GEN_8301 : _GEN_8141; // @[executor.scala 308:60]
  wire [7:0] _GEN_8462 = 8'h0 < length_3 ? _GEN_8302 : _GEN_8142; // @[executor.scala 308:60]
  wire [7:0] _GEN_8463 = 8'h0 < length_3 ? _GEN_8303 : _GEN_8143; // @[executor.scala 308:60]
  wire [7:0] _GEN_8464 = 8'h0 < length_3 ? _GEN_8304 : _GEN_8144; // @[executor.scala 308:60]
  wire [7:0] _GEN_8465 = 8'h0 < length_3 ? _GEN_8305 : _GEN_8145; // @[executor.scala 308:60]
  wire [7:0] _GEN_8466 = 8'h0 < length_3 ? _GEN_8306 : _GEN_8146; // @[executor.scala 308:60]
  wire [7:0] _GEN_8467 = 8'h0 < length_3 ? _GEN_8307 : _GEN_8147; // @[executor.scala 308:60]
  wire [7:0] _GEN_8468 = 8'h0 < length_3 ? _GEN_8308 : _GEN_8148; // @[executor.scala 308:60]
  wire [7:0] _GEN_8469 = 8'h0 < length_3 ? _GEN_8309 : _GEN_8149; // @[executor.scala 308:60]
  wire [7:0] _GEN_8470 = 8'h0 < length_3 ? _GEN_8310 : _GEN_8150; // @[executor.scala 308:60]
  wire [7:0] _GEN_8471 = 8'h0 < length_3 ? _GEN_8311 : _GEN_8151; // @[executor.scala 308:60]
  wire [7:0] _GEN_8472 = 8'h0 < length_3 ? _GEN_8312 : _GEN_8152; // @[executor.scala 308:60]
  wire [7:0] _GEN_8473 = 8'h0 < length_3 ? _GEN_8313 : _GEN_8153; // @[executor.scala 308:60]
  wire [7:0] _GEN_8474 = 8'h0 < length_3 ? _GEN_8314 : _GEN_8154; // @[executor.scala 308:60]
  wire [7:0] _GEN_8475 = 8'h0 < length_3 ? _GEN_8315 : _GEN_8155; // @[executor.scala 308:60]
  wire [7:0] _GEN_8476 = 8'h0 < length_3 ? _GEN_8316 : _GEN_8156; // @[executor.scala 308:60]
  wire [7:0] _GEN_8477 = 8'h0 < length_3 ? _GEN_8317 : _GEN_8157; // @[executor.scala 308:60]
  wire [7:0] _GEN_8478 = 8'h0 < length_3 ? _GEN_8318 : _GEN_8158; // @[executor.scala 308:60]
  wire [7:0] _GEN_8479 = 8'h0 < length_3 ? _GEN_8319 : _GEN_8159; // @[executor.scala 308:60]
  wire [7:0] _GEN_8480 = 8'h0 < length_3 ? _GEN_8320 : _GEN_8160; // @[executor.scala 308:60]
  wire [7:0] _GEN_8481 = 8'h0 < length_3 ? _GEN_8321 : _GEN_8161; // @[executor.scala 308:60]
  wire [7:0] _GEN_8482 = 8'h0 < length_3 ? _GEN_8322 : _GEN_8162; // @[executor.scala 308:60]
  wire [7:0] _GEN_8483 = 8'h0 < length_3 ? _GEN_8323 : _GEN_8163; // @[executor.scala 308:60]
  wire [7:0] _GEN_8484 = 8'h0 < length_3 ? _GEN_8324 : _GEN_8164; // @[executor.scala 308:60]
  wire [7:0] _GEN_8485 = 8'h0 < length_3 ? _GEN_8325 : _GEN_8165; // @[executor.scala 308:60]
  wire [7:0] field_byte_25 = field_3[55:48]; // @[executor.scala 305:57]
  wire [7:0] total_offset_25 = offset_3 + 8'h1; // @[executor.scala 307:57]
  wire [7:0] _GEN_8486 = 8'h0 == total_offset_25 ? field_byte_25 : _GEN_8326; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8487 = 8'h1 == total_offset_25 ? field_byte_25 : _GEN_8327; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8488 = 8'h2 == total_offset_25 ? field_byte_25 : _GEN_8328; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8489 = 8'h3 == total_offset_25 ? field_byte_25 : _GEN_8329; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8490 = 8'h4 == total_offset_25 ? field_byte_25 : _GEN_8330; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8491 = 8'h5 == total_offset_25 ? field_byte_25 : _GEN_8331; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8492 = 8'h6 == total_offset_25 ? field_byte_25 : _GEN_8332; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8493 = 8'h7 == total_offset_25 ? field_byte_25 : _GEN_8333; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8494 = 8'h8 == total_offset_25 ? field_byte_25 : _GEN_8334; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8495 = 8'h9 == total_offset_25 ? field_byte_25 : _GEN_8335; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8496 = 8'ha == total_offset_25 ? field_byte_25 : _GEN_8336; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8497 = 8'hb == total_offset_25 ? field_byte_25 : _GEN_8337; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8498 = 8'hc == total_offset_25 ? field_byte_25 : _GEN_8338; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8499 = 8'hd == total_offset_25 ? field_byte_25 : _GEN_8339; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8500 = 8'he == total_offset_25 ? field_byte_25 : _GEN_8340; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8501 = 8'hf == total_offset_25 ? field_byte_25 : _GEN_8341; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8502 = 8'h10 == total_offset_25 ? field_byte_25 : _GEN_8342; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8503 = 8'h11 == total_offset_25 ? field_byte_25 : _GEN_8343; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8504 = 8'h12 == total_offset_25 ? field_byte_25 : _GEN_8344; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8505 = 8'h13 == total_offset_25 ? field_byte_25 : _GEN_8345; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8506 = 8'h14 == total_offset_25 ? field_byte_25 : _GEN_8346; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8507 = 8'h15 == total_offset_25 ? field_byte_25 : _GEN_8347; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8508 = 8'h16 == total_offset_25 ? field_byte_25 : _GEN_8348; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8509 = 8'h17 == total_offset_25 ? field_byte_25 : _GEN_8349; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8510 = 8'h18 == total_offset_25 ? field_byte_25 : _GEN_8350; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8511 = 8'h19 == total_offset_25 ? field_byte_25 : _GEN_8351; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8512 = 8'h1a == total_offset_25 ? field_byte_25 : _GEN_8352; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8513 = 8'h1b == total_offset_25 ? field_byte_25 : _GEN_8353; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8514 = 8'h1c == total_offset_25 ? field_byte_25 : _GEN_8354; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8515 = 8'h1d == total_offset_25 ? field_byte_25 : _GEN_8355; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8516 = 8'h1e == total_offset_25 ? field_byte_25 : _GEN_8356; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8517 = 8'h1f == total_offset_25 ? field_byte_25 : _GEN_8357; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8518 = 8'h20 == total_offset_25 ? field_byte_25 : _GEN_8358; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8519 = 8'h21 == total_offset_25 ? field_byte_25 : _GEN_8359; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8520 = 8'h22 == total_offset_25 ? field_byte_25 : _GEN_8360; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8521 = 8'h23 == total_offset_25 ? field_byte_25 : _GEN_8361; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8522 = 8'h24 == total_offset_25 ? field_byte_25 : _GEN_8362; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8523 = 8'h25 == total_offset_25 ? field_byte_25 : _GEN_8363; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8524 = 8'h26 == total_offset_25 ? field_byte_25 : _GEN_8364; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8525 = 8'h27 == total_offset_25 ? field_byte_25 : _GEN_8365; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8526 = 8'h28 == total_offset_25 ? field_byte_25 : _GEN_8366; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8527 = 8'h29 == total_offset_25 ? field_byte_25 : _GEN_8367; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8528 = 8'h2a == total_offset_25 ? field_byte_25 : _GEN_8368; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8529 = 8'h2b == total_offset_25 ? field_byte_25 : _GEN_8369; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8530 = 8'h2c == total_offset_25 ? field_byte_25 : _GEN_8370; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8531 = 8'h2d == total_offset_25 ? field_byte_25 : _GEN_8371; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8532 = 8'h2e == total_offset_25 ? field_byte_25 : _GEN_8372; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8533 = 8'h2f == total_offset_25 ? field_byte_25 : _GEN_8373; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8534 = 8'h30 == total_offset_25 ? field_byte_25 : _GEN_8374; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8535 = 8'h31 == total_offset_25 ? field_byte_25 : _GEN_8375; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8536 = 8'h32 == total_offset_25 ? field_byte_25 : _GEN_8376; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8537 = 8'h33 == total_offset_25 ? field_byte_25 : _GEN_8377; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8538 = 8'h34 == total_offset_25 ? field_byte_25 : _GEN_8378; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8539 = 8'h35 == total_offset_25 ? field_byte_25 : _GEN_8379; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8540 = 8'h36 == total_offset_25 ? field_byte_25 : _GEN_8380; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8541 = 8'h37 == total_offset_25 ? field_byte_25 : _GEN_8381; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8542 = 8'h38 == total_offset_25 ? field_byte_25 : _GEN_8382; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8543 = 8'h39 == total_offset_25 ? field_byte_25 : _GEN_8383; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8544 = 8'h3a == total_offset_25 ? field_byte_25 : _GEN_8384; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8545 = 8'h3b == total_offset_25 ? field_byte_25 : _GEN_8385; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8546 = 8'h3c == total_offset_25 ? field_byte_25 : _GEN_8386; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8547 = 8'h3d == total_offset_25 ? field_byte_25 : _GEN_8387; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8548 = 8'h3e == total_offset_25 ? field_byte_25 : _GEN_8388; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8549 = 8'h3f == total_offset_25 ? field_byte_25 : _GEN_8389; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8550 = 8'h40 == total_offset_25 ? field_byte_25 : _GEN_8390; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8551 = 8'h41 == total_offset_25 ? field_byte_25 : _GEN_8391; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8552 = 8'h42 == total_offset_25 ? field_byte_25 : _GEN_8392; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8553 = 8'h43 == total_offset_25 ? field_byte_25 : _GEN_8393; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8554 = 8'h44 == total_offset_25 ? field_byte_25 : _GEN_8394; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8555 = 8'h45 == total_offset_25 ? field_byte_25 : _GEN_8395; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8556 = 8'h46 == total_offset_25 ? field_byte_25 : _GEN_8396; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8557 = 8'h47 == total_offset_25 ? field_byte_25 : _GEN_8397; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8558 = 8'h48 == total_offset_25 ? field_byte_25 : _GEN_8398; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8559 = 8'h49 == total_offset_25 ? field_byte_25 : _GEN_8399; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8560 = 8'h4a == total_offset_25 ? field_byte_25 : _GEN_8400; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8561 = 8'h4b == total_offset_25 ? field_byte_25 : _GEN_8401; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8562 = 8'h4c == total_offset_25 ? field_byte_25 : _GEN_8402; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8563 = 8'h4d == total_offset_25 ? field_byte_25 : _GEN_8403; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8564 = 8'h4e == total_offset_25 ? field_byte_25 : _GEN_8404; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8565 = 8'h4f == total_offset_25 ? field_byte_25 : _GEN_8405; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8566 = 8'h50 == total_offset_25 ? field_byte_25 : _GEN_8406; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8567 = 8'h51 == total_offset_25 ? field_byte_25 : _GEN_8407; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8568 = 8'h52 == total_offset_25 ? field_byte_25 : _GEN_8408; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8569 = 8'h53 == total_offset_25 ? field_byte_25 : _GEN_8409; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8570 = 8'h54 == total_offset_25 ? field_byte_25 : _GEN_8410; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8571 = 8'h55 == total_offset_25 ? field_byte_25 : _GEN_8411; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8572 = 8'h56 == total_offset_25 ? field_byte_25 : _GEN_8412; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8573 = 8'h57 == total_offset_25 ? field_byte_25 : _GEN_8413; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8574 = 8'h58 == total_offset_25 ? field_byte_25 : _GEN_8414; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8575 = 8'h59 == total_offset_25 ? field_byte_25 : _GEN_8415; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8576 = 8'h5a == total_offset_25 ? field_byte_25 : _GEN_8416; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8577 = 8'h5b == total_offset_25 ? field_byte_25 : _GEN_8417; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8578 = 8'h5c == total_offset_25 ? field_byte_25 : _GEN_8418; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8579 = 8'h5d == total_offset_25 ? field_byte_25 : _GEN_8419; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8580 = 8'h5e == total_offset_25 ? field_byte_25 : _GEN_8420; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8581 = 8'h5f == total_offset_25 ? field_byte_25 : _GEN_8421; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8582 = 8'h60 == total_offset_25 ? field_byte_25 : _GEN_8422; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8583 = 8'h61 == total_offset_25 ? field_byte_25 : _GEN_8423; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8584 = 8'h62 == total_offset_25 ? field_byte_25 : _GEN_8424; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8585 = 8'h63 == total_offset_25 ? field_byte_25 : _GEN_8425; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8586 = 8'h64 == total_offset_25 ? field_byte_25 : _GEN_8426; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8587 = 8'h65 == total_offset_25 ? field_byte_25 : _GEN_8427; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8588 = 8'h66 == total_offset_25 ? field_byte_25 : _GEN_8428; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8589 = 8'h67 == total_offset_25 ? field_byte_25 : _GEN_8429; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8590 = 8'h68 == total_offset_25 ? field_byte_25 : _GEN_8430; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8591 = 8'h69 == total_offset_25 ? field_byte_25 : _GEN_8431; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8592 = 8'h6a == total_offset_25 ? field_byte_25 : _GEN_8432; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8593 = 8'h6b == total_offset_25 ? field_byte_25 : _GEN_8433; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8594 = 8'h6c == total_offset_25 ? field_byte_25 : _GEN_8434; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8595 = 8'h6d == total_offset_25 ? field_byte_25 : _GEN_8435; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8596 = 8'h6e == total_offset_25 ? field_byte_25 : _GEN_8436; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8597 = 8'h6f == total_offset_25 ? field_byte_25 : _GEN_8437; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8598 = 8'h70 == total_offset_25 ? field_byte_25 : _GEN_8438; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8599 = 8'h71 == total_offset_25 ? field_byte_25 : _GEN_8439; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8600 = 8'h72 == total_offset_25 ? field_byte_25 : _GEN_8440; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8601 = 8'h73 == total_offset_25 ? field_byte_25 : _GEN_8441; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8602 = 8'h74 == total_offset_25 ? field_byte_25 : _GEN_8442; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8603 = 8'h75 == total_offset_25 ? field_byte_25 : _GEN_8443; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8604 = 8'h76 == total_offset_25 ? field_byte_25 : _GEN_8444; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8605 = 8'h77 == total_offset_25 ? field_byte_25 : _GEN_8445; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8606 = 8'h78 == total_offset_25 ? field_byte_25 : _GEN_8446; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8607 = 8'h79 == total_offset_25 ? field_byte_25 : _GEN_8447; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8608 = 8'h7a == total_offset_25 ? field_byte_25 : _GEN_8448; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8609 = 8'h7b == total_offset_25 ? field_byte_25 : _GEN_8449; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8610 = 8'h7c == total_offset_25 ? field_byte_25 : _GEN_8450; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8611 = 8'h7d == total_offset_25 ? field_byte_25 : _GEN_8451; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8612 = 8'h7e == total_offset_25 ? field_byte_25 : _GEN_8452; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8613 = 8'h7f == total_offset_25 ? field_byte_25 : _GEN_8453; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8614 = 8'h80 == total_offset_25 ? field_byte_25 : _GEN_8454; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8615 = 8'h81 == total_offset_25 ? field_byte_25 : _GEN_8455; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8616 = 8'h82 == total_offset_25 ? field_byte_25 : _GEN_8456; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8617 = 8'h83 == total_offset_25 ? field_byte_25 : _GEN_8457; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8618 = 8'h84 == total_offset_25 ? field_byte_25 : _GEN_8458; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8619 = 8'h85 == total_offset_25 ? field_byte_25 : _GEN_8459; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8620 = 8'h86 == total_offset_25 ? field_byte_25 : _GEN_8460; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8621 = 8'h87 == total_offset_25 ? field_byte_25 : _GEN_8461; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8622 = 8'h88 == total_offset_25 ? field_byte_25 : _GEN_8462; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8623 = 8'h89 == total_offset_25 ? field_byte_25 : _GEN_8463; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8624 = 8'h8a == total_offset_25 ? field_byte_25 : _GEN_8464; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8625 = 8'h8b == total_offset_25 ? field_byte_25 : _GEN_8465; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8626 = 8'h8c == total_offset_25 ? field_byte_25 : _GEN_8466; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8627 = 8'h8d == total_offset_25 ? field_byte_25 : _GEN_8467; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8628 = 8'h8e == total_offset_25 ? field_byte_25 : _GEN_8468; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8629 = 8'h8f == total_offset_25 ? field_byte_25 : _GEN_8469; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8630 = 8'h90 == total_offset_25 ? field_byte_25 : _GEN_8470; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8631 = 8'h91 == total_offset_25 ? field_byte_25 : _GEN_8471; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8632 = 8'h92 == total_offset_25 ? field_byte_25 : _GEN_8472; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8633 = 8'h93 == total_offset_25 ? field_byte_25 : _GEN_8473; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8634 = 8'h94 == total_offset_25 ? field_byte_25 : _GEN_8474; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8635 = 8'h95 == total_offset_25 ? field_byte_25 : _GEN_8475; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8636 = 8'h96 == total_offset_25 ? field_byte_25 : _GEN_8476; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8637 = 8'h97 == total_offset_25 ? field_byte_25 : _GEN_8477; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8638 = 8'h98 == total_offset_25 ? field_byte_25 : _GEN_8478; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8639 = 8'h99 == total_offset_25 ? field_byte_25 : _GEN_8479; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8640 = 8'h9a == total_offset_25 ? field_byte_25 : _GEN_8480; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8641 = 8'h9b == total_offset_25 ? field_byte_25 : _GEN_8481; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8642 = 8'h9c == total_offset_25 ? field_byte_25 : _GEN_8482; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8643 = 8'h9d == total_offset_25 ? field_byte_25 : _GEN_8483; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8644 = 8'h9e == total_offset_25 ? field_byte_25 : _GEN_8484; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8645 = 8'h9f == total_offset_25 ? field_byte_25 : _GEN_8485; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8646 = 8'h1 < length_3 ? _GEN_8486 : _GEN_8326; // @[executor.scala 308:60]
  wire [7:0] _GEN_8647 = 8'h1 < length_3 ? _GEN_8487 : _GEN_8327; // @[executor.scala 308:60]
  wire [7:0] _GEN_8648 = 8'h1 < length_3 ? _GEN_8488 : _GEN_8328; // @[executor.scala 308:60]
  wire [7:0] _GEN_8649 = 8'h1 < length_3 ? _GEN_8489 : _GEN_8329; // @[executor.scala 308:60]
  wire [7:0] _GEN_8650 = 8'h1 < length_3 ? _GEN_8490 : _GEN_8330; // @[executor.scala 308:60]
  wire [7:0] _GEN_8651 = 8'h1 < length_3 ? _GEN_8491 : _GEN_8331; // @[executor.scala 308:60]
  wire [7:0] _GEN_8652 = 8'h1 < length_3 ? _GEN_8492 : _GEN_8332; // @[executor.scala 308:60]
  wire [7:0] _GEN_8653 = 8'h1 < length_3 ? _GEN_8493 : _GEN_8333; // @[executor.scala 308:60]
  wire [7:0] _GEN_8654 = 8'h1 < length_3 ? _GEN_8494 : _GEN_8334; // @[executor.scala 308:60]
  wire [7:0] _GEN_8655 = 8'h1 < length_3 ? _GEN_8495 : _GEN_8335; // @[executor.scala 308:60]
  wire [7:0] _GEN_8656 = 8'h1 < length_3 ? _GEN_8496 : _GEN_8336; // @[executor.scala 308:60]
  wire [7:0] _GEN_8657 = 8'h1 < length_3 ? _GEN_8497 : _GEN_8337; // @[executor.scala 308:60]
  wire [7:0] _GEN_8658 = 8'h1 < length_3 ? _GEN_8498 : _GEN_8338; // @[executor.scala 308:60]
  wire [7:0] _GEN_8659 = 8'h1 < length_3 ? _GEN_8499 : _GEN_8339; // @[executor.scala 308:60]
  wire [7:0] _GEN_8660 = 8'h1 < length_3 ? _GEN_8500 : _GEN_8340; // @[executor.scala 308:60]
  wire [7:0] _GEN_8661 = 8'h1 < length_3 ? _GEN_8501 : _GEN_8341; // @[executor.scala 308:60]
  wire [7:0] _GEN_8662 = 8'h1 < length_3 ? _GEN_8502 : _GEN_8342; // @[executor.scala 308:60]
  wire [7:0] _GEN_8663 = 8'h1 < length_3 ? _GEN_8503 : _GEN_8343; // @[executor.scala 308:60]
  wire [7:0] _GEN_8664 = 8'h1 < length_3 ? _GEN_8504 : _GEN_8344; // @[executor.scala 308:60]
  wire [7:0] _GEN_8665 = 8'h1 < length_3 ? _GEN_8505 : _GEN_8345; // @[executor.scala 308:60]
  wire [7:0] _GEN_8666 = 8'h1 < length_3 ? _GEN_8506 : _GEN_8346; // @[executor.scala 308:60]
  wire [7:0] _GEN_8667 = 8'h1 < length_3 ? _GEN_8507 : _GEN_8347; // @[executor.scala 308:60]
  wire [7:0] _GEN_8668 = 8'h1 < length_3 ? _GEN_8508 : _GEN_8348; // @[executor.scala 308:60]
  wire [7:0] _GEN_8669 = 8'h1 < length_3 ? _GEN_8509 : _GEN_8349; // @[executor.scala 308:60]
  wire [7:0] _GEN_8670 = 8'h1 < length_3 ? _GEN_8510 : _GEN_8350; // @[executor.scala 308:60]
  wire [7:0] _GEN_8671 = 8'h1 < length_3 ? _GEN_8511 : _GEN_8351; // @[executor.scala 308:60]
  wire [7:0] _GEN_8672 = 8'h1 < length_3 ? _GEN_8512 : _GEN_8352; // @[executor.scala 308:60]
  wire [7:0] _GEN_8673 = 8'h1 < length_3 ? _GEN_8513 : _GEN_8353; // @[executor.scala 308:60]
  wire [7:0] _GEN_8674 = 8'h1 < length_3 ? _GEN_8514 : _GEN_8354; // @[executor.scala 308:60]
  wire [7:0] _GEN_8675 = 8'h1 < length_3 ? _GEN_8515 : _GEN_8355; // @[executor.scala 308:60]
  wire [7:0] _GEN_8676 = 8'h1 < length_3 ? _GEN_8516 : _GEN_8356; // @[executor.scala 308:60]
  wire [7:0] _GEN_8677 = 8'h1 < length_3 ? _GEN_8517 : _GEN_8357; // @[executor.scala 308:60]
  wire [7:0] _GEN_8678 = 8'h1 < length_3 ? _GEN_8518 : _GEN_8358; // @[executor.scala 308:60]
  wire [7:0] _GEN_8679 = 8'h1 < length_3 ? _GEN_8519 : _GEN_8359; // @[executor.scala 308:60]
  wire [7:0] _GEN_8680 = 8'h1 < length_3 ? _GEN_8520 : _GEN_8360; // @[executor.scala 308:60]
  wire [7:0] _GEN_8681 = 8'h1 < length_3 ? _GEN_8521 : _GEN_8361; // @[executor.scala 308:60]
  wire [7:0] _GEN_8682 = 8'h1 < length_3 ? _GEN_8522 : _GEN_8362; // @[executor.scala 308:60]
  wire [7:0] _GEN_8683 = 8'h1 < length_3 ? _GEN_8523 : _GEN_8363; // @[executor.scala 308:60]
  wire [7:0] _GEN_8684 = 8'h1 < length_3 ? _GEN_8524 : _GEN_8364; // @[executor.scala 308:60]
  wire [7:0] _GEN_8685 = 8'h1 < length_3 ? _GEN_8525 : _GEN_8365; // @[executor.scala 308:60]
  wire [7:0] _GEN_8686 = 8'h1 < length_3 ? _GEN_8526 : _GEN_8366; // @[executor.scala 308:60]
  wire [7:0] _GEN_8687 = 8'h1 < length_3 ? _GEN_8527 : _GEN_8367; // @[executor.scala 308:60]
  wire [7:0] _GEN_8688 = 8'h1 < length_3 ? _GEN_8528 : _GEN_8368; // @[executor.scala 308:60]
  wire [7:0] _GEN_8689 = 8'h1 < length_3 ? _GEN_8529 : _GEN_8369; // @[executor.scala 308:60]
  wire [7:0] _GEN_8690 = 8'h1 < length_3 ? _GEN_8530 : _GEN_8370; // @[executor.scala 308:60]
  wire [7:0] _GEN_8691 = 8'h1 < length_3 ? _GEN_8531 : _GEN_8371; // @[executor.scala 308:60]
  wire [7:0] _GEN_8692 = 8'h1 < length_3 ? _GEN_8532 : _GEN_8372; // @[executor.scala 308:60]
  wire [7:0] _GEN_8693 = 8'h1 < length_3 ? _GEN_8533 : _GEN_8373; // @[executor.scala 308:60]
  wire [7:0] _GEN_8694 = 8'h1 < length_3 ? _GEN_8534 : _GEN_8374; // @[executor.scala 308:60]
  wire [7:0] _GEN_8695 = 8'h1 < length_3 ? _GEN_8535 : _GEN_8375; // @[executor.scala 308:60]
  wire [7:0] _GEN_8696 = 8'h1 < length_3 ? _GEN_8536 : _GEN_8376; // @[executor.scala 308:60]
  wire [7:0] _GEN_8697 = 8'h1 < length_3 ? _GEN_8537 : _GEN_8377; // @[executor.scala 308:60]
  wire [7:0] _GEN_8698 = 8'h1 < length_3 ? _GEN_8538 : _GEN_8378; // @[executor.scala 308:60]
  wire [7:0] _GEN_8699 = 8'h1 < length_3 ? _GEN_8539 : _GEN_8379; // @[executor.scala 308:60]
  wire [7:0] _GEN_8700 = 8'h1 < length_3 ? _GEN_8540 : _GEN_8380; // @[executor.scala 308:60]
  wire [7:0] _GEN_8701 = 8'h1 < length_3 ? _GEN_8541 : _GEN_8381; // @[executor.scala 308:60]
  wire [7:0] _GEN_8702 = 8'h1 < length_3 ? _GEN_8542 : _GEN_8382; // @[executor.scala 308:60]
  wire [7:0] _GEN_8703 = 8'h1 < length_3 ? _GEN_8543 : _GEN_8383; // @[executor.scala 308:60]
  wire [7:0] _GEN_8704 = 8'h1 < length_3 ? _GEN_8544 : _GEN_8384; // @[executor.scala 308:60]
  wire [7:0] _GEN_8705 = 8'h1 < length_3 ? _GEN_8545 : _GEN_8385; // @[executor.scala 308:60]
  wire [7:0] _GEN_8706 = 8'h1 < length_3 ? _GEN_8546 : _GEN_8386; // @[executor.scala 308:60]
  wire [7:0] _GEN_8707 = 8'h1 < length_3 ? _GEN_8547 : _GEN_8387; // @[executor.scala 308:60]
  wire [7:0] _GEN_8708 = 8'h1 < length_3 ? _GEN_8548 : _GEN_8388; // @[executor.scala 308:60]
  wire [7:0] _GEN_8709 = 8'h1 < length_3 ? _GEN_8549 : _GEN_8389; // @[executor.scala 308:60]
  wire [7:0] _GEN_8710 = 8'h1 < length_3 ? _GEN_8550 : _GEN_8390; // @[executor.scala 308:60]
  wire [7:0] _GEN_8711 = 8'h1 < length_3 ? _GEN_8551 : _GEN_8391; // @[executor.scala 308:60]
  wire [7:0] _GEN_8712 = 8'h1 < length_3 ? _GEN_8552 : _GEN_8392; // @[executor.scala 308:60]
  wire [7:0] _GEN_8713 = 8'h1 < length_3 ? _GEN_8553 : _GEN_8393; // @[executor.scala 308:60]
  wire [7:0] _GEN_8714 = 8'h1 < length_3 ? _GEN_8554 : _GEN_8394; // @[executor.scala 308:60]
  wire [7:0] _GEN_8715 = 8'h1 < length_3 ? _GEN_8555 : _GEN_8395; // @[executor.scala 308:60]
  wire [7:0] _GEN_8716 = 8'h1 < length_3 ? _GEN_8556 : _GEN_8396; // @[executor.scala 308:60]
  wire [7:0] _GEN_8717 = 8'h1 < length_3 ? _GEN_8557 : _GEN_8397; // @[executor.scala 308:60]
  wire [7:0] _GEN_8718 = 8'h1 < length_3 ? _GEN_8558 : _GEN_8398; // @[executor.scala 308:60]
  wire [7:0] _GEN_8719 = 8'h1 < length_3 ? _GEN_8559 : _GEN_8399; // @[executor.scala 308:60]
  wire [7:0] _GEN_8720 = 8'h1 < length_3 ? _GEN_8560 : _GEN_8400; // @[executor.scala 308:60]
  wire [7:0] _GEN_8721 = 8'h1 < length_3 ? _GEN_8561 : _GEN_8401; // @[executor.scala 308:60]
  wire [7:0] _GEN_8722 = 8'h1 < length_3 ? _GEN_8562 : _GEN_8402; // @[executor.scala 308:60]
  wire [7:0] _GEN_8723 = 8'h1 < length_3 ? _GEN_8563 : _GEN_8403; // @[executor.scala 308:60]
  wire [7:0] _GEN_8724 = 8'h1 < length_3 ? _GEN_8564 : _GEN_8404; // @[executor.scala 308:60]
  wire [7:0] _GEN_8725 = 8'h1 < length_3 ? _GEN_8565 : _GEN_8405; // @[executor.scala 308:60]
  wire [7:0] _GEN_8726 = 8'h1 < length_3 ? _GEN_8566 : _GEN_8406; // @[executor.scala 308:60]
  wire [7:0] _GEN_8727 = 8'h1 < length_3 ? _GEN_8567 : _GEN_8407; // @[executor.scala 308:60]
  wire [7:0] _GEN_8728 = 8'h1 < length_3 ? _GEN_8568 : _GEN_8408; // @[executor.scala 308:60]
  wire [7:0] _GEN_8729 = 8'h1 < length_3 ? _GEN_8569 : _GEN_8409; // @[executor.scala 308:60]
  wire [7:0] _GEN_8730 = 8'h1 < length_3 ? _GEN_8570 : _GEN_8410; // @[executor.scala 308:60]
  wire [7:0] _GEN_8731 = 8'h1 < length_3 ? _GEN_8571 : _GEN_8411; // @[executor.scala 308:60]
  wire [7:0] _GEN_8732 = 8'h1 < length_3 ? _GEN_8572 : _GEN_8412; // @[executor.scala 308:60]
  wire [7:0] _GEN_8733 = 8'h1 < length_3 ? _GEN_8573 : _GEN_8413; // @[executor.scala 308:60]
  wire [7:0] _GEN_8734 = 8'h1 < length_3 ? _GEN_8574 : _GEN_8414; // @[executor.scala 308:60]
  wire [7:0] _GEN_8735 = 8'h1 < length_3 ? _GEN_8575 : _GEN_8415; // @[executor.scala 308:60]
  wire [7:0] _GEN_8736 = 8'h1 < length_3 ? _GEN_8576 : _GEN_8416; // @[executor.scala 308:60]
  wire [7:0] _GEN_8737 = 8'h1 < length_3 ? _GEN_8577 : _GEN_8417; // @[executor.scala 308:60]
  wire [7:0] _GEN_8738 = 8'h1 < length_3 ? _GEN_8578 : _GEN_8418; // @[executor.scala 308:60]
  wire [7:0] _GEN_8739 = 8'h1 < length_3 ? _GEN_8579 : _GEN_8419; // @[executor.scala 308:60]
  wire [7:0] _GEN_8740 = 8'h1 < length_3 ? _GEN_8580 : _GEN_8420; // @[executor.scala 308:60]
  wire [7:0] _GEN_8741 = 8'h1 < length_3 ? _GEN_8581 : _GEN_8421; // @[executor.scala 308:60]
  wire [7:0] _GEN_8742 = 8'h1 < length_3 ? _GEN_8582 : _GEN_8422; // @[executor.scala 308:60]
  wire [7:0] _GEN_8743 = 8'h1 < length_3 ? _GEN_8583 : _GEN_8423; // @[executor.scala 308:60]
  wire [7:0] _GEN_8744 = 8'h1 < length_3 ? _GEN_8584 : _GEN_8424; // @[executor.scala 308:60]
  wire [7:0] _GEN_8745 = 8'h1 < length_3 ? _GEN_8585 : _GEN_8425; // @[executor.scala 308:60]
  wire [7:0] _GEN_8746 = 8'h1 < length_3 ? _GEN_8586 : _GEN_8426; // @[executor.scala 308:60]
  wire [7:0] _GEN_8747 = 8'h1 < length_3 ? _GEN_8587 : _GEN_8427; // @[executor.scala 308:60]
  wire [7:0] _GEN_8748 = 8'h1 < length_3 ? _GEN_8588 : _GEN_8428; // @[executor.scala 308:60]
  wire [7:0] _GEN_8749 = 8'h1 < length_3 ? _GEN_8589 : _GEN_8429; // @[executor.scala 308:60]
  wire [7:0] _GEN_8750 = 8'h1 < length_3 ? _GEN_8590 : _GEN_8430; // @[executor.scala 308:60]
  wire [7:0] _GEN_8751 = 8'h1 < length_3 ? _GEN_8591 : _GEN_8431; // @[executor.scala 308:60]
  wire [7:0] _GEN_8752 = 8'h1 < length_3 ? _GEN_8592 : _GEN_8432; // @[executor.scala 308:60]
  wire [7:0] _GEN_8753 = 8'h1 < length_3 ? _GEN_8593 : _GEN_8433; // @[executor.scala 308:60]
  wire [7:0] _GEN_8754 = 8'h1 < length_3 ? _GEN_8594 : _GEN_8434; // @[executor.scala 308:60]
  wire [7:0] _GEN_8755 = 8'h1 < length_3 ? _GEN_8595 : _GEN_8435; // @[executor.scala 308:60]
  wire [7:0] _GEN_8756 = 8'h1 < length_3 ? _GEN_8596 : _GEN_8436; // @[executor.scala 308:60]
  wire [7:0] _GEN_8757 = 8'h1 < length_3 ? _GEN_8597 : _GEN_8437; // @[executor.scala 308:60]
  wire [7:0] _GEN_8758 = 8'h1 < length_3 ? _GEN_8598 : _GEN_8438; // @[executor.scala 308:60]
  wire [7:0] _GEN_8759 = 8'h1 < length_3 ? _GEN_8599 : _GEN_8439; // @[executor.scala 308:60]
  wire [7:0] _GEN_8760 = 8'h1 < length_3 ? _GEN_8600 : _GEN_8440; // @[executor.scala 308:60]
  wire [7:0] _GEN_8761 = 8'h1 < length_3 ? _GEN_8601 : _GEN_8441; // @[executor.scala 308:60]
  wire [7:0] _GEN_8762 = 8'h1 < length_3 ? _GEN_8602 : _GEN_8442; // @[executor.scala 308:60]
  wire [7:0] _GEN_8763 = 8'h1 < length_3 ? _GEN_8603 : _GEN_8443; // @[executor.scala 308:60]
  wire [7:0] _GEN_8764 = 8'h1 < length_3 ? _GEN_8604 : _GEN_8444; // @[executor.scala 308:60]
  wire [7:0] _GEN_8765 = 8'h1 < length_3 ? _GEN_8605 : _GEN_8445; // @[executor.scala 308:60]
  wire [7:0] _GEN_8766 = 8'h1 < length_3 ? _GEN_8606 : _GEN_8446; // @[executor.scala 308:60]
  wire [7:0] _GEN_8767 = 8'h1 < length_3 ? _GEN_8607 : _GEN_8447; // @[executor.scala 308:60]
  wire [7:0] _GEN_8768 = 8'h1 < length_3 ? _GEN_8608 : _GEN_8448; // @[executor.scala 308:60]
  wire [7:0] _GEN_8769 = 8'h1 < length_3 ? _GEN_8609 : _GEN_8449; // @[executor.scala 308:60]
  wire [7:0] _GEN_8770 = 8'h1 < length_3 ? _GEN_8610 : _GEN_8450; // @[executor.scala 308:60]
  wire [7:0] _GEN_8771 = 8'h1 < length_3 ? _GEN_8611 : _GEN_8451; // @[executor.scala 308:60]
  wire [7:0] _GEN_8772 = 8'h1 < length_3 ? _GEN_8612 : _GEN_8452; // @[executor.scala 308:60]
  wire [7:0] _GEN_8773 = 8'h1 < length_3 ? _GEN_8613 : _GEN_8453; // @[executor.scala 308:60]
  wire [7:0] _GEN_8774 = 8'h1 < length_3 ? _GEN_8614 : _GEN_8454; // @[executor.scala 308:60]
  wire [7:0] _GEN_8775 = 8'h1 < length_3 ? _GEN_8615 : _GEN_8455; // @[executor.scala 308:60]
  wire [7:0] _GEN_8776 = 8'h1 < length_3 ? _GEN_8616 : _GEN_8456; // @[executor.scala 308:60]
  wire [7:0] _GEN_8777 = 8'h1 < length_3 ? _GEN_8617 : _GEN_8457; // @[executor.scala 308:60]
  wire [7:0] _GEN_8778 = 8'h1 < length_3 ? _GEN_8618 : _GEN_8458; // @[executor.scala 308:60]
  wire [7:0] _GEN_8779 = 8'h1 < length_3 ? _GEN_8619 : _GEN_8459; // @[executor.scala 308:60]
  wire [7:0] _GEN_8780 = 8'h1 < length_3 ? _GEN_8620 : _GEN_8460; // @[executor.scala 308:60]
  wire [7:0] _GEN_8781 = 8'h1 < length_3 ? _GEN_8621 : _GEN_8461; // @[executor.scala 308:60]
  wire [7:0] _GEN_8782 = 8'h1 < length_3 ? _GEN_8622 : _GEN_8462; // @[executor.scala 308:60]
  wire [7:0] _GEN_8783 = 8'h1 < length_3 ? _GEN_8623 : _GEN_8463; // @[executor.scala 308:60]
  wire [7:0] _GEN_8784 = 8'h1 < length_3 ? _GEN_8624 : _GEN_8464; // @[executor.scala 308:60]
  wire [7:0] _GEN_8785 = 8'h1 < length_3 ? _GEN_8625 : _GEN_8465; // @[executor.scala 308:60]
  wire [7:0] _GEN_8786 = 8'h1 < length_3 ? _GEN_8626 : _GEN_8466; // @[executor.scala 308:60]
  wire [7:0] _GEN_8787 = 8'h1 < length_3 ? _GEN_8627 : _GEN_8467; // @[executor.scala 308:60]
  wire [7:0] _GEN_8788 = 8'h1 < length_3 ? _GEN_8628 : _GEN_8468; // @[executor.scala 308:60]
  wire [7:0] _GEN_8789 = 8'h1 < length_3 ? _GEN_8629 : _GEN_8469; // @[executor.scala 308:60]
  wire [7:0] _GEN_8790 = 8'h1 < length_3 ? _GEN_8630 : _GEN_8470; // @[executor.scala 308:60]
  wire [7:0] _GEN_8791 = 8'h1 < length_3 ? _GEN_8631 : _GEN_8471; // @[executor.scala 308:60]
  wire [7:0] _GEN_8792 = 8'h1 < length_3 ? _GEN_8632 : _GEN_8472; // @[executor.scala 308:60]
  wire [7:0] _GEN_8793 = 8'h1 < length_3 ? _GEN_8633 : _GEN_8473; // @[executor.scala 308:60]
  wire [7:0] _GEN_8794 = 8'h1 < length_3 ? _GEN_8634 : _GEN_8474; // @[executor.scala 308:60]
  wire [7:0] _GEN_8795 = 8'h1 < length_3 ? _GEN_8635 : _GEN_8475; // @[executor.scala 308:60]
  wire [7:0] _GEN_8796 = 8'h1 < length_3 ? _GEN_8636 : _GEN_8476; // @[executor.scala 308:60]
  wire [7:0] _GEN_8797 = 8'h1 < length_3 ? _GEN_8637 : _GEN_8477; // @[executor.scala 308:60]
  wire [7:0] _GEN_8798 = 8'h1 < length_3 ? _GEN_8638 : _GEN_8478; // @[executor.scala 308:60]
  wire [7:0] _GEN_8799 = 8'h1 < length_3 ? _GEN_8639 : _GEN_8479; // @[executor.scala 308:60]
  wire [7:0] _GEN_8800 = 8'h1 < length_3 ? _GEN_8640 : _GEN_8480; // @[executor.scala 308:60]
  wire [7:0] _GEN_8801 = 8'h1 < length_3 ? _GEN_8641 : _GEN_8481; // @[executor.scala 308:60]
  wire [7:0] _GEN_8802 = 8'h1 < length_3 ? _GEN_8642 : _GEN_8482; // @[executor.scala 308:60]
  wire [7:0] _GEN_8803 = 8'h1 < length_3 ? _GEN_8643 : _GEN_8483; // @[executor.scala 308:60]
  wire [7:0] _GEN_8804 = 8'h1 < length_3 ? _GEN_8644 : _GEN_8484; // @[executor.scala 308:60]
  wire [7:0] _GEN_8805 = 8'h1 < length_3 ? _GEN_8645 : _GEN_8485; // @[executor.scala 308:60]
  wire [7:0] field_byte_26 = field_3[47:40]; // @[executor.scala 305:57]
  wire [7:0] total_offset_26 = offset_3 + 8'h2; // @[executor.scala 307:57]
  wire [7:0] _GEN_8806 = 8'h0 == total_offset_26 ? field_byte_26 : _GEN_8646; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8807 = 8'h1 == total_offset_26 ? field_byte_26 : _GEN_8647; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8808 = 8'h2 == total_offset_26 ? field_byte_26 : _GEN_8648; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8809 = 8'h3 == total_offset_26 ? field_byte_26 : _GEN_8649; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8810 = 8'h4 == total_offset_26 ? field_byte_26 : _GEN_8650; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8811 = 8'h5 == total_offset_26 ? field_byte_26 : _GEN_8651; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8812 = 8'h6 == total_offset_26 ? field_byte_26 : _GEN_8652; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8813 = 8'h7 == total_offset_26 ? field_byte_26 : _GEN_8653; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8814 = 8'h8 == total_offset_26 ? field_byte_26 : _GEN_8654; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8815 = 8'h9 == total_offset_26 ? field_byte_26 : _GEN_8655; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8816 = 8'ha == total_offset_26 ? field_byte_26 : _GEN_8656; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8817 = 8'hb == total_offset_26 ? field_byte_26 : _GEN_8657; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8818 = 8'hc == total_offset_26 ? field_byte_26 : _GEN_8658; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8819 = 8'hd == total_offset_26 ? field_byte_26 : _GEN_8659; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8820 = 8'he == total_offset_26 ? field_byte_26 : _GEN_8660; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8821 = 8'hf == total_offset_26 ? field_byte_26 : _GEN_8661; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8822 = 8'h10 == total_offset_26 ? field_byte_26 : _GEN_8662; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8823 = 8'h11 == total_offset_26 ? field_byte_26 : _GEN_8663; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8824 = 8'h12 == total_offset_26 ? field_byte_26 : _GEN_8664; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8825 = 8'h13 == total_offset_26 ? field_byte_26 : _GEN_8665; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8826 = 8'h14 == total_offset_26 ? field_byte_26 : _GEN_8666; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8827 = 8'h15 == total_offset_26 ? field_byte_26 : _GEN_8667; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8828 = 8'h16 == total_offset_26 ? field_byte_26 : _GEN_8668; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8829 = 8'h17 == total_offset_26 ? field_byte_26 : _GEN_8669; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8830 = 8'h18 == total_offset_26 ? field_byte_26 : _GEN_8670; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8831 = 8'h19 == total_offset_26 ? field_byte_26 : _GEN_8671; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8832 = 8'h1a == total_offset_26 ? field_byte_26 : _GEN_8672; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8833 = 8'h1b == total_offset_26 ? field_byte_26 : _GEN_8673; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8834 = 8'h1c == total_offset_26 ? field_byte_26 : _GEN_8674; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8835 = 8'h1d == total_offset_26 ? field_byte_26 : _GEN_8675; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8836 = 8'h1e == total_offset_26 ? field_byte_26 : _GEN_8676; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8837 = 8'h1f == total_offset_26 ? field_byte_26 : _GEN_8677; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8838 = 8'h20 == total_offset_26 ? field_byte_26 : _GEN_8678; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8839 = 8'h21 == total_offset_26 ? field_byte_26 : _GEN_8679; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8840 = 8'h22 == total_offset_26 ? field_byte_26 : _GEN_8680; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8841 = 8'h23 == total_offset_26 ? field_byte_26 : _GEN_8681; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8842 = 8'h24 == total_offset_26 ? field_byte_26 : _GEN_8682; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8843 = 8'h25 == total_offset_26 ? field_byte_26 : _GEN_8683; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8844 = 8'h26 == total_offset_26 ? field_byte_26 : _GEN_8684; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8845 = 8'h27 == total_offset_26 ? field_byte_26 : _GEN_8685; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8846 = 8'h28 == total_offset_26 ? field_byte_26 : _GEN_8686; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8847 = 8'h29 == total_offset_26 ? field_byte_26 : _GEN_8687; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8848 = 8'h2a == total_offset_26 ? field_byte_26 : _GEN_8688; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8849 = 8'h2b == total_offset_26 ? field_byte_26 : _GEN_8689; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8850 = 8'h2c == total_offset_26 ? field_byte_26 : _GEN_8690; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8851 = 8'h2d == total_offset_26 ? field_byte_26 : _GEN_8691; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8852 = 8'h2e == total_offset_26 ? field_byte_26 : _GEN_8692; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8853 = 8'h2f == total_offset_26 ? field_byte_26 : _GEN_8693; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8854 = 8'h30 == total_offset_26 ? field_byte_26 : _GEN_8694; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8855 = 8'h31 == total_offset_26 ? field_byte_26 : _GEN_8695; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8856 = 8'h32 == total_offset_26 ? field_byte_26 : _GEN_8696; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8857 = 8'h33 == total_offset_26 ? field_byte_26 : _GEN_8697; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8858 = 8'h34 == total_offset_26 ? field_byte_26 : _GEN_8698; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8859 = 8'h35 == total_offset_26 ? field_byte_26 : _GEN_8699; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8860 = 8'h36 == total_offset_26 ? field_byte_26 : _GEN_8700; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8861 = 8'h37 == total_offset_26 ? field_byte_26 : _GEN_8701; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8862 = 8'h38 == total_offset_26 ? field_byte_26 : _GEN_8702; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8863 = 8'h39 == total_offset_26 ? field_byte_26 : _GEN_8703; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8864 = 8'h3a == total_offset_26 ? field_byte_26 : _GEN_8704; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8865 = 8'h3b == total_offset_26 ? field_byte_26 : _GEN_8705; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8866 = 8'h3c == total_offset_26 ? field_byte_26 : _GEN_8706; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8867 = 8'h3d == total_offset_26 ? field_byte_26 : _GEN_8707; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8868 = 8'h3e == total_offset_26 ? field_byte_26 : _GEN_8708; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8869 = 8'h3f == total_offset_26 ? field_byte_26 : _GEN_8709; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8870 = 8'h40 == total_offset_26 ? field_byte_26 : _GEN_8710; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8871 = 8'h41 == total_offset_26 ? field_byte_26 : _GEN_8711; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8872 = 8'h42 == total_offset_26 ? field_byte_26 : _GEN_8712; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8873 = 8'h43 == total_offset_26 ? field_byte_26 : _GEN_8713; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8874 = 8'h44 == total_offset_26 ? field_byte_26 : _GEN_8714; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8875 = 8'h45 == total_offset_26 ? field_byte_26 : _GEN_8715; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8876 = 8'h46 == total_offset_26 ? field_byte_26 : _GEN_8716; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8877 = 8'h47 == total_offset_26 ? field_byte_26 : _GEN_8717; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8878 = 8'h48 == total_offset_26 ? field_byte_26 : _GEN_8718; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8879 = 8'h49 == total_offset_26 ? field_byte_26 : _GEN_8719; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8880 = 8'h4a == total_offset_26 ? field_byte_26 : _GEN_8720; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8881 = 8'h4b == total_offset_26 ? field_byte_26 : _GEN_8721; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8882 = 8'h4c == total_offset_26 ? field_byte_26 : _GEN_8722; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8883 = 8'h4d == total_offset_26 ? field_byte_26 : _GEN_8723; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8884 = 8'h4e == total_offset_26 ? field_byte_26 : _GEN_8724; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8885 = 8'h4f == total_offset_26 ? field_byte_26 : _GEN_8725; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8886 = 8'h50 == total_offset_26 ? field_byte_26 : _GEN_8726; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8887 = 8'h51 == total_offset_26 ? field_byte_26 : _GEN_8727; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8888 = 8'h52 == total_offset_26 ? field_byte_26 : _GEN_8728; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8889 = 8'h53 == total_offset_26 ? field_byte_26 : _GEN_8729; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8890 = 8'h54 == total_offset_26 ? field_byte_26 : _GEN_8730; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8891 = 8'h55 == total_offset_26 ? field_byte_26 : _GEN_8731; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8892 = 8'h56 == total_offset_26 ? field_byte_26 : _GEN_8732; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8893 = 8'h57 == total_offset_26 ? field_byte_26 : _GEN_8733; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8894 = 8'h58 == total_offset_26 ? field_byte_26 : _GEN_8734; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8895 = 8'h59 == total_offset_26 ? field_byte_26 : _GEN_8735; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8896 = 8'h5a == total_offset_26 ? field_byte_26 : _GEN_8736; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8897 = 8'h5b == total_offset_26 ? field_byte_26 : _GEN_8737; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8898 = 8'h5c == total_offset_26 ? field_byte_26 : _GEN_8738; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8899 = 8'h5d == total_offset_26 ? field_byte_26 : _GEN_8739; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8900 = 8'h5e == total_offset_26 ? field_byte_26 : _GEN_8740; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8901 = 8'h5f == total_offset_26 ? field_byte_26 : _GEN_8741; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8902 = 8'h60 == total_offset_26 ? field_byte_26 : _GEN_8742; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8903 = 8'h61 == total_offset_26 ? field_byte_26 : _GEN_8743; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8904 = 8'h62 == total_offset_26 ? field_byte_26 : _GEN_8744; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8905 = 8'h63 == total_offset_26 ? field_byte_26 : _GEN_8745; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8906 = 8'h64 == total_offset_26 ? field_byte_26 : _GEN_8746; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8907 = 8'h65 == total_offset_26 ? field_byte_26 : _GEN_8747; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8908 = 8'h66 == total_offset_26 ? field_byte_26 : _GEN_8748; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8909 = 8'h67 == total_offset_26 ? field_byte_26 : _GEN_8749; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8910 = 8'h68 == total_offset_26 ? field_byte_26 : _GEN_8750; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8911 = 8'h69 == total_offset_26 ? field_byte_26 : _GEN_8751; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8912 = 8'h6a == total_offset_26 ? field_byte_26 : _GEN_8752; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8913 = 8'h6b == total_offset_26 ? field_byte_26 : _GEN_8753; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8914 = 8'h6c == total_offset_26 ? field_byte_26 : _GEN_8754; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8915 = 8'h6d == total_offset_26 ? field_byte_26 : _GEN_8755; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8916 = 8'h6e == total_offset_26 ? field_byte_26 : _GEN_8756; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8917 = 8'h6f == total_offset_26 ? field_byte_26 : _GEN_8757; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8918 = 8'h70 == total_offset_26 ? field_byte_26 : _GEN_8758; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8919 = 8'h71 == total_offset_26 ? field_byte_26 : _GEN_8759; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8920 = 8'h72 == total_offset_26 ? field_byte_26 : _GEN_8760; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8921 = 8'h73 == total_offset_26 ? field_byte_26 : _GEN_8761; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8922 = 8'h74 == total_offset_26 ? field_byte_26 : _GEN_8762; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8923 = 8'h75 == total_offset_26 ? field_byte_26 : _GEN_8763; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8924 = 8'h76 == total_offset_26 ? field_byte_26 : _GEN_8764; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8925 = 8'h77 == total_offset_26 ? field_byte_26 : _GEN_8765; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8926 = 8'h78 == total_offset_26 ? field_byte_26 : _GEN_8766; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8927 = 8'h79 == total_offset_26 ? field_byte_26 : _GEN_8767; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8928 = 8'h7a == total_offset_26 ? field_byte_26 : _GEN_8768; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8929 = 8'h7b == total_offset_26 ? field_byte_26 : _GEN_8769; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8930 = 8'h7c == total_offset_26 ? field_byte_26 : _GEN_8770; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8931 = 8'h7d == total_offset_26 ? field_byte_26 : _GEN_8771; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8932 = 8'h7e == total_offset_26 ? field_byte_26 : _GEN_8772; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8933 = 8'h7f == total_offset_26 ? field_byte_26 : _GEN_8773; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8934 = 8'h80 == total_offset_26 ? field_byte_26 : _GEN_8774; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8935 = 8'h81 == total_offset_26 ? field_byte_26 : _GEN_8775; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8936 = 8'h82 == total_offset_26 ? field_byte_26 : _GEN_8776; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8937 = 8'h83 == total_offset_26 ? field_byte_26 : _GEN_8777; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8938 = 8'h84 == total_offset_26 ? field_byte_26 : _GEN_8778; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8939 = 8'h85 == total_offset_26 ? field_byte_26 : _GEN_8779; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8940 = 8'h86 == total_offset_26 ? field_byte_26 : _GEN_8780; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8941 = 8'h87 == total_offset_26 ? field_byte_26 : _GEN_8781; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8942 = 8'h88 == total_offset_26 ? field_byte_26 : _GEN_8782; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8943 = 8'h89 == total_offset_26 ? field_byte_26 : _GEN_8783; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8944 = 8'h8a == total_offset_26 ? field_byte_26 : _GEN_8784; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8945 = 8'h8b == total_offset_26 ? field_byte_26 : _GEN_8785; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8946 = 8'h8c == total_offset_26 ? field_byte_26 : _GEN_8786; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8947 = 8'h8d == total_offset_26 ? field_byte_26 : _GEN_8787; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8948 = 8'h8e == total_offset_26 ? field_byte_26 : _GEN_8788; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8949 = 8'h8f == total_offset_26 ? field_byte_26 : _GEN_8789; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8950 = 8'h90 == total_offset_26 ? field_byte_26 : _GEN_8790; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8951 = 8'h91 == total_offset_26 ? field_byte_26 : _GEN_8791; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8952 = 8'h92 == total_offset_26 ? field_byte_26 : _GEN_8792; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8953 = 8'h93 == total_offset_26 ? field_byte_26 : _GEN_8793; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8954 = 8'h94 == total_offset_26 ? field_byte_26 : _GEN_8794; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8955 = 8'h95 == total_offset_26 ? field_byte_26 : _GEN_8795; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8956 = 8'h96 == total_offset_26 ? field_byte_26 : _GEN_8796; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8957 = 8'h97 == total_offset_26 ? field_byte_26 : _GEN_8797; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8958 = 8'h98 == total_offset_26 ? field_byte_26 : _GEN_8798; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8959 = 8'h99 == total_offset_26 ? field_byte_26 : _GEN_8799; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8960 = 8'h9a == total_offset_26 ? field_byte_26 : _GEN_8800; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8961 = 8'h9b == total_offset_26 ? field_byte_26 : _GEN_8801; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8962 = 8'h9c == total_offset_26 ? field_byte_26 : _GEN_8802; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8963 = 8'h9d == total_offset_26 ? field_byte_26 : _GEN_8803; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8964 = 8'h9e == total_offset_26 ? field_byte_26 : _GEN_8804; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8965 = 8'h9f == total_offset_26 ? field_byte_26 : _GEN_8805; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_8966 = 8'h2 < length_3 ? _GEN_8806 : _GEN_8646; // @[executor.scala 308:60]
  wire [7:0] _GEN_8967 = 8'h2 < length_3 ? _GEN_8807 : _GEN_8647; // @[executor.scala 308:60]
  wire [7:0] _GEN_8968 = 8'h2 < length_3 ? _GEN_8808 : _GEN_8648; // @[executor.scala 308:60]
  wire [7:0] _GEN_8969 = 8'h2 < length_3 ? _GEN_8809 : _GEN_8649; // @[executor.scala 308:60]
  wire [7:0] _GEN_8970 = 8'h2 < length_3 ? _GEN_8810 : _GEN_8650; // @[executor.scala 308:60]
  wire [7:0] _GEN_8971 = 8'h2 < length_3 ? _GEN_8811 : _GEN_8651; // @[executor.scala 308:60]
  wire [7:0] _GEN_8972 = 8'h2 < length_3 ? _GEN_8812 : _GEN_8652; // @[executor.scala 308:60]
  wire [7:0] _GEN_8973 = 8'h2 < length_3 ? _GEN_8813 : _GEN_8653; // @[executor.scala 308:60]
  wire [7:0] _GEN_8974 = 8'h2 < length_3 ? _GEN_8814 : _GEN_8654; // @[executor.scala 308:60]
  wire [7:0] _GEN_8975 = 8'h2 < length_3 ? _GEN_8815 : _GEN_8655; // @[executor.scala 308:60]
  wire [7:0] _GEN_8976 = 8'h2 < length_3 ? _GEN_8816 : _GEN_8656; // @[executor.scala 308:60]
  wire [7:0] _GEN_8977 = 8'h2 < length_3 ? _GEN_8817 : _GEN_8657; // @[executor.scala 308:60]
  wire [7:0] _GEN_8978 = 8'h2 < length_3 ? _GEN_8818 : _GEN_8658; // @[executor.scala 308:60]
  wire [7:0] _GEN_8979 = 8'h2 < length_3 ? _GEN_8819 : _GEN_8659; // @[executor.scala 308:60]
  wire [7:0] _GEN_8980 = 8'h2 < length_3 ? _GEN_8820 : _GEN_8660; // @[executor.scala 308:60]
  wire [7:0] _GEN_8981 = 8'h2 < length_3 ? _GEN_8821 : _GEN_8661; // @[executor.scala 308:60]
  wire [7:0] _GEN_8982 = 8'h2 < length_3 ? _GEN_8822 : _GEN_8662; // @[executor.scala 308:60]
  wire [7:0] _GEN_8983 = 8'h2 < length_3 ? _GEN_8823 : _GEN_8663; // @[executor.scala 308:60]
  wire [7:0] _GEN_8984 = 8'h2 < length_3 ? _GEN_8824 : _GEN_8664; // @[executor.scala 308:60]
  wire [7:0] _GEN_8985 = 8'h2 < length_3 ? _GEN_8825 : _GEN_8665; // @[executor.scala 308:60]
  wire [7:0] _GEN_8986 = 8'h2 < length_3 ? _GEN_8826 : _GEN_8666; // @[executor.scala 308:60]
  wire [7:0] _GEN_8987 = 8'h2 < length_3 ? _GEN_8827 : _GEN_8667; // @[executor.scala 308:60]
  wire [7:0] _GEN_8988 = 8'h2 < length_3 ? _GEN_8828 : _GEN_8668; // @[executor.scala 308:60]
  wire [7:0] _GEN_8989 = 8'h2 < length_3 ? _GEN_8829 : _GEN_8669; // @[executor.scala 308:60]
  wire [7:0] _GEN_8990 = 8'h2 < length_3 ? _GEN_8830 : _GEN_8670; // @[executor.scala 308:60]
  wire [7:0] _GEN_8991 = 8'h2 < length_3 ? _GEN_8831 : _GEN_8671; // @[executor.scala 308:60]
  wire [7:0] _GEN_8992 = 8'h2 < length_3 ? _GEN_8832 : _GEN_8672; // @[executor.scala 308:60]
  wire [7:0] _GEN_8993 = 8'h2 < length_3 ? _GEN_8833 : _GEN_8673; // @[executor.scala 308:60]
  wire [7:0] _GEN_8994 = 8'h2 < length_3 ? _GEN_8834 : _GEN_8674; // @[executor.scala 308:60]
  wire [7:0] _GEN_8995 = 8'h2 < length_3 ? _GEN_8835 : _GEN_8675; // @[executor.scala 308:60]
  wire [7:0] _GEN_8996 = 8'h2 < length_3 ? _GEN_8836 : _GEN_8676; // @[executor.scala 308:60]
  wire [7:0] _GEN_8997 = 8'h2 < length_3 ? _GEN_8837 : _GEN_8677; // @[executor.scala 308:60]
  wire [7:0] _GEN_8998 = 8'h2 < length_3 ? _GEN_8838 : _GEN_8678; // @[executor.scala 308:60]
  wire [7:0] _GEN_8999 = 8'h2 < length_3 ? _GEN_8839 : _GEN_8679; // @[executor.scala 308:60]
  wire [7:0] _GEN_9000 = 8'h2 < length_3 ? _GEN_8840 : _GEN_8680; // @[executor.scala 308:60]
  wire [7:0] _GEN_9001 = 8'h2 < length_3 ? _GEN_8841 : _GEN_8681; // @[executor.scala 308:60]
  wire [7:0] _GEN_9002 = 8'h2 < length_3 ? _GEN_8842 : _GEN_8682; // @[executor.scala 308:60]
  wire [7:0] _GEN_9003 = 8'h2 < length_3 ? _GEN_8843 : _GEN_8683; // @[executor.scala 308:60]
  wire [7:0] _GEN_9004 = 8'h2 < length_3 ? _GEN_8844 : _GEN_8684; // @[executor.scala 308:60]
  wire [7:0] _GEN_9005 = 8'h2 < length_3 ? _GEN_8845 : _GEN_8685; // @[executor.scala 308:60]
  wire [7:0] _GEN_9006 = 8'h2 < length_3 ? _GEN_8846 : _GEN_8686; // @[executor.scala 308:60]
  wire [7:0] _GEN_9007 = 8'h2 < length_3 ? _GEN_8847 : _GEN_8687; // @[executor.scala 308:60]
  wire [7:0] _GEN_9008 = 8'h2 < length_3 ? _GEN_8848 : _GEN_8688; // @[executor.scala 308:60]
  wire [7:0] _GEN_9009 = 8'h2 < length_3 ? _GEN_8849 : _GEN_8689; // @[executor.scala 308:60]
  wire [7:0] _GEN_9010 = 8'h2 < length_3 ? _GEN_8850 : _GEN_8690; // @[executor.scala 308:60]
  wire [7:0] _GEN_9011 = 8'h2 < length_3 ? _GEN_8851 : _GEN_8691; // @[executor.scala 308:60]
  wire [7:0] _GEN_9012 = 8'h2 < length_3 ? _GEN_8852 : _GEN_8692; // @[executor.scala 308:60]
  wire [7:0] _GEN_9013 = 8'h2 < length_3 ? _GEN_8853 : _GEN_8693; // @[executor.scala 308:60]
  wire [7:0] _GEN_9014 = 8'h2 < length_3 ? _GEN_8854 : _GEN_8694; // @[executor.scala 308:60]
  wire [7:0] _GEN_9015 = 8'h2 < length_3 ? _GEN_8855 : _GEN_8695; // @[executor.scala 308:60]
  wire [7:0] _GEN_9016 = 8'h2 < length_3 ? _GEN_8856 : _GEN_8696; // @[executor.scala 308:60]
  wire [7:0] _GEN_9017 = 8'h2 < length_3 ? _GEN_8857 : _GEN_8697; // @[executor.scala 308:60]
  wire [7:0] _GEN_9018 = 8'h2 < length_3 ? _GEN_8858 : _GEN_8698; // @[executor.scala 308:60]
  wire [7:0] _GEN_9019 = 8'h2 < length_3 ? _GEN_8859 : _GEN_8699; // @[executor.scala 308:60]
  wire [7:0] _GEN_9020 = 8'h2 < length_3 ? _GEN_8860 : _GEN_8700; // @[executor.scala 308:60]
  wire [7:0] _GEN_9021 = 8'h2 < length_3 ? _GEN_8861 : _GEN_8701; // @[executor.scala 308:60]
  wire [7:0] _GEN_9022 = 8'h2 < length_3 ? _GEN_8862 : _GEN_8702; // @[executor.scala 308:60]
  wire [7:0] _GEN_9023 = 8'h2 < length_3 ? _GEN_8863 : _GEN_8703; // @[executor.scala 308:60]
  wire [7:0] _GEN_9024 = 8'h2 < length_3 ? _GEN_8864 : _GEN_8704; // @[executor.scala 308:60]
  wire [7:0] _GEN_9025 = 8'h2 < length_3 ? _GEN_8865 : _GEN_8705; // @[executor.scala 308:60]
  wire [7:0] _GEN_9026 = 8'h2 < length_3 ? _GEN_8866 : _GEN_8706; // @[executor.scala 308:60]
  wire [7:0] _GEN_9027 = 8'h2 < length_3 ? _GEN_8867 : _GEN_8707; // @[executor.scala 308:60]
  wire [7:0] _GEN_9028 = 8'h2 < length_3 ? _GEN_8868 : _GEN_8708; // @[executor.scala 308:60]
  wire [7:0] _GEN_9029 = 8'h2 < length_3 ? _GEN_8869 : _GEN_8709; // @[executor.scala 308:60]
  wire [7:0] _GEN_9030 = 8'h2 < length_3 ? _GEN_8870 : _GEN_8710; // @[executor.scala 308:60]
  wire [7:0] _GEN_9031 = 8'h2 < length_3 ? _GEN_8871 : _GEN_8711; // @[executor.scala 308:60]
  wire [7:0] _GEN_9032 = 8'h2 < length_3 ? _GEN_8872 : _GEN_8712; // @[executor.scala 308:60]
  wire [7:0] _GEN_9033 = 8'h2 < length_3 ? _GEN_8873 : _GEN_8713; // @[executor.scala 308:60]
  wire [7:0] _GEN_9034 = 8'h2 < length_3 ? _GEN_8874 : _GEN_8714; // @[executor.scala 308:60]
  wire [7:0] _GEN_9035 = 8'h2 < length_3 ? _GEN_8875 : _GEN_8715; // @[executor.scala 308:60]
  wire [7:0] _GEN_9036 = 8'h2 < length_3 ? _GEN_8876 : _GEN_8716; // @[executor.scala 308:60]
  wire [7:0] _GEN_9037 = 8'h2 < length_3 ? _GEN_8877 : _GEN_8717; // @[executor.scala 308:60]
  wire [7:0] _GEN_9038 = 8'h2 < length_3 ? _GEN_8878 : _GEN_8718; // @[executor.scala 308:60]
  wire [7:0] _GEN_9039 = 8'h2 < length_3 ? _GEN_8879 : _GEN_8719; // @[executor.scala 308:60]
  wire [7:0] _GEN_9040 = 8'h2 < length_3 ? _GEN_8880 : _GEN_8720; // @[executor.scala 308:60]
  wire [7:0] _GEN_9041 = 8'h2 < length_3 ? _GEN_8881 : _GEN_8721; // @[executor.scala 308:60]
  wire [7:0] _GEN_9042 = 8'h2 < length_3 ? _GEN_8882 : _GEN_8722; // @[executor.scala 308:60]
  wire [7:0] _GEN_9043 = 8'h2 < length_3 ? _GEN_8883 : _GEN_8723; // @[executor.scala 308:60]
  wire [7:0] _GEN_9044 = 8'h2 < length_3 ? _GEN_8884 : _GEN_8724; // @[executor.scala 308:60]
  wire [7:0] _GEN_9045 = 8'h2 < length_3 ? _GEN_8885 : _GEN_8725; // @[executor.scala 308:60]
  wire [7:0] _GEN_9046 = 8'h2 < length_3 ? _GEN_8886 : _GEN_8726; // @[executor.scala 308:60]
  wire [7:0] _GEN_9047 = 8'h2 < length_3 ? _GEN_8887 : _GEN_8727; // @[executor.scala 308:60]
  wire [7:0] _GEN_9048 = 8'h2 < length_3 ? _GEN_8888 : _GEN_8728; // @[executor.scala 308:60]
  wire [7:0] _GEN_9049 = 8'h2 < length_3 ? _GEN_8889 : _GEN_8729; // @[executor.scala 308:60]
  wire [7:0] _GEN_9050 = 8'h2 < length_3 ? _GEN_8890 : _GEN_8730; // @[executor.scala 308:60]
  wire [7:0] _GEN_9051 = 8'h2 < length_3 ? _GEN_8891 : _GEN_8731; // @[executor.scala 308:60]
  wire [7:0] _GEN_9052 = 8'h2 < length_3 ? _GEN_8892 : _GEN_8732; // @[executor.scala 308:60]
  wire [7:0] _GEN_9053 = 8'h2 < length_3 ? _GEN_8893 : _GEN_8733; // @[executor.scala 308:60]
  wire [7:0] _GEN_9054 = 8'h2 < length_3 ? _GEN_8894 : _GEN_8734; // @[executor.scala 308:60]
  wire [7:0] _GEN_9055 = 8'h2 < length_3 ? _GEN_8895 : _GEN_8735; // @[executor.scala 308:60]
  wire [7:0] _GEN_9056 = 8'h2 < length_3 ? _GEN_8896 : _GEN_8736; // @[executor.scala 308:60]
  wire [7:0] _GEN_9057 = 8'h2 < length_3 ? _GEN_8897 : _GEN_8737; // @[executor.scala 308:60]
  wire [7:0] _GEN_9058 = 8'h2 < length_3 ? _GEN_8898 : _GEN_8738; // @[executor.scala 308:60]
  wire [7:0] _GEN_9059 = 8'h2 < length_3 ? _GEN_8899 : _GEN_8739; // @[executor.scala 308:60]
  wire [7:0] _GEN_9060 = 8'h2 < length_3 ? _GEN_8900 : _GEN_8740; // @[executor.scala 308:60]
  wire [7:0] _GEN_9061 = 8'h2 < length_3 ? _GEN_8901 : _GEN_8741; // @[executor.scala 308:60]
  wire [7:0] _GEN_9062 = 8'h2 < length_3 ? _GEN_8902 : _GEN_8742; // @[executor.scala 308:60]
  wire [7:0] _GEN_9063 = 8'h2 < length_3 ? _GEN_8903 : _GEN_8743; // @[executor.scala 308:60]
  wire [7:0] _GEN_9064 = 8'h2 < length_3 ? _GEN_8904 : _GEN_8744; // @[executor.scala 308:60]
  wire [7:0] _GEN_9065 = 8'h2 < length_3 ? _GEN_8905 : _GEN_8745; // @[executor.scala 308:60]
  wire [7:0] _GEN_9066 = 8'h2 < length_3 ? _GEN_8906 : _GEN_8746; // @[executor.scala 308:60]
  wire [7:0] _GEN_9067 = 8'h2 < length_3 ? _GEN_8907 : _GEN_8747; // @[executor.scala 308:60]
  wire [7:0] _GEN_9068 = 8'h2 < length_3 ? _GEN_8908 : _GEN_8748; // @[executor.scala 308:60]
  wire [7:0] _GEN_9069 = 8'h2 < length_3 ? _GEN_8909 : _GEN_8749; // @[executor.scala 308:60]
  wire [7:0] _GEN_9070 = 8'h2 < length_3 ? _GEN_8910 : _GEN_8750; // @[executor.scala 308:60]
  wire [7:0] _GEN_9071 = 8'h2 < length_3 ? _GEN_8911 : _GEN_8751; // @[executor.scala 308:60]
  wire [7:0] _GEN_9072 = 8'h2 < length_3 ? _GEN_8912 : _GEN_8752; // @[executor.scala 308:60]
  wire [7:0] _GEN_9073 = 8'h2 < length_3 ? _GEN_8913 : _GEN_8753; // @[executor.scala 308:60]
  wire [7:0] _GEN_9074 = 8'h2 < length_3 ? _GEN_8914 : _GEN_8754; // @[executor.scala 308:60]
  wire [7:0] _GEN_9075 = 8'h2 < length_3 ? _GEN_8915 : _GEN_8755; // @[executor.scala 308:60]
  wire [7:0] _GEN_9076 = 8'h2 < length_3 ? _GEN_8916 : _GEN_8756; // @[executor.scala 308:60]
  wire [7:0] _GEN_9077 = 8'h2 < length_3 ? _GEN_8917 : _GEN_8757; // @[executor.scala 308:60]
  wire [7:0] _GEN_9078 = 8'h2 < length_3 ? _GEN_8918 : _GEN_8758; // @[executor.scala 308:60]
  wire [7:0] _GEN_9079 = 8'h2 < length_3 ? _GEN_8919 : _GEN_8759; // @[executor.scala 308:60]
  wire [7:0] _GEN_9080 = 8'h2 < length_3 ? _GEN_8920 : _GEN_8760; // @[executor.scala 308:60]
  wire [7:0] _GEN_9081 = 8'h2 < length_3 ? _GEN_8921 : _GEN_8761; // @[executor.scala 308:60]
  wire [7:0] _GEN_9082 = 8'h2 < length_3 ? _GEN_8922 : _GEN_8762; // @[executor.scala 308:60]
  wire [7:0] _GEN_9083 = 8'h2 < length_3 ? _GEN_8923 : _GEN_8763; // @[executor.scala 308:60]
  wire [7:0] _GEN_9084 = 8'h2 < length_3 ? _GEN_8924 : _GEN_8764; // @[executor.scala 308:60]
  wire [7:0] _GEN_9085 = 8'h2 < length_3 ? _GEN_8925 : _GEN_8765; // @[executor.scala 308:60]
  wire [7:0] _GEN_9086 = 8'h2 < length_3 ? _GEN_8926 : _GEN_8766; // @[executor.scala 308:60]
  wire [7:0] _GEN_9087 = 8'h2 < length_3 ? _GEN_8927 : _GEN_8767; // @[executor.scala 308:60]
  wire [7:0] _GEN_9088 = 8'h2 < length_3 ? _GEN_8928 : _GEN_8768; // @[executor.scala 308:60]
  wire [7:0] _GEN_9089 = 8'h2 < length_3 ? _GEN_8929 : _GEN_8769; // @[executor.scala 308:60]
  wire [7:0] _GEN_9090 = 8'h2 < length_3 ? _GEN_8930 : _GEN_8770; // @[executor.scala 308:60]
  wire [7:0] _GEN_9091 = 8'h2 < length_3 ? _GEN_8931 : _GEN_8771; // @[executor.scala 308:60]
  wire [7:0] _GEN_9092 = 8'h2 < length_3 ? _GEN_8932 : _GEN_8772; // @[executor.scala 308:60]
  wire [7:0] _GEN_9093 = 8'h2 < length_3 ? _GEN_8933 : _GEN_8773; // @[executor.scala 308:60]
  wire [7:0] _GEN_9094 = 8'h2 < length_3 ? _GEN_8934 : _GEN_8774; // @[executor.scala 308:60]
  wire [7:0] _GEN_9095 = 8'h2 < length_3 ? _GEN_8935 : _GEN_8775; // @[executor.scala 308:60]
  wire [7:0] _GEN_9096 = 8'h2 < length_3 ? _GEN_8936 : _GEN_8776; // @[executor.scala 308:60]
  wire [7:0] _GEN_9097 = 8'h2 < length_3 ? _GEN_8937 : _GEN_8777; // @[executor.scala 308:60]
  wire [7:0] _GEN_9098 = 8'h2 < length_3 ? _GEN_8938 : _GEN_8778; // @[executor.scala 308:60]
  wire [7:0] _GEN_9099 = 8'h2 < length_3 ? _GEN_8939 : _GEN_8779; // @[executor.scala 308:60]
  wire [7:0] _GEN_9100 = 8'h2 < length_3 ? _GEN_8940 : _GEN_8780; // @[executor.scala 308:60]
  wire [7:0] _GEN_9101 = 8'h2 < length_3 ? _GEN_8941 : _GEN_8781; // @[executor.scala 308:60]
  wire [7:0] _GEN_9102 = 8'h2 < length_3 ? _GEN_8942 : _GEN_8782; // @[executor.scala 308:60]
  wire [7:0] _GEN_9103 = 8'h2 < length_3 ? _GEN_8943 : _GEN_8783; // @[executor.scala 308:60]
  wire [7:0] _GEN_9104 = 8'h2 < length_3 ? _GEN_8944 : _GEN_8784; // @[executor.scala 308:60]
  wire [7:0] _GEN_9105 = 8'h2 < length_3 ? _GEN_8945 : _GEN_8785; // @[executor.scala 308:60]
  wire [7:0] _GEN_9106 = 8'h2 < length_3 ? _GEN_8946 : _GEN_8786; // @[executor.scala 308:60]
  wire [7:0] _GEN_9107 = 8'h2 < length_3 ? _GEN_8947 : _GEN_8787; // @[executor.scala 308:60]
  wire [7:0] _GEN_9108 = 8'h2 < length_3 ? _GEN_8948 : _GEN_8788; // @[executor.scala 308:60]
  wire [7:0] _GEN_9109 = 8'h2 < length_3 ? _GEN_8949 : _GEN_8789; // @[executor.scala 308:60]
  wire [7:0] _GEN_9110 = 8'h2 < length_3 ? _GEN_8950 : _GEN_8790; // @[executor.scala 308:60]
  wire [7:0] _GEN_9111 = 8'h2 < length_3 ? _GEN_8951 : _GEN_8791; // @[executor.scala 308:60]
  wire [7:0] _GEN_9112 = 8'h2 < length_3 ? _GEN_8952 : _GEN_8792; // @[executor.scala 308:60]
  wire [7:0] _GEN_9113 = 8'h2 < length_3 ? _GEN_8953 : _GEN_8793; // @[executor.scala 308:60]
  wire [7:0] _GEN_9114 = 8'h2 < length_3 ? _GEN_8954 : _GEN_8794; // @[executor.scala 308:60]
  wire [7:0] _GEN_9115 = 8'h2 < length_3 ? _GEN_8955 : _GEN_8795; // @[executor.scala 308:60]
  wire [7:0] _GEN_9116 = 8'h2 < length_3 ? _GEN_8956 : _GEN_8796; // @[executor.scala 308:60]
  wire [7:0] _GEN_9117 = 8'h2 < length_3 ? _GEN_8957 : _GEN_8797; // @[executor.scala 308:60]
  wire [7:0] _GEN_9118 = 8'h2 < length_3 ? _GEN_8958 : _GEN_8798; // @[executor.scala 308:60]
  wire [7:0] _GEN_9119 = 8'h2 < length_3 ? _GEN_8959 : _GEN_8799; // @[executor.scala 308:60]
  wire [7:0] _GEN_9120 = 8'h2 < length_3 ? _GEN_8960 : _GEN_8800; // @[executor.scala 308:60]
  wire [7:0] _GEN_9121 = 8'h2 < length_3 ? _GEN_8961 : _GEN_8801; // @[executor.scala 308:60]
  wire [7:0] _GEN_9122 = 8'h2 < length_3 ? _GEN_8962 : _GEN_8802; // @[executor.scala 308:60]
  wire [7:0] _GEN_9123 = 8'h2 < length_3 ? _GEN_8963 : _GEN_8803; // @[executor.scala 308:60]
  wire [7:0] _GEN_9124 = 8'h2 < length_3 ? _GEN_8964 : _GEN_8804; // @[executor.scala 308:60]
  wire [7:0] _GEN_9125 = 8'h2 < length_3 ? _GEN_8965 : _GEN_8805; // @[executor.scala 308:60]
  wire [7:0] field_byte_27 = field_3[39:32]; // @[executor.scala 305:57]
  wire [7:0] total_offset_27 = offset_3 + 8'h3; // @[executor.scala 307:57]
  wire [7:0] _GEN_9126 = 8'h0 == total_offset_27 ? field_byte_27 : _GEN_8966; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9127 = 8'h1 == total_offset_27 ? field_byte_27 : _GEN_8967; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9128 = 8'h2 == total_offset_27 ? field_byte_27 : _GEN_8968; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9129 = 8'h3 == total_offset_27 ? field_byte_27 : _GEN_8969; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9130 = 8'h4 == total_offset_27 ? field_byte_27 : _GEN_8970; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9131 = 8'h5 == total_offset_27 ? field_byte_27 : _GEN_8971; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9132 = 8'h6 == total_offset_27 ? field_byte_27 : _GEN_8972; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9133 = 8'h7 == total_offset_27 ? field_byte_27 : _GEN_8973; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9134 = 8'h8 == total_offset_27 ? field_byte_27 : _GEN_8974; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9135 = 8'h9 == total_offset_27 ? field_byte_27 : _GEN_8975; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9136 = 8'ha == total_offset_27 ? field_byte_27 : _GEN_8976; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9137 = 8'hb == total_offset_27 ? field_byte_27 : _GEN_8977; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9138 = 8'hc == total_offset_27 ? field_byte_27 : _GEN_8978; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9139 = 8'hd == total_offset_27 ? field_byte_27 : _GEN_8979; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9140 = 8'he == total_offset_27 ? field_byte_27 : _GEN_8980; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9141 = 8'hf == total_offset_27 ? field_byte_27 : _GEN_8981; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9142 = 8'h10 == total_offset_27 ? field_byte_27 : _GEN_8982; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9143 = 8'h11 == total_offset_27 ? field_byte_27 : _GEN_8983; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9144 = 8'h12 == total_offset_27 ? field_byte_27 : _GEN_8984; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9145 = 8'h13 == total_offset_27 ? field_byte_27 : _GEN_8985; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9146 = 8'h14 == total_offset_27 ? field_byte_27 : _GEN_8986; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9147 = 8'h15 == total_offset_27 ? field_byte_27 : _GEN_8987; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9148 = 8'h16 == total_offset_27 ? field_byte_27 : _GEN_8988; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9149 = 8'h17 == total_offset_27 ? field_byte_27 : _GEN_8989; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9150 = 8'h18 == total_offset_27 ? field_byte_27 : _GEN_8990; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9151 = 8'h19 == total_offset_27 ? field_byte_27 : _GEN_8991; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9152 = 8'h1a == total_offset_27 ? field_byte_27 : _GEN_8992; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9153 = 8'h1b == total_offset_27 ? field_byte_27 : _GEN_8993; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9154 = 8'h1c == total_offset_27 ? field_byte_27 : _GEN_8994; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9155 = 8'h1d == total_offset_27 ? field_byte_27 : _GEN_8995; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9156 = 8'h1e == total_offset_27 ? field_byte_27 : _GEN_8996; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9157 = 8'h1f == total_offset_27 ? field_byte_27 : _GEN_8997; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9158 = 8'h20 == total_offset_27 ? field_byte_27 : _GEN_8998; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9159 = 8'h21 == total_offset_27 ? field_byte_27 : _GEN_8999; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9160 = 8'h22 == total_offset_27 ? field_byte_27 : _GEN_9000; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9161 = 8'h23 == total_offset_27 ? field_byte_27 : _GEN_9001; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9162 = 8'h24 == total_offset_27 ? field_byte_27 : _GEN_9002; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9163 = 8'h25 == total_offset_27 ? field_byte_27 : _GEN_9003; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9164 = 8'h26 == total_offset_27 ? field_byte_27 : _GEN_9004; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9165 = 8'h27 == total_offset_27 ? field_byte_27 : _GEN_9005; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9166 = 8'h28 == total_offset_27 ? field_byte_27 : _GEN_9006; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9167 = 8'h29 == total_offset_27 ? field_byte_27 : _GEN_9007; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9168 = 8'h2a == total_offset_27 ? field_byte_27 : _GEN_9008; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9169 = 8'h2b == total_offset_27 ? field_byte_27 : _GEN_9009; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9170 = 8'h2c == total_offset_27 ? field_byte_27 : _GEN_9010; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9171 = 8'h2d == total_offset_27 ? field_byte_27 : _GEN_9011; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9172 = 8'h2e == total_offset_27 ? field_byte_27 : _GEN_9012; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9173 = 8'h2f == total_offset_27 ? field_byte_27 : _GEN_9013; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9174 = 8'h30 == total_offset_27 ? field_byte_27 : _GEN_9014; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9175 = 8'h31 == total_offset_27 ? field_byte_27 : _GEN_9015; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9176 = 8'h32 == total_offset_27 ? field_byte_27 : _GEN_9016; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9177 = 8'h33 == total_offset_27 ? field_byte_27 : _GEN_9017; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9178 = 8'h34 == total_offset_27 ? field_byte_27 : _GEN_9018; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9179 = 8'h35 == total_offset_27 ? field_byte_27 : _GEN_9019; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9180 = 8'h36 == total_offset_27 ? field_byte_27 : _GEN_9020; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9181 = 8'h37 == total_offset_27 ? field_byte_27 : _GEN_9021; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9182 = 8'h38 == total_offset_27 ? field_byte_27 : _GEN_9022; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9183 = 8'h39 == total_offset_27 ? field_byte_27 : _GEN_9023; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9184 = 8'h3a == total_offset_27 ? field_byte_27 : _GEN_9024; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9185 = 8'h3b == total_offset_27 ? field_byte_27 : _GEN_9025; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9186 = 8'h3c == total_offset_27 ? field_byte_27 : _GEN_9026; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9187 = 8'h3d == total_offset_27 ? field_byte_27 : _GEN_9027; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9188 = 8'h3e == total_offset_27 ? field_byte_27 : _GEN_9028; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9189 = 8'h3f == total_offset_27 ? field_byte_27 : _GEN_9029; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9190 = 8'h40 == total_offset_27 ? field_byte_27 : _GEN_9030; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9191 = 8'h41 == total_offset_27 ? field_byte_27 : _GEN_9031; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9192 = 8'h42 == total_offset_27 ? field_byte_27 : _GEN_9032; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9193 = 8'h43 == total_offset_27 ? field_byte_27 : _GEN_9033; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9194 = 8'h44 == total_offset_27 ? field_byte_27 : _GEN_9034; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9195 = 8'h45 == total_offset_27 ? field_byte_27 : _GEN_9035; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9196 = 8'h46 == total_offset_27 ? field_byte_27 : _GEN_9036; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9197 = 8'h47 == total_offset_27 ? field_byte_27 : _GEN_9037; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9198 = 8'h48 == total_offset_27 ? field_byte_27 : _GEN_9038; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9199 = 8'h49 == total_offset_27 ? field_byte_27 : _GEN_9039; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9200 = 8'h4a == total_offset_27 ? field_byte_27 : _GEN_9040; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9201 = 8'h4b == total_offset_27 ? field_byte_27 : _GEN_9041; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9202 = 8'h4c == total_offset_27 ? field_byte_27 : _GEN_9042; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9203 = 8'h4d == total_offset_27 ? field_byte_27 : _GEN_9043; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9204 = 8'h4e == total_offset_27 ? field_byte_27 : _GEN_9044; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9205 = 8'h4f == total_offset_27 ? field_byte_27 : _GEN_9045; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9206 = 8'h50 == total_offset_27 ? field_byte_27 : _GEN_9046; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9207 = 8'h51 == total_offset_27 ? field_byte_27 : _GEN_9047; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9208 = 8'h52 == total_offset_27 ? field_byte_27 : _GEN_9048; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9209 = 8'h53 == total_offset_27 ? field_byte_27 : _GEN_9049; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9210 = 8'h54 == total_offset_27 ? field_byte_27 : _GEN_9050; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9211 = 8'h55 == total_offset_27 ? field_byte_27 : _GEN_9051; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9212 = 8'h56 == total_offset_27 ? field_byte_27 : _GEN_9052; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9213 = 8'h57 == total_offset_27 ? field_byte_27 : _GEN_9053; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9214 = 8'h58 == total_offset_27 ? field_byte_27 : _GEN_9054; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9215 = 8'h59 == total_offset_27 ? field_byte_27 : _GEN_9055; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9216 = 8'h5a == total_offset_27 ? field_byte_27 : _GEN_9056; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9217 = 8'h5b == total_offset_27 ? field_byte_27 : _GEN_9057; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9218 = 8'h5c == total_offset_27 ? field_byte_27 : _GEN_9058; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9219 = 8'h5d == total_offset_27 ? field_byte_27 : _GEN_9059; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9220 = 8'h5e == total_offset_27 ? field_byte_27 : _GEN_9060; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9221 = 8'h5f == total_offset_27 ? field_byte_27 : _GEN_9061; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9222 = 8'h60 == total_offset_27 ? field_byte_27 : _GEN_9062; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9223 = 8'h61 == total_offset_27 ? field_byte_27 : _GEN_9063; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9224 = 8'h62 == total_offset_27 ? field_byte_27 : _GEN_9064; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9225 = 8'h63 == total_offset_27 ? field_byte_27 : _GEN_9065; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9226 = 8'h64 == total_offset_27 ? field_byte_27 : _GEN_9066; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9227 = 8'h65 == total_offset_27 ? field_byte_27 : _GEN_9067; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9228 = 8'h66 == total_offset_27 ? field_byte_27 : _GEN_9068; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9229 = 8'h67 == total_offset_27 ? field_byte_27 : _GEN_9069; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9230 = 8'h68 == total_offset_27 ? field_byte_27 : _GEN_9070; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9231 = 8'h69 == total_offset_27 ? field_byte_27 : _GEN_9071; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9232 = 8'h6a == total_offset_27 ? field_byte_27 : _GEN_9072; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9233 = 8'h6b == total_offset_27 ? field_byte_27 : _GEN_9073; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9234 = 8'h6c == total_offset_27 ? field_byte_27 : _GEN_9074; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9235 = 8'h6d == total_offset_27 ? field_byte_27 : _GEN_9075; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9236 = 8'h6e == total_offset_27 ? field_byte_27 : _GEN_9076; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9237 = 8'h6f == total_offset_27 ? field_byte_27 : _GEN_9077; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9238 = 8'h70 == total_offset_27 ? field_byte_27 : _GEN_9078; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9239 = 8'h71 == total_offset_27 ? field_byte_27 : _GEN_9079; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9240 = 8'h72 == total_offset_27 ? field_byte_27 : _GEN_9080; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9241 = 8'h73 == total_offset_27 ? field_byte_27 : _GEN_9081; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9242 = 8'h74 == total_offset_27 ? field_byte_27 : _GEN_9082; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9243 = 8'h75 == total_offset_27 ? field_byte_27 : _GEN_9083; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9244 = 8'h76 == total_offset_27 ? field_byte_27 : _GEN_9084; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9245 = 8'h77 == total_offset_27 ? field_byte_27 : _GEN_9085; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9246 = 8'h78 == total_offset_27 ? field_byte_27 : _GEN_9086; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9247 = 8'h79 == total_offset_27 ? field_byte_27 : _GEN_9087; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9248 = 8'h7a == total_offset_27 ? field_byte_27 : _GEN_9088; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9249 = 8'h7b == total_offset_27 ? field_byte_27 : _GEN_9089; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9250 = 8'h7c == total_offset_27 ? field_byte_27 : _GEN_9090; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9251 = 8'h7d == total_offset_27 ? field_byte_27 : _GEN_9091; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9252 = 8'h7e == total_offset_27 ? field_byte_27 : _GEN_9092; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9253 = 8'h7f == total_offset_27 ? field_byte_27 : _GEN_9093; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9254 = 8'h80 == total_offset_27 ? field_byte_27 : _GEN_9094; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9255 = 8'h81 == total_offset_27 ? field_byte_27 : _GEN_9095; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9256 = 8'h82 == total_offset_27 ? field_byte_27 : _GEN_9096; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9257 = 8'h83 == total_offset_27 ? field_byte_27 : _GEN_9097; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9258 = 8'h84 == total_offset_27 ? field_byte_27 : _GEN_9098; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9259 = 8'h85 == total_offset_27 ? field_byte_27 : _GEN_9099; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9260 = 8'h86 == total_offset_27 ? field_byte_27 : _GEN_9100; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9261 = 8'h87 == total_offset_27 ? field_byte_27 : _GEN_9101; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9262 = 8'h88 == total_offset_27 ? field_byte_27 : _GEN_9102; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9263 = 8'h89 == total_offset_27 ? field_byte_27 : _GEN_9103; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9264 = 8'h8a == total_offset_27 ? field_byte_27 : _GEN_9104; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9265 = 8'h8b == total_offset_27 ? field_byte_27 : _GEN_9105; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9266 = 8'h8c == total_offset_27 ? field_byte_27 : _GEN_9106; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9267 = 8'h8d == total_offset_27 ? field_byte_27 : _GEN_9107; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9268 = 8'h8e == total_offset_27 ? field_byte_27 : _GEN_9108; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9269 = 8'h8f == total_offset_27 ? field_byte_27 : _GEN_9109; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9270 = 8'h90 == total_offset_27 ? field_byte_27 : _GEN_9110; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9271 = 8'h91 == total_offset_27 ? field_byte_27 : _GEN_9111; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9272 = 8'h92 == total_offset_27 ? field_byte_27 : _GEN_9112; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9273 = 8'h93 == total_offset_27 ? field_byte_27 : _GEN_9113; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9274 = 8'h94 == total_offset_27 ? field_byte_27 : _GEN_9114; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9275 = 8'h95 == total_offset_27 ? field_byte_27 : _GEN_9115; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9276 = 8'h96 == total_offset_27 ? field_byte_27 : _GEN_9116; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9277 = 8'h97 == total_offset_27 ? field_byte_27 : _GEN_9117; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9278 = 8'h98 == total_offset_27 ? field_byte_27 : _GEN_9118; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9279 = 8'h99 == total_offset_27 ? field_byte_27 : _GEN_9119; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9280 = 8'h9a == total_offset_27 ? field_byte_27 : _GEN_9120; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9281 = 8'h9b == total_offset_27 ? field_byte_27 : _GEN_9121; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9282 = 8'h9c == total_offset_27 ? field_byte_27 : _GEN_9122; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9283 = 8'h9d == total_offset_27 ? field_byte_27 : _GEN_9123; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9284 = 8'h9e == total_offset_27 ? field_byte_27 : _GEN_9124; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9285 = 8'h9f == total_offset_27 ? field_byte_27 : _GEN_9125; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9286 = 8'h3 < length_3 ? _GEN_9126 : _GEN_8966; // @[executor.scala 308:60]
  wire [7:0] _GEN_9287 = 8'h3 < length_3 ? _GEN_9127 : _GEN_8967; // @[executor.scala 308:60]
  wire [7:0] _GEN_9288 = 8'h3 < length_3 ? _GEN_9128 : _GEN_8968; // @[executor.scala 308:60]
  wire [7:0] _GEN_9289 = 8'h3 < length_3 ? _GEN_9129 : _GEN_8969; // @[executor.scala 308:60]
  wire [7:0] _GEN_9290 = 8'h3 < length_3 ? _GEN_9130 : _GEN_8970; // @[executor.scala 308:60]
  wire [7:0] _GEN_9291 = 8'h3 < length_3 ? _GEN_9131 : _GEN_8971; // @[executor.scala 308:60]
  wire [7:0] _GEN_9292 = 8'h3 < length_3 ? _GEN_9132 : _GEN_8972; // @[executor.scala 308:60]
  wire [7:0] _GEN_9293 = 8'h3 < length_3 ? _GEN_9133 : _GEN_8973; // @[executor.scala 308:60]
  wire [7:0] _GEN_9294 = 8'h3 < length_3 ? _GEN_9134 : _GEN_8974; // @[executor.scala 308:60]
  wire [7:0] _GEN_9295 = 8'h3 < length_3 ? _GEN_9135 : _GEN_8975; // @[executor.scala 308:60]
  wire [7:0] _GEN_9296 = 8'h3 < length_3 ? _GEN_9136 : _GEN_8976; // @[executor.scala 308:60]
  wire [7:0] _GEN_9297 = 8'h3 < length_3 ? _GEN_9137 : _GEN_8977; // @[executor.scala 308:60]
  wire [7:0] _GEN_9298 = 8'h3 < length_3 ? _GEN_9138 : _GEN_8978; // @[executor.scala 308:60]
  wire [7:0] _GEN_9299 = 8'h3 < length_3 ? _GEN_9139 : _GEN_8979; // @[executor.scala 308:60]
  wire [7:0] _GEN_9300 = 8'h3 < length_3 ? _GEN_9140 : _GEN_8980; // @[executor.scala 308:60]
  wire [7:0] _GEN_9301 = 8'h3 < length_3 ? _GEN_9141 : _GEN_8981; // @[executor.scala 308:60]
  wire [7:0] _GEN_9302 = 8'h3 < length_3 ? _GEN_9142 : _GEN_8982; // @[executor.scala 308:60]
  wire [7:0] _GEN_9303 = 8'h3 < length_3 ? _GEN_9143 : _GEN_8983; // @[executor.scala 308:60]
  wire [7:0] _GEN_9304 = 8'h3 < length_3 ? _GEN_9144 : _GEN_8984; // @[executor.scala 308:60]
  wire [7:0] _GEN_9305 = 8'h3 < length_3 ? _GEN_9145 : _GEN_8985; // @[executor.scala 308:60]
  wire [7:0] _GEN_9306 = 8'h3 < length_3 ? _GEN_9146 : _GEN_8986; // @[executor.scala 308:60]
  wire [7:0] _GEN_9307 = 8'h3 < length_3 ? _GEN_9147 : _GEN_8987; // @[executor.scala 308:60]
  wire [7:0] _GEN_9308 = 8'h3 < length_3 ? _GEN_9148 : _GEN_8988; // @[executor.scala 308:60]
  wire [7:0] _GEN_9309 = 8'h3 < length_3 ? _GEN_9149 : _GEN_8989; // @[executor.scala 308:60]
  wire [7:0] _GEN_9310 = 8'h3 < length_3 ? _GEN_9150 : _GEN_8990; // @[executor.scala 308:60]
  wire [7:0] _GEN_9311 = 8'h3 < length_3 ? _GEN_9151 : _GEN_8991; // @[executor.scala 308:60]
  wire [7:0] _GEN_9312 = 8'h3 < length_3 ? _GEN_9152 : _GEN_8992; // @[executor.scala 308:60]
  wire [7:0] _GEN_9313 = 8'h3 < length_3 ? _GEN_9153 : _GEN_8993; // @[executor.scala 308:60]
  wire [7:0] _GEN_9314 = 8'h3 < length_3 ? _GEN_9154 : _GEN_8994; // @[executor.scala 308:60]
  wire [7:0] _GEN_9315 = 8'h3 < length_3 ? _GEN_9155 : _GEN_8995; // @[executor.scala 308:60]
  wire [7:0] _GEN_9316 = 8'h3 < length_3 ? _GEN_9156 : _GEN_8996; // @[executor.scala 308:60]
  wire [7:0] _GEN_9317 = 8'h3 < length_3 ? _GEN_9157 : _GEN_8997; // @[executor.scala 308:60]
  wire [7:0] _GEN_9318 = 8'h3 < length_3 ? _GEN_9158 : _GEN_8998; // @[executor.scala 308:60]
  wire [7:0] _GEN_9319 = 8'h3 < length_3 ? _GEN_9159 : _GEN_8999; // @[executor.scala 308:60]
  wire [7:0] _GEN_9320 = 8'h3 < length_3 ? _GEN_9160 : _GEN_9000; // @[executor.scala 308:60]
  wire [7:0] _GEN_9321 = 8'h3 < length_3 ? _GEN_9161 : _GEN_9001; // @[executor.scala 308:60]
  wire [7:0] _GEN_9322 = 8'h3 < length_3 ? _GEN_9162 : _GEN_9002; // @[executor.scala 308:60]
  wire [7:0] _GEN_9323 = 8'h3 < length_3 ? _GEN_9163 : _GEN_9003; // @[executor.scala 308:60]
  wire [7:0] _GEN_9324 = 8'h3 < length_3 ? _GEN_9164 : _GEN_9004; // @[executor.scala 308:60]
  wire [7:0] _GEN_9325 = 8'h3 < length_3 ? _GEN_9165 : _GEN_9005; // @[executor.scala 308:60]
  wire [7:0] _GEN_9326 = 8'h3 < length_3 ? _GEN_9166 : _GEN_9006; // @[executor.scala 308:60]
  wire [7:0] _GEN_9327 = 8'h3 < length_3 ? _GEN_9167 : _GEN_9007; // @[executor.scala 308:60]
  wire [7:0] _GEN_9328 = 8'h3 < length_3 ? _GEN_9168 : _GEN_9008; // @[executor.scala 308:60]
  wire [7:0] _GEN_9329 = 8'h3 < length_3 ? _GEN_9169 : _GEN_9009; // @[executor.scala 308:60]
  wire [7:0] _GEN_9330 = 8'h3 < length_3 ? _GEN_9170 : _GEN_9010; // @[executor.scala 308:60]
  wire [7:0] _GEN_9331 = 8'h3 < length_3 ? _GEN_9171 : _GEN_9011; // @[executor.scala 308:60]
  wire [7:0] _GEN_9332 = 8'h3 < length_3 ? _GEN_9172 : _GEN_9012; // @[executor.scala 308:60]
  wire [7:0] _GEN_9333 = 8'h3 < length_3 ? _GEN_9173 : _GEN_9013; // @[executor.scala 308:60]
  wire [7:0] _GEN_9334 = 8'h3 < length_3 ? _GEN_9174 : _GEN_9014; // @[executor.scala 308:60]
  wire [7:0] _GEN_9335 = 8'h3 < length_3 ? _GEN_9175 : _GEN_9015; // @[executor.scala 308:60]
  wire [7:0] _GEN_9336 = 8'h3 < length_3 ? _GEN_9176 : _GEN_9016; // @[executor.scala 308:60]
  wire [7:0] _GEN_9337 = 8'h3 < length_3 ? _GEN_9177 : _GEN_9017; // @[executor.scala 308:60]
  wire [7:0] _GEN_9338 = 8'h3 < length_3 ? _GEN_9178 : _GEN_9018; // @[executor.scala 308:60]
  wire [7:0] _GEN_9339 = 8'h3 < length_3 ? _GEN_9179 : _GEN_9019; // @[executor.scala 308:60]
  wire [7:0] _GEN_9340 = 8'h3 < length_3 ? _GEN_9180 : _GEN_9020; // @[executor.scala 308:60]
  wire [7:0] _GEN_9341 = 8'h3 < length_3 ? _GEN_9181 : _GEN_9021; // @[executor.scala 308:60]
  wire [7:0] _GEN_9342 = 8'h3 < length_3 ? _GEN_9182 : _GEN_9022; // @[executor.scala 308:60]
  wire [7:0] _GEN_9343 = 8'h3 < length_3 ? _GEN_9183 : _GEN_9023; // @[executor.scala 308:60]
  wire [7:0] _GEN_9344 = 8'h3 < length_3 ? _GEN_9184 : _GEN_9024; // @[executor.scala 308:60]
  wire [7:0] _GEN_9345 = 8'h3 < length_3 ? _GEN_9185 : _GEN_9025; // @[executor.scala 308:60]
  wire [7:0] _GEN_9346 = 8'h3 < length_3 ? _GEN_9186 : _GEN_9026; // @[executor.scala 308:60]
  wire [7:0] _GEN_9347 = 8'h3 < length_3 ? _GEN_9187 : _GEN_9027; // @[executor.scala 308:60]
  wire [7:0] _GEN_9348 = 8'h3 < length_3 ? _GEN_9188 : _GEN_9028; // @[executor.scala 308:60]
  wire [7:0] _GEN_9349 = 8'h3 < length_3 ? _GEN_9189 : _GEN_9029; // @[executor.scala 308:60]
  wire [7:0] _GEN_9350 = 8'h3 < length_3 ? _GEN_9190 : _GEN_9030; // @[executor.scala 308:60]
  wire [7:0] _GEN_9351 = 8'h3 < length_3 ? _GEN_9191 : _GEN_9031; // @[executor.scala 308:60]
  wire [7:0] _GEN_9352 = 8'h3 < length_3 ? _GEN_9192 : _GEN_9032; // @[executor.scala 308:60]
  wire [7:0] _GEN_9353 = 8'h3 < length_3 ? _GEN_9193 : _GEN_9033; // @[executor.scala 308:60]
  wire [7:0] _GEN_9354 = 8'h3 < length_3 ? _GEN_9194 : _GEN_9034; // @[executor.scala 308:60]
  wire [7:0] _GEN_9355 = 8'h3 < length_3 ? _GEN_9195 : _GEN_9035; // @[executor.scala 308:60]
  wire [7:0] _GEN_9356 = 8'h3 < length_3 ? _GEN_9196 : _GEN_9036; // @[executor.scala 308:60]
  wire [7:0] _GEN_9357 = 8'h3 < length_3 ? _GEN_9197 : _GEN_9037; // @[executor.scala 308:60]
  wire [7:0] _GEN_9358 = 8'h3 < length_3 ? _GEN_9198 : _GEN_9038; // @[executor.scala 308:60]
  wire [7:0] _GEN_9359 = 8'h3 < length_3 ? _GEN_9199 : _GEN_9039; // @[executor.scala 308:60]
  wire [7:0] _GEN_9360 = 8'h3 < length_3 ? _GEN_9200 : _GEN_9040; // @[executor.scala 308:60]
  wire [7:0] _GEN_9361 = 8'h3 < length_3 ? _GEN_9201 : _GEN_9041; // @[executor.scala 308:60]
  wire [7:0] _GEN_9362 = 8'h3 < length_3 ? _GEN_9202 : _GEN_9042; // @[executor.scala 308:60]
  wire [7:0] _GEN_9363 = 8'h3 < length_3 ? _GEN_9203 : _GEN_9043; // @[executor.scala 308:60]
  wire [7:0] _GEN_9364 = 8'h3 < length_3 ? _GEN_9204 : _GEN_9044; // @[executor.scala 308:60]
  wire [7:0] _GEN_9365 = 8'h3 < length_3 ? _GEN_9205 : _GEN_9045; // @[executor.scala 308:60]
  wire [7:0] _GEN_9366 = 8'h3 < length_3 ? _GEN_9206 : _GEN_9046; // @[executor.scala 308:60]
  wire [7:0] _GEN_9367 = 8'h3 < length_3 ? _GEN_9207 : _GEN_9047; // @[executor.scala 308:60]
  wire [7:0] _GEN_9368 = 8'h3 < length_3 ? _GEN_9208 : _GEN_9048; // @[executor.scala 308:60]
  wire [7:0] _GEN_9369 = 8'h3 < length_3 ? _GEN_9209 : _GEN_9049; // @[executor.scala 308:60]
  wire [7:0] _GEN_9370 = 8'h3 < length_3 ? _GEN_9210 : _GEN_9050; // @[executor.scala 308:60]
  wire [7:0] _GEN_9371 = 8'h3 < length_3 ? _GEN_9211 : _GEN_9051; // @[executor.scala 308:60]
  wire [7:0] _GEN_9372 = 8'h3 < length_3 ? _GEN_9212 : _GEN_9052; // @[executor.scala 308:60]
  wire [7:0] _GEN_9373 = 8'h3 < length_3 ? _GEN_9213 : _GEN_9053; // @[executor.scala 308:60]
  wire [7:0] _GEN_9374 = 8'h3 < length_3 ? _GEN_9214 : _GEN_9054; // @[executor.scala 308:60]
  wire [7:0] _GEN_9375 = 8'h3 < length_3 ? _GEN_9215 : _GEN_9055; // @[executor.scala 308:60]
  wire [7:0] _GEN_9376 = 8'h3 < length_3 ? _GEN_9216 : _GEN_9056; // @[executor.scala 308:60]
  wire [7:0] _GEN_9377 = 8'h3 < length_3 ? _GEN_9217 : _GEN_9057; // @[executor.scala 308:60]
  wire [7:0] _GEN_9378 = 8'h3 < length_3 ? _GEN_9218 : _GEN_9058; // @[executor.scala 308:60]
  wire [7:0] _GEN_9379 = 8'h3 < length_3 ? _GEN_9219 : _GEN_9059; // @[executor.scala 308:60]
  wire [7:0] _GEN_9380 = 8'h3 < length_3 ? _GEN_9220 : _GEN_9060; // @[executor.scala 308:60]
  wire [7:0] _GEN_9381 = 8'h3 < length_3 ? _GEN_9221 : _GEN_9061; // @[executor.scala 308:60]
  wire [7:0] _GEN_9382 = 8'h3 < length_3 ? _GEN_9222 : _GEN_9062; // @[executor.scala 308:60]
  wire [7:0] _GEN_9383 = 8'h3 < length_3 ? _GEN_9223 : _GEN_9063; // @[executor.scala 308:60]
  wire [7:0] _GEN_9384 = 8'h3 < length_3 ? _GEN_9224 : _GEN_9064; // @[executor.scala 308:60]
  wire [7:0] _GEN_9385 = 8'h3 < length_3 ? _GEN_9225 : _GEN_9065; // @[executor.scala 308:60]
  wire [7:0] _GEN_9386 = 8'h3 < length_3 ? _GEN_9226 : _GEN_9066; // @[executor.scala 308:60]
  wire [7:0] _GEN_9387 = 8'h3 < length_3 ? _GEN_9227 : _GEN_9067; // @[executor.scala 308:60]
  wire [7:0] _GEN_9388 = 8'h3 < length_3 ? _GEN_9228 : _GEN_9068; // @[executor.scala 308:60]
  wire [7:0] _GEN_9389 = 8'h3 < length_3 ? _GEN_9229 : _GEN_9069; // @[executor.scala 308:60]
  wire [7:0] _GEN_9390 = 8'h3 < length_3 ? _GEN_9230 : _GEN_9070; // @[executor.scala 308:60]
  wire [7:0] _GEN_9391 = 8'h3 < length_3 ? _GEN_9231 : _GEN_9071; // @[executor.scala 308:60]
  wire [7:0] _GEN_9392 = 8'h3 < length_3 ? _GEN_9232 : _GEN_9072; // @[executor.scala 308:60]
  wire [7:0] _GEN_9393 = 8'h3 < length_3 ? _GEN_9233 : _GEN_9073; // @[executor.scala 308:60]
  wire [7:0] _GEN_9394 = 8'h3 < length_3 ? _GEN_9234 : _GEN_9074; // @[executor.scala 308:60]
  wire [7:0] _GEN_9395 = 8'h3 < length_3 ? _GEN_9235 : _GEN_9075; // @[executor.scala 308:60]
  wire [7:0] _GEN_9396 = 8'h3 < length_3 ? _GEN_9236 : _GEN_9076; // @[executor.scala 308:60]
  wire [7:0] _GEN_9397 = 8'h3 < length_3 ? _GEN_9237 : _GEN_9077; // @[executor.scala 308:60]
  wire [7:0] _GEN_9398 = 8'h3 < length_3 ? _GEN_9238 : _GEN_9078; // @[executor.scala 308:60]
  wire [7:0] _GEN_9399 = 8'h3 < length_3 ? _GEN_9239 : _GEN_9079; // @[executor.scala 308:60]
  wire [7:0] _GEN_9400 = 8'h3 < length_3 ? _GEN_9240 : _GEN_9080; // @[executor.scala 308:60]
  wire [7:0] _GEN_9401 = 8'h3 < length_3 ? _GEN_9241 : _GEN_9081; // @[executor.scala 308:60]
  wire [7:0] _GEN_9402 = 8'h3 < length_3 ? _GEN_9242 : _GEN_9082; // @[executor.scala 308:60]
  wire [7:0] _GEN_9403 = 8'h3 < length_3 ? _GEN_9243 : _GEN_9083; // @[executor.scala 308:60]
  wire [7:0] _GEN_9404 = 8'h3 < length_3 ? _GEN_9244 : _GEN_9084; // @[executor.scala 308:60]
  wire [7:0] _GEN_9405 = 8'h3 < length_3 ? _GEN_9245 : _GEN_9085; // @[executor.scala 308:60]
  wire [7:0] _GEN_9406 = 8'h3 < length_3 ? _GEN_9246 : _GEN_9086; // @[executor.scala 308:60]
  wire [7:0] _GEN_9407 = 8'h3 < length_3 ? _GEN_9247 : _GEN_9087; // @[executor.scala 308:60]
  wire [7:0] _GEN_9408 = 8'h3 < length_3 ? _GEN_9248 : _GEN_9088; // @[executor.scala 308:60]
  wire [7:0] _GEN_9409 = 8'h3 < length_3 ? _GEN_9249 : _GEN_9089; // @[executor.scala 308:60]
  wire [7:0] _GEN_9410 = 8'h3 < length_3 ? _GEN_9250 : _GEN_9090; // @[executor.scala 308:60]
  wire [7:0] _GEN_9411 = 8'h3 < length_3 ? _GEN_9251 : _GEN_9091; // @[executor.scala 308:60]
  wire [7:0] _GEN_9412 = 8'h3 < length_3 ? _GEN_9252 : _GEN_9092; // @[executor.scala 308:60]
  wire [7:0] _GEN_9413 = 8'h3 < length_3 ? _GEN_9253 : _GEN_9093; // @[executor.scala 308:60]
  wire [7:0] _GEN_9414 = 8'h3 < length_3 ? _GEN_9254 : _GEN_9094; // @[executor.scala 308:60]
  wire [7:0] _GEN_9415 = 8'h3 < length_3 ? _GEN_9255 : _GEN_9095; // @[executor.scala 308:60]
  wire [7:0] _GEN_9416 = 8'h3 < length_3 ? _GEN_9256 : _GEN_9096; // @[executor.scala 308:60]
  wire [7:0] _GEN_9417 = 8'h3 < length_3 ? _GEN_9257 : _GEN_9097; // @[executor.scala 308:60]
  wire [7:0] _GEN_9418 = 8'h3 < length_3 ? _GEN_9258 : _GEN_9098; // @[executor.scala 308:60]
  wire [7:0] _GEN_9419 = 8'h3 < length_3 ? _GEN_9259 : _GEN_9099; // @[executor.scala 308:60]
  wire [7:0] _GEN_9420 = 8'h3 < length_3 ? _GEN_9260 : _GEN_9100; // @[executor.scala 308:60]
  wire [7:0] _GEN_9421 = 8'h3 < length_3 ? _GEN_9261 : _GEN_9101; // @[executor.scala 308:60]
  wire [7:0] _GEN_9422 = 8'h3 < length_3 ? _GEN_9262 : _GEN_9102; // @[executor.scala 308:60]
  wire [7:0] _GEN_9423 = 8'h3 < length_3 ? _GEN_9263 : _GEN_9103; // @[executor.scala 308:60]
  wire [7:0] _GEN_9424 = 8'h3 < length_3 ? _GEN_9264 : _GEN_9104; // @[executor.scala 308:60]
  wire [7:0] _GEN_9425 = 8'h3 < length_3 ? _GEN_9265 : _GEN_9105; // @[executor.scala 308:60]
  wire [7:0] _GEN_9426 = 8'h3 < length_3 ? _GEN_9266 : _GEN_9106; // @[executor.scala 308:60]
  wire [7:0] _GEN_9427 = 8'h3 < length_3 ? _GEN_9267 : _GEN_9107; // @[executor.scala 308:60]
  wire [7:0] _GEN_9428 = 8'h3 < length_3 ? _GEN_9268 : _GEN_9108; // @[executor.scala 308:60]
  wire [7:0] _GEN_9429 = 8'h3 < length_3 ? _GEN_9269 : _GEN_9109; // @[executor.scala 308:60]
  wire [7:0] _GEN_9430 = 8'h3 < length_3 ? _GEN_9270 : _GEN_9110; // @[executor.scala 308:60]
  wire [7:0] _GEN_9431 = 8'h3 < length_3 ? _GEN_9271 : _GEN_9111; // @[executor.scala 308:60]
  wire [7:0] _GEN_9432 = 8'h3 < length_3 ? _GEN_9272 : _GEN_9112; // @[executor.scala 308:60]
  wire [7:0] _GEN_9433 = 8'h3 < length_3 ? _GEN_9273 : _GEN_9113; // @[executor.scala 308:60]
  wire [7:0] _GEN_9434 = 8'h3 < length_3 ? _GEN_9274 : _GEN_9114; // @[executor.scala 308:60]
  wire [7:0] _GEN_9435 = 8'h3 < length_3 ? _GEN_9275 : _GEN_9115; // @[executor.scala 308:60]
  wire [7:0] _GEN_9436 = 8'h3 < length_3 ? _GEN_9276 : _GEN_9116; // @[executor.scala 308:60]
  wire [7:0] _GEN_9437 = 8'h3 < length_3 ? _GEN_9277 : _GEN_9117; // @[executor.scala 308:60]
  wire [7:0] _GEN_9438 = 8'h3 < length_3 ? _GEN_9278 : _GEN_9118; // @[executor.scala 308:60]
  wire [7:0] _GEN_9439 = 8'h3 < length_3 ? _GEN_9279 : _GEN_9119; // @[executor.scala 308:60]
  wire [7:0] _GEN_9440 = 8'h3 < length_3 ? _GEN_9280 : _GEN_9120; // @[executor.scala 308:60]
  wire [7:0] _GEN_9441 = 8'h3 < length_3 ? _GEN_9281 : _GEN_9121; // @[executor.scala 308:60]
  wire [7:0] _GEN_9442 = 8'h3 < length_3 ? _GEN_9282 : _GEN_9122; // @[executor.scala 308:60]
  wire [7:0] _GEN_9443 = 8'h3 < length_3 ? _GEN_9283 : _GEN_9123; // @[executor.scala 308:60]
  wire [7:0] _GEN_9444 = 8'h3 < length_3 ? _GEN_9284 : _GEN_9124; // @[executor.scala 308:60]
  wire [7:0] _GEN_9445 = 8'h3 < length_3 ? _GEN_9285 : _GEN_9125; // @[executor.scala 308:60]
  wire [7:0] field_byte_28 = field_3[31:24]; // @[executor.scala 305:57]
  wire [7:0] total_offset_28 = offset_3 + 8'h4; // @[executor.scala 307:57]
  wire [7:0] _GEN_9446 = 8'h0 == total_offset_28 ? field_byte_28 : _GEN_9286; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9447 = 8'h1 == total_offset_28 ? field_byte_28 : _GEN_9287; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9448 = 8'h2 == total_offset_28 ? field_byte_28 : _GEN_9288; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9449 = 8'h3 == total_offset_28 ? field_byte_28 : _GEN_9289; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9450 = 8'h4 == total_offset_28 ? field_byte_28 : _GEN_9290; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9451 = 8'h5 == total_offset_28 ? field_byte_28 : _GEN_9291; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9452 = 8'h6 == total_offset_28 ? field_byte_28 : _GEN_9292; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9453 = 8'h7 == total_offset_28 ? field_byte_28 : _GEN_9293; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9454 = 8'h8 == total_offset_28 ? field_byte_28 : _GEN_9294; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9455 = 8'h9 == total_offset_28 ? field_byte_28 : _GEN_9295; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9456 = 8'ha == total_offset_28 ? field_byte_28 : _GEN_9296; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9457 = 8'hb == total_offset_28 ? field_byte_28 : _GEN_9297; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9458 = 8'hc == total_offset_28 ? field_byte_28 : _GEN_9298; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9459 = 8'hd == total_offset_28 ? field_byte_28 : _GEN_9299; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9460 = 8'he == total_offset_28 ? field_byte_28 : _GEN_9300; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9461 = 8'hf == total_offset_28 ? field_byte_28 : _GEN_9301; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9462 = 8'h10 == total_offset_28 ? field_byte_28 : _GEN_9302; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9463 = 8'h11 == total_offset_28 ? field_byte_28 : _GEN_9303; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9464 = 8'h12 == total_offset_28 ? field_byte_28 : _GEN_9304; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9465 = 8'h13 == total_offset_28 ? field_byte_28 : _GEN_9305; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9466 = 8'h14 == total_offset_28 ? field_byte_28 : _GEN_9306; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9467 = 8'h15 == total_offset_28 ? field_byte_28 : _GEN_9307; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9468 = 8'h16 == total_offset_28 ? field_byte_28 : _GEN_9308; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9469 = 8'h17 == total_offset_28 ? field_byte_28 : _GEN_9309; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9470 = 8'h18 == total_offset_28 ? field_byte_28 : _GEN_9310; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9471 = 8'h19 == total_offset_28 ? field_byte_28 : _GEN_9311; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9472 = 8'h1a == total_offset_28 ? field_byte_28 : _GEN_9312; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9473 = 8'h1b == total_offset_28 ? field_byte_28 : _GEN_9313; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9474 = 8'h1c == total_offset_28 ? field_byte_28 : _GEN_9314; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9475 = 8'h1d == total_offset_28 ? field_byte_28 : _GEN_9315; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9476 = 8'h1e == total_offset_28 ? field_byte_28 : _GEN_9316; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9477 = 8'h1f == total_offset_28 ? field_byte_28 : _GEN_9317; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9478 = 8'h20 == total_offset_28 ? field_byte_28 : _GEN_9318; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9479 = 8'h21 == total_offset_28 ? field_byte_28 : _GEN_9319; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9480 = 8'h22 == total_offset_28 ? field_byte_28 : _GEN_9320; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9481 = 8'h23 == total_offset_28 ? field_byte_28 : _GEN_9321; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9482 = 8'h24 == total_offset_28 ? field_byte_28 : _GEN_9322; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9483 = 8'h25 == total_offset_28 ? field_byte_28 : _GEN_9323; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9484 = 8'h26 == total_offset_28 ? field_byte_28 : _GEN_9324; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9485 = 8'h27 == total_offset_28 ? field_byte_28 : _GEN_9325; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9486 = 8'h28 == total_offset_28 ? field_byte_28 : _GEN_9326; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9487 = 8'h29 == total_offset_28 ? field_byte_28 : _GEN_9327; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9488 = 8'h2a == total_offset_28 ? field_byte_28 : _GEN_9328; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9489 = 8'h2b == total_offset_28 ? field_byte_28 : _GEN_9329; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9490 = 8'h2c == total_offset_28 ? field_byte_28 : _GEN_9330; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9491 = 8'h2d == total_offset_28 ? field_byte_28 : _GEN_9331; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9492 = 8'h2e == total_offset_28 ? field_byte_28 : _GEN_9332; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9493 = 8'h2f == total_offset_28 ? field_byte_28 : _GEN_9333; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9494 = 8'h30 == total_offset_28 ? field_byte_28 : _GEN_9334; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9495 = 8'h31 == total_offset_28 ? field_byte_28 : _GEN_9335; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9496 = 8'h32 == total_offset_28 ? field_byte_28 : _GEN_9336; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9497 = 8'h33 == total_offset_28 ? field_byte_28 : _GEN_9337; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9498 = 8'h34 == total_offset_28 ? field_byte_28 : _GEN_9338; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9499 = 8'h35 == total_offset_28 ? field_byte_28 : _GEN_9339; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9500 = 8'h36 == total_offset_28 ? field_byte_28 : _GEN_9340; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9501 = 8'h37 == total_offset_28 ? field_byte_28 : _GEN_9341; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9502 = 8'h38 == total_offset_28 ? field_byte_28 : _GEN_9342; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9503 = 8'h39 == total_offset_28 ? field_byte_28 : _GEN_9343; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9504 = 8'h3a == total_offset_28 ? field_byte_28 : _GEN_9344; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9505 = 8'h3b == total_offset_28 ? field_byte_28 : _GEN_9345; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9506 = 8'h3c == total_offset_28 ? field_byte_28 : _GEN_9346; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9507 = 8'h3d == total_offset_28 ? field_byte_28 : _GEN_9347; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9508 = 8'h3e == total_offset_28 ? field_byte_28 : _GEN_9348; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9509 = 8'h3f == total_offset_28 ? field_byte_28 : _GEN_9349; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9510 = 8'h40 == total_offset_28 ? field_byte_28 : _GEN_9350; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9511 = 8'h41 == total_offset_28 ? field_byte_28 : _GEN_9351; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9512 = 8'h42 == total_offset_28 ? field_byte_28 : _GEN_9352; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9513 = 8'h43 == total_offset_28 ? field_byte_28 : _GEN_9353; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9514 = 8'h44 == total_offset_28 ? field_byte_28 : _GEN_9354; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9515 = 8'h45 == total_offset_28 ? field_byte_28 : _GEN_9355; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9516 = 8'h46 == total_offset_28 ? field_byte_28 : _GEN_9356; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9517 = 8'h47 == total_offset_28 ? field_byte_28 : _GEN_9357; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9518 = 8'h48 == total_offset_28 ? field_byte_28 : _GEN_9358; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9519 = 8'h49 == total_offset_28 ? field_byte_28 : _GEN_9359; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9520 = 8'h4a == total_offset_28 ? field_byte_28 : _GEN_9360; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9521 = 8'h4b == total_offset_28 ? field_byte_28 : _GEN_9361; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9522 = 8'h4c == total_offset_28 ? field_byte_28 : _GEN_9362; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9523 = 8'h4d == total_offset_28 ? field_byte_28 : _GEN_9363; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9524 = 8'h4e == total_offset_28 ? field_byte_28 : _GEN_9364; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9525 = 8'h4f == total_offset_28 ? field_byte_28 : _GEN_9365; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9526 = 8'h50 == total_offset_28 ? field_byte_28 : _GEN_9366; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9527 = 8'h51 == total_offset_28 ? field_byte_28 : _GEN_9367; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9528 = 8'h52 == total_offset_28 ? field_byte_28 : _GEN_9368; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9529 = 8'h53 == total_offset_28 ? field_byte_28 : _GEN_9369; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9530 = 8'h54 == total_offset_28 ? field_byte_28 : _GEN_9370; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9531 = 8'h55 == total_offset_28 ? field_byte_28 : _GEN_9371; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9532 = 8'h56 == total_offset_28 ? field_byte_28 : _GEN_9372; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9533 = 8'h57 == total_offset_28 ? field_byte_28 : _GEN_9373; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9534 = 8'h58 == total_offset_28 ? field_byte_28 : _GEN_9374; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9535 = 8'h59 == total_offset_28 ? field_byte_28 : _GEN_9375; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9536 = 8'h5a == total_offset_28 ? field_byte_28 : _GEN_9376; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9537 = 8'h5b == total_offset_28 ? field_byte_28 : _GEN_9377; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9538 = 8'h5c == total_offset_28 ? field_byte_28 : _GEN_9378; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9539 = 8'h5d == total_offset_28 ? field_byte_28 : _GEN_9379; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9540 = 8'h5e == total_offset_28 ? field_byte_28 : _GEN_9380; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9541 = 8'h5f == total_offset_28 ? field_byte_28 : _GEN_9381; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9542 = 8'h60 == total_offset_28 ? field_byte_28 : _GEN_9382; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9543 = 8'h61 == total_offset_28 ? field_byte_28 : _GEN_9383; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9544 = 8'h62 == total_offset_28 ? field_byte_28 : _GEN_9384; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9545 = 8'h63 == total_offset_28 ? field_byte_28 : _GEN_9385; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9546 = 8'h64 == total_offset_28 ? field_byte_28 : _GEN_9386; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9547 = 8'h65 == total_offset_28 ? field_byte_28 : _GEN_9387; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9548 = 8'h66 == total_offset_28 ? field_byte_28 : _GEN_9388; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9549 = 8'h67 == total_offset_28 ? field_byte_28 : _GEN_9389; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9550 = 8'h68 == total_offset_28 ? field_byte_28 : _GEN_9390; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9551 = 8'h69 == total_offset_28 ? field_byte_28 : _GEN_9391; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9552 = 8'h6a == total_offset_28 ? field_byte_28 : _GEN_9392; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9553 = 8'h6b == total_offset_28 ? field_byte_28 : _GEN_9393; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9554 = 8'h6c == total_offset_28 ? field_byte_28 : _GEN_9394; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9555 = 8'h6d == total_offset_28 ? field_byte_28 : _GEN_9395; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9556 = 8'h6e == total_offset_28 ? field_byte_28 : _GEN_9396; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9557 = 8'h6f == total_offset_28 ? field_byte_28 : _GEN_9397; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9558 = 8'h70 == total_offset_28 ? field_byte_28 : _GEN_9398; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9559 = 8'h71 == total_offset_28 ? field_byte_28 : _GEN_9399; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9560 = 8'h72 == total_offset_28 ? field_byte_28 : _GEN_9400; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9561 = 8'h73 == total_offset_28 ? field_byte_28 : _GEN_9401; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9562 = 8'h74 == total_offset_28 ? field_byte_28 : _GEN_9402; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9563 = 8'h75 == total_offset_28 ? field_byte_28 : _GEN_9403; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9564 = 8'h76 == total_offset_28 ? field_byte_28 : _GEN_9404; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9565 = 8'h77 == total_offset_28 ? field_byte_28 : _GEN_9405; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9566 = 8'h78 == total_offset_28 ? field_byte_28 : _GEN_9406; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9567 = 8'h79 == total_offset_28 ? field_byte_28 : _GEN_9407; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9568 = 8'h7a == total_offset_28 ? field_byte_28 : _GEN_9408; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9569 = 8'h7b == total_offset_28 ? field_byte_28 : _GEN_9409; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9570 = 8'h7c == total_offset_28 ? field_byte_28 : _GEN_9410; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9571 = 8'h7d == total_offset_28 ? field_byte_28 : _GEN_9411; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9572 = 8'h7e == total_offset_28 ? field_byte_28 : _GEN_9412; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9573 = 8'h7f == total_offset_28 ? field_byte_28 : _GEN_9413; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9574 = 8'h80 == total_offset_28 ? field_byte_28 : _GEN_9414; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9575 = 8'h81 == total_offset_28 ? field_byte_28 : _GEN_9415; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9576 = 8'h82 == total_offset_28 ? field_byte_28 : _GEN_9416; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9577 = 8'h83 == total_offset_28 ? field_byte_28 : _GEN_9417; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9578 = 8'h84 == total_offset_28 ? field_byte_28 : _GEN_9418; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9579 = 8'h85 == total_offset_28 ? field_byte_28 : _GEN_9419; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9580 = 8'h86 == total_offset_28 ? field_byte_28 : _GEN_9420; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9581 = 8'h87 == total_offset_28 ? field_byte_28 : _GEN_9421; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9582 = 8'h88 == total_offset_28 ? field_byte_28 : _GEN_9422; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9583 = 8'h89 == total_offset_28 ? field_byte_28 : _GEN_9423; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9584 = 8'h8a == total_offset_28 ? field_byte_28 : _GEN_9424; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9585 = 8'h8b == total_offset_28 ? field_byte_28 : _GEN_9425; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9586 = 8'h8c == total_offset_28 ? field_byte_28 : _GEN_9426; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9587 = 8'h8d == total_offset_28 ? field_byte_28 : _GEN_9427; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9588 = 8'h8e == total_offset_28 ? field_byte_28 : _GEN_9428; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9589 = 8'h8f == total_offset_28 ? field_byte_28 : _GEN_9429; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9590 = 8'h90 == total_offset_28 ? field_byte_28 : _GEN_9430; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9591 = 8'h91 == total_offset_28 ? field_byte_28 : _GEN_9431; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9592 = 8'h92 == total_offset_28 ? field_byte_28 : _GEN_9432; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9593 = 8'h93 == total_offset_28 ? field_byte_28 : _GEN_9433; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9594 = 8'h94 == total_offset_28 ? field_byte_28 : _GEN_9434; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9595 = 8'h95 == total_offset_28 ? field_byte_28 : _GEN_9435; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9596 = 8'h96 == total_offset_28 ? field_byte_28 : _GEN_9436; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9597 = 8'h97 == total_offset_28 ? field_byte_28 : _GEN_9437; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9598 = 8'h98 == total_offset_28 ? field_byte_28 : _GEN_9438; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9599 = 8'h99 == total_offset_28 ? field_byte_28 : _GEN_9439; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9600 = 8'h9a == total_offset_28 ? field_byte_28 : _GEN_9440; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9601 = 8'h9b == total_offset_28 ? field_byte_28 : _GEN_9441; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9602 = 8'h9c == total_offset_28 ? field_byte_28 : _GEN_9442; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9603 = 8'h9d == total_offset_28 ? field_byte_28 : _GEN_9443; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9604 = 8'h9e == total_offset_28 ? field_byte_28 : _GEN_9444; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9605 = 8'h9f == total_offset_28 ? field_byte_28 : _GEN_9445; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9606 = 8'h4 < length_3 ? _GEN_9446 : _GEN_9286; // @[executor.scala 308:60]
  wire [7:0] _GEN_9607 = 8'h4 < length_3 ? _GEN_9447 : _GEN_9287; // @[executor.scala 308:60]
  wire [7:0] _GEN_9608 = 8'h4 < length_3 ? _GEN_9448 : _GEN_9288; // @[executor.scala 308:60]
  wire [7:0] _GEN_9609 = 8'h4 < length_3 ? _GEN_9449 : _GEN_9289; // @[executor.scala 308:60]
  wire [7:0] _GEN_9610 = 8'h4 < length_3 ? _GEN_9450 : _GEN_9290; // @[executor.scala 308:60]
  wire [7:0] _GEN_9611 = 8'h4 < length_3 ? _GEN_9451 : _GEN_9291; // @[executor.scala 308:60]
  wire [7:0] _GEN_9612 = 8'h4 < length_3 ? _GEN_9452 : _GEN_9292; // @[executor.scala 308:60]
  wire [7:0] _GEN_9613 = 8'h4 < length_3 ? _GEN_9453 : _GEN_9293; // @[executor.scala 308:60]
  wire [7:0] _GEN_9614 = 8'h4 < length_3 ? _GEN_9454 : _GEN_9294; // @[executor.scala 308:60]
  wire [7:0] _GEN_9615 = 8'h4 < length_3 ? _GEN_9455 : _GEN_9295; // @[executor.scala 308:60]
  wire [7:0] _GEN_9616 = 8'h4 < length_3 ? _GEN_9456 : _GEN_9296; // @[executor.scala 308:60]
  wire [7:0] _GEN_9617 = 8'h4 < length_3 ? _GEN_9457 : _GEN_9297; // @[executor.scala 308:60]
  wire [7:0] _GEN_9618 = 8'h4 < length_3 ? _GEN_9458 : _GEN_9298; // @[executor.scala 308:60]
  wire [7:0] _GEN_9619 = 8'h4 < length_3 ? _GEN_9459 : _GEN_9299; // @[executor.scala 308:60]
  wire [7:0] _GEN_9620 = 8'h4 < length_3 ? _GEN_9460 : _GEN_9300; // @[executor.scala 308:60]
  wire [7:0] _GEN_9621 = 8'h4 < length_3 ? _GEN_9461 : _GEN_9301; // @[executor.scala 308:60]
  wire [7:0] _GEN_9622 = 8'h4 < length_3 ? _GEN_9462 : _GEN_9302; // @[executor.scala 308:60]
  wire [7:0] _GEN_9623 = 8'h4 < length_3 ? _GEN_9463 : _GEN_9303; // @[executor.scala 308:60]
  wire [7:0] _GEN_9624 = 8'h4 < length_3 ? _GEN_9464 : _GEN_9304; // @[executor.scala 308:60]
  wire [7:0] _GEN_9625 = 8'h4 < length_3 ? _GEN_9465 : _GEN_9305; // @[executor.scala 308:60]
  wire [7:0] _GEN_9626 = 8'h4 < length_3 ? _GEN_9466 : _GEN_9306; // @[executor.scala 308:60]
  wire [7:0] _GEN_9627 = 8'h4 < length_3 ? _GEN_9467 : _GEN_9307; // @[executor.scala 308:60]
  wire [7:0] _GEN_9628 = 8'h4 < length_3 ? _GEN_9468 : _GEN_9308; // @[executor.scala 308:60]
  wire [7:0] _GEN_9629 = 8'h4 < length_3 ? _GEN_9469 : _GEN_9309; // @[executor.scala 308:60]
  wire [7:0] _GEN_9630 = 8'h4 < length_3 ? _GEN_9470 : _GEN_9310; // @[executor.scala 308:60]
  wire [7:0] _GEN_9631 = 8'h4 < length_3 ? _GEN_9471 : _GEN_9311; // @[executor.scala 308:60]
  wire [7:0] _GEN_9632 = 8'h4 < length_3 ? _GEN_9472 : _GEN_9312; // @[executor.scala 308:60]
  wire [7:0] _GEN_9633 = 8'h4 < length_3 ? _GEN_9473 : _GEN_9313; // @[executor.scala 308:60]
  wire [7:0] _GEN_9634 = 8'h4 < length_3 ? _GEN_9474 : _GEN_9314; // @[executor.scala 308:60]
  wire [7:0] _GEN_9635 = 8'h4 < length_3 ? _GEN_9475 : _GEN_9315; // @[executor.scala 308:60]
  wire [7:0] _GEN_9636 = 8'h4 < length_3 ? _GEN_9476 : _GEN_9316; // @[executor.scala 308:60]
  wire [7:0] _GEN_9637 = 8'h4 < length_3 ? _GEN_9477 : _GEN_9317; // @[executor.scala 308:60]
  wire [7:0] _GEN_9638 = 8'h4 < length_3 ? _GEN_9478 : _GEN_9318; // @[executor.scala 308:60]
  wire [7:0] _GEN_9639 = 8'h4 < length_3 ? _GEN_9479 : _GEN_9319; // @[executor.scala 308:60]
  wire [7:0] _GEN_9640 = 8'h4 < length_3 ? _GEN_9480 : _GEN_9320; // @[executor.scala 308:60]
  wire [7:0] _GEN_9641 = 8'h4 < length_3 ? _GEN_9481 : _GEN_9321; // @[executor.scala 308:60]
  wire [7:0] _GEN_9642 = 8'h4 < length_3 ? _GEN_9482 : _GEN_9322; // @[executor.scala 308:60]
  wire [7:0] _GEN_9643 = 8'h4 < length_3 ? _GEN_9483 : _GEN_9323; // @[executor.scala 308:60]
  wire [7:0] _GEN_9644 = 8'h4 < length_3 ? _GEN_9484 : _GEN_9324; // @[executor.scala 308:60]
  wire [7:0] _GEN_9645 = 8'h4 < length_3 ? _GEN_9485 : _GEN_9325; // @[executor.scala 308:60]
  wire [7:0] _GEN_9646 = 8'h4 < length_3 ? _GEN_9486 : _GEN_9326; // @[executor.scala 308:60]
  wire [7:0] _GEN_9647 = 8'h4 < length_3 ? _GEN_9487 : _GEN_9327; // @[executor.scala 308:60]
  wire [7:0] _GEN_9648 = 8'h4 < length_3 ? _GEN_9488 : _GEN_9328; // @[executor.scala 308:60]
  wire [7:0] _GEN_9649 = 8'h4 < length_3 ? _GEN_9489 : _GEN_9329; // @[executor.scala 308:60]
  wire [7:0] _GEN_9650 = 8'h4 < length_3 ? _GEN_9490 : _GEN_9330; // @[executor.scala 308:60]
  wire [7:0] _GEN_9651 = 8'h4 < length_3 ? _GEN_9491 : _GEN_9331; // @[executor.scala 308:60]
  wire [7:0] _GEN_9652 = 8'h4 < length_3 ? _GEN_9492 : _GEN_9332; // @[executor.scala 308:60]
  wire [7:0] _GEN_9653 = 8'h4 < length_3 ? _GEN_9493 : _GEN_9333; // @[executor.scala 308:60]
  wire [7:0] _GEN_9654 = 8'h4 < length_3 ? _GEN_9494 : _GEN_9334; // @[executor.scala 308:60]
  wire [7:0] _GEN_9655 = 8'h4 < length_3 ? _GEN_9495 : _GEN_9335; // @[executor.scala 308:60]
  wire [7:0] _GEN_9656 = 8'h4 < length_3 ? _GEN_9496 : _GEN_9336; // @[executor.scala 308:60]
  wire [7:0] _GEN_9657 = 8'h4 < length_3 ? _GEN_9497 : _GEN_9337; // @[executor.scala 308:60]
  wire [7:0] _GEN_9658 = 8'h4 < length_3 ? _GEN_9498 : _GEN_9338; // @[executor.scala 308:60]
  wire [7:0] _GEN_9659 = 8'h4 < length_3 ? _GEN_9499 : _GEN_9339; // @[executor.scala 308:60]
  wire [7:0] _GEN_9660 = 8'h4 < length_3 ? _GEN_9500 : _GEN_9340; // @[executor.scala 308:60]
  wire [7:0] _GEN_9661 = 8'h4 < length_3 ? _GEN_9501 : _GEN_9341; // @[executor.scala 308:60]
  wire [7:0] _GEN_9662 = 8'h4 < length_3 ? _GEN_9502 : _GEN_9342; // @[executor.scala 308:60]
  wire [7:0] _GEN_9663 = 8'h4 < length_3 ? _GEN_9503 : _GEN_9343; // @[executor.scala 308:60]
  wire [7:0] _GEN_9664 = 8'h4 < length_3 ? _GEN_9504 : _GEN_9344; // @[executor.scala 308:60]
  wire [7:0] _GEN_9665 = 8'h4 < length_3 ? _GEN_9505 : _GEN_9345; // @[executor.scala 308:60]
  wire [7:0] _GEN_9666 = 8'h4 < length_3 ? _GEN_9506 : _GEN_9346; // @[executor.scala 308:60]
  wire [7:0] _GEN_9667 = 8'h4 < length_3 ? _GEN_9507 : _GEN_9347; // @[executor.scala 308:60]
  wire [7:0] _GEN_9668 = 8'h4 < length_3 ? _GEN_9508 : _GEN_9348; // @[executor.scala 308:60]
  wire [7:0] _GEN_9669 = 8'h4 < length_3 ? _GEN_9509 : _GEN_9349; // @[executor.scala 308:60]
  wire [7:0] _GEN_9670 = 8'h4 < length_3 ? _GEN_9510 : _GEN_9350; // @[executor.scala 308:60]
  wire [7:0] _GEN_9671 = 8'h4 < length_3 ? _GEN_9511 : _GEN_9351; // @[executor.scala 308:60]
  wire [7:0] _GEN_9672 = 8'h4 < length_3 ? _GEN_9512 : _GEN_9352; // @[executor.scala 308:60]
  wire [7:0] _GEN_9673 = 8'h4 < length_3 ? _GEN_9513 : _GEN_9353; // @[executor.scala 308:60]
  wire [7:0] _GEN_9674 = 8'h4 < length_3 ? _GEN_9514 : _GEN_9354; // @[executor.scala 308:60]
  wire [7:0] _GEN_9675 = 8'h4 < length_3 ? _GEN_9515 : _GEN_9355; // @[executor.scala 308:60]
  wire [7:0] _GEN_9676 = 8'h4 < length_3 ? _GEN_9516 : _GEN_9356; // @[executor.scala 308:60]
  wire [7:0] _GEN_9677 = 8'h4 < length_3 ? _GEN_9517 : _GEN_9357; // @[executor.scala 308:60]
  wire [7:0] _GEN_9678 = 8'h4 < length_3 ? _GEN_9518 : _GEN_9358; // @[executor.scala 308:60]
  wire [7:0] _GEN_9679 = 8'h4 < length_3 ? _GEN_9519 : _GEN_9359; // @[executor.scala 308:60]
  wire [7:0] _GEN_9680 = 8'h4 < length_3 ? _GEN_9520 : _GEN_9360; // @[executor.scala 308:60]
  wire [7:0] _GEN_9681 = 8'h4 < length_3 ? _GEN_9521 : _GEN_9361; // @[executor.scala 308:60]
  wire [7:0] _GEN_9682 = 8'h4 < length_3 ? _GEN_9522 : _GEN_9362; // @[executor.scala 308:60]
  wire [7:0] _GEN_9683 = 8'h4 < length_3 ? _GEN_9523 : _GEN_9363; // @[executor.scala 308:60]
  wire [7:0] _GEN_9684 = 8'h4 < length_3 ? _GEN_9524 : _GEN_9364; // @[executor.scala 308:60]
  wire [7:0] _GEN_9685 = 8'h4 < length_3 ? _GEN_9525 : _GEN_9365; // @[executor.scala 308:60]
  wire [7:0] _GEN_9686 = 8'h4 < length_3 ? _GEN_9526 : _GEN_9366; // @[executor.scala 308:60]
  wire [7:0] _GEN_9687 = 8'h4 < length_3 ? _GEN_9527 : _GEN_9367; // @[executor.scala 308:60]
  wire [7:0] _GEN_9688 = 8'h4 < length_3 ? _GEN_9528 : _GEN_9368; // @[executor.scala 308:60]
  wire [7:0] _GEN_9689 = 8'h4 < length_3 ? _GEN_9529 : _GEN_9369; // @[executor.scala 308:60]
  wire [7:0] _GEN_9690 = 8'h4 < length_3 ? _GEN_9530 : _GEN_9370; // @[executor.scala 308:60]
  wire [7:0] _GEN_9691 = 8'h4 < length_3 ? _GEN_9531 : _GEN_9371; // @[executor.scala 308:60]
  wire [7:0] _GEN_9692 = 8'h4 < length_3 ? _GEN_9532 : _GEN_9372; // @[executor.scala 308:60]
  wire [7:0] _GEN_9693 = 8'h4 < length_3 ? _GEN_9533 : _GEN_9373; // @[executor.scala 308:60]
  wire [7:0] _GEN_9694 = 8'h4 < length_3 ? _GEN_9534 : _GEN_9374; // @[executor.scala 308:60]
  wire [7:0] _GEN_9695 = 8'h4 < length_3 ? _GEN_9535 : _GEN_9375; // @[executor.scala 308:60]
  wire [7:0] _GEN_9696 = 8'h4 < length_3 ? _GEN_9536 : _GEN_9376; // @[executor.scala 308:60]
  wire [7:0] _GEN_9697 = 8'h4 < length_3 ? _GEN_9537 : _GEN_9377; // @[executor.scala 308:60]
  wire [7:0] _GEN_9698 = 8'h4 < length_3 ? _GEN_9538 : _GEN_9378; // @[executor.scala 308:60]
  wire [7:0] _GEN_9699 = 8'h4 < length_3 ? _GEN_9539 : _GEN_9379; // @[executor.scala 308:60]
  wire [7:0] _GEN_9700 = 8'h4 < length_3 ? _GEN_9540 : _GEN_9380; // @[executor.scala 308:60]
  wire [7:0] _GEN_9701 = 8'h4 < length_3 ? _GEN_9541 : _GEN_9381; // @[executor.scala 308:60]
  wire [7:0] _GEN_9702 = 8'h4 < length_3 ? _GEN_9542 : _GEN_9382; // @[executor.scala 308:60]
  wire [7:0] _GEN_9703 = 8'h4 < length_3 ? _GEN_9543 : _GEN_9383; // @[executor.scala 308:60]
  wire [7:0] _GEN_9704 = 8'h4 < length_3 ? _GEN_9544 : _GEN_9384; // @[executor.scala 308:60]
  wire [7:0] _GEN_9705 = 8'h4 < length_3 ? _GEN_9545 : _GEN_9385; // @[executor.scala 308:60]
  wire [7:0] _GEN_9706 = 8'h4 < length_3 ? _GEN_9546 : _GEN_9386; // @[executor.scala 308:60]
  wire [7:0] _GEN_9707 = 8'h4 < length_3 ? _GEN_9547 : _GEN_9387; // @[executor.scala 308:60]
  wire [7:0] _GEN_9708 = 8'h4 < length_3 ? _GEN_9548 : _GEN_9388; // @[executor.scala 308:60]
  wire [7:0] _GEN_9709 = 8'h4 < length_3 ? _GEN_9549 : _GEN_9389; // @[executor.scala 308:60]
  wire [7:0] _GEN_9710 = 8'h4 < length_3 ? _GEN_9550 : _GEN_9390; // @[executor.scala 308:60]
  wire [7:0] _GEN_9711 = 8'h4 < length_3 ? _GEN_9551 : _GEN_9391; // @[executor.scala 308:60]
  wire [7:0] _GEN_9712 = 8'h4 < length_3 ? _GEN_9552 : _GEN_9392; // @[executor.scala 308:60]
  wire [7:0] _GEN_9713 = 8'h4 < length_3 ? _GEN_9553 : _GEN_9393; // @[executor.scala 308:60]
  wire [7:0] _GEN_9714 = 8'h4 < length_3 ? _GEN_9554 : _GEN_9394; // @[executor.scala 308:60]
  wire [7:0] _GEN_9715 = 8'h4 < length_3 ? _GEN_9555 : _GEN_9395; // @[executor.scala 308:60]
  wire [7:0] _GEN_9716 = 8'h4 < length_3 ? _GEN_9556 : _GEN_9396; // @[executor.scala 308:60]
  wire [7:0] _GEN_9717 = 8'h4 < length_3 ? _GEN_9557 : _GEN_9397; // @[executor.scala 308:60]
  wire [7:0] _GEN_9718 = 8'h4 < length_3 ? _GEN_9558 : _GEN_9398; // @[executor.scala 308:60]
  wire [7:0] _GEN_9719 = 8'h4 < length_3 ? _GEN_9559 : _GEN_9399; // @[executor.scala 308:60]
  wire [7:0] _GEN_9720 = 8'h4 < length_3 ? _GEN_9560 : _GEN_9400; // @[executor.scala 308:60]
  wire [7:0] _GEN_9721 = 8'h4 < length_3 ? _GEN_9561 : _GEN_9401; // @[executor.scala 308:60]
  wire [7:0] _GEN_9722 = 8'h4 < length_3 ? _GEN_9562 : _GEN_9402; // @[executor.scala 308:60]
  wire [7:0] _GEN_9723 = 8'h4 < length_3 ? _GEN_9563 : _GEN_9403; // @[executor.scala 308:60]
  wire [7:0] _GEN_9724 = 8'h4 < length_3 ? _GEN_9564 : _GEN_9404; // @[executor.scala 308:60]
  wire [7:0] _GEN_9725 = 8'h4 < length_3 ? _GEN_9565 : _GEN_9405; // @[executor.scala 308:60]
  wire [7:0] _GEN_9726 = 8'h4 < length_3 ? _GEN_9566 : _GEN_9406; // @[executor.scala 308:60]
  wire [7:0] _GEN_9727 = 8'h4 < length_3 ? _GEN_9567 : _GEN_9407; // @[executor.scala 308:60]
  wire [7:0] _GEN_9728 = 8'h4 < length_3 ? _GEN_9568 : _GEN_9408; // @[executor.scala 308:60]
  wire [7:0] _GEN_9729 = 8'h4 < length_3 ? _GEN_9569 : _GEN_9409; // @[executor.scala 308:60]
  wire [7:0] _GEN_9730 = 8'h4 < length_3 ? _GEN_9570 : _GEN_9410; // @[executor.scala 308:60]
  wire [7:0] _GEN_9731 = 8'h4 < length_3 ? _GEN_9571 : _GEN_9411; // @[executor.scala 308:60]
  wire [7:0] _GEN_9732 = 8'h4 < length_3 ? _GEN_9572 : _GEN_9412; // @[executor.scala 308:60]
  wire [7:0] _GEN_9733 = 8'h4 < length_3 ? _GEN_9573 : _GEN_9413; // @[executor.scala 308:60]
  wire [7:0] _GEN_9734 = 8'h4 < length_3 ? _GEN_9574 : _GEN_9414; // @[executor.scala 308:60]
  wire [7:0] _GEN_9735 = 8'h4 < length_3 ? _GEN_9575 : _GEN_9415; // @[executor.scala 308:60]
  wire [7:0] _GEN_9736 = 8'h4 < length_3 ? _GEN_9576 : _GEN_9416; // @[executor.scala 308:60]
  wire [7:0] _GEN_9737 = 8'h4 < length_3 ? _GEN_9577 : _GEN_9417; // @[executor.scala 308:60]
  wire [7:0] _GEN_9738 = 8'h4 < length_3 ? _GEN_9578 : _GEN_9418; // @[executor.scala 308:60]
  wire [7:0] _GEN_9739 = 8'h4 < length_3 ? _GEN_9579 : _GEN_9419; // @[executor.scala 308:60]
  wire [7:0] _GEN_9740 = 8'h4 < length_3 ? _GEN_9580 : _GEN_9420; // @[executor.scala 308:60]
  wire [7:0] _GEN_9741 = 8'h4 < length_3 ? _GEN_9581 : _GEN_9421; // @[executor.scala 308:60]
  wire [7:0] _GEN_9742 = 8'h4 < length_3 ? _GEN_9582 : _GEN_9422; // @[executor.scala 308:60]
  wire [7:0] _GEN_9743 = 8'h4 < length_3 ? _GEN_9583 : _GEN_9423; // @[executor.scala 308:60]
  wire [7:0] _GEN_9744 = 8'h4 < length_3 ? _GEN_9584 : _GEN_9424; // @[executor.scala 308:60]
  wire [7:0] _GEN_9745 = 8'h4 < length_3 ? _GEN_9585 : _GEN_9425; // @[executor.scala 308:60]
  wire [7:0] _GEN_9746 = 8'h4 < length_3 ? _GEN_9586 : _GEN_9426; // @[executor.scala 308:60]
  wire [7:0] _GEN_9747 = 8'h4 < length_3 ? _GEN_9587 : _GEN_9427; // @[executor.scala 308:60]
  wire [7:0] _GEN_9748 = 8'h4 < length_3 ? _GEN_9588 : _GEN_9428; // @[executor.scala 308:60]
  wire [7:0] _GEN_9749 = 8'h4 < length_3 ? _GEN_9589 : _GEN_9429; // @[executor.scala 308:60]
  wire [7:0] _GEN_9750 = 8'h4 < length_3 ? _GEN_9590 : _GEN_9430; // @[executor.scala 308:60]
  wire [7:0] _GEN_9751 = 8'h4 < length_3 ? _GEN_9591 : _GEN_9431; // @[executor.scala 308:60]
  wire [7:0] _GEN_9752 = 8'h4 < length_3 ? _GEN_9592 : _GEN_9432; // @[executor.scala 308:60]
  wire [7:0] _GEN_9753 = 8'h4 < length_3 ? _GEN_9593 : _GEN_9433; // @[executor.scala 308:60]
  wire [7:0] _GEN_9754 = 8'h4 < length_3 ? _GEN_9594 : _GEN_9434; // @[executor.scala 308:60]
  wire [7:0] _GEN_9755 = 8'h4 < length_3 ? _GEN_9595 : _GEN_9435; // @[executor.scala 308:60]
  wire [7:0] _GEN_9756 = 8'h4 < length_3 ? _GEN_9596 : _GEN_9436; // @[executor.scala 308:60]
  wire [7:0] _GEN_9757 = 8'h4 < length_3 ? _GEN_9597 : _GEN_9437; // @[executor.scala 308:60]
  wire [7:0] _GEN_9758 = 8'h4 < length_3 ? _GEN_9598 : _GEN_9438; // @[executor.scala 308:60]
  wire [7:0] _GEN_9759 = 8'h4 < length_3 ? _GEN_9599 : _GEN_9439; // @[executor.scala 308:60]
  wire [7:0] _GEN_9760 = 8'h4 < length_3 ? _GEN_9600 : _GEN_9440; // @[executor.scala 308:60]
  wire [7:0] _GEN_9761 = 8'h4 < length_3 ? _GEN_9601 : _GEN_9441; // @[executor.scala 308:60]
  wire [7:0] _GEN_9762 = 8'h4 < length_3 ? _GEN_9602 : _GEN_9442; // @[executor.scala 308:60]
  wire [7:0] _GEN_9763 = 8'h4 < length_3 ? _GEN_9603 : _GEN_9443; // @[executor.scala 308:60]
  wire [7:0] _GEN_9764 = 8'h4 < length_3 ? _GEN_9604 : _GEN_9444; // @[executor.scala 308:60]
  wire [7:0] _GEN_9765 = 8'h4 < length_3 ? _GEN_9605 : _GEN_9445; // @[executor.scala 308:60]
  wire [7:0] field_byte_29 = field_3[23:16]; // @[executor.scala 305:57]
  wire [7:0] total_offset_29 = offset_3 + 8'h5; // @[executor.scala 307:57]
  wire [7:0] _GEN_9766 = 8'h0 == total_offset_29 ? field_byte_29 : _GEN_9606; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9767 = 8'h1 == total_offset_29 ? field_byte_29 : _GEN_9607; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9768 = 8'h2 == total_offset_29 ? field_byte_29 : _GEN_9608; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9769 = 8'h3 == total_offset_29 ? field_byte_29 : _GEN_9609; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9770 = 8'h4 == total_offset_29 ? field_byte_29 : _GEN_9610; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9771 = 8'h5 == total_offset_29 ? field_byte_29 : _GEN_9611; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9772 = 8'h6 == total_offset_29 ? field_byte_29 : _GEN_9612; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9773 = 8'h7 == total_offset_29 ? field_byte_29 : _GEN_9613; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9774 = 8'h8 == total_offset_29 ? field_byte_29 : _GEN_9614; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9775 = 8'h9 == total_offset_29 ? field_byte_29 : _GEN_9615; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9776 = 8'ha == total_offset_29 ? field_byte_29 : _GEN_9616; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9777 = 8'hb == total_offset_29 ? field_byte_29 : _GEN_9617; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9778 = 8'hc == total_offset_29 ? field_byte_29 : _GEN_9618; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9779 = 8'hd == total_offset_29 ? field_byte_29 : _GEN_9619; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9780 = 8'he == total_offset_29 ? field_byte_29 : _GEN_9620; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9781 = 8'hf == total_offset_29 ? field_byte_29 : _GEN_9621; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9782 = 8'h10 == total_offset_29 ? field_byte_29 : _GEN_9622; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9783 = 8'h11 == total_offset_29 ? field_byte_29 : _GEN_9623; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9784 = 8'h12 == total_offset_29 ? field_byte_29 : _GEN_9624; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9785 = 8'h13 == total_offset_29 ? field_byte_29 : _GEN_9625; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9786 = 8'h14 == total_offset_29 ? field_byte_29 : _GEN_9626; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9787 = 8'h15 == total_offset_29 ? field_byte_29 : _GEN_9627; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9788 = 8'h16 == total_offset_29 ? field_byte_29 : _GEN_9628; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9789 = 8'h17 == total_offset_29 ? field_byte_29 : _GEN_9629; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9790 = 8'h18 == total_offset_29 ? field_byte_29 : _GEN_9630; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9791 = 8'h19 == total_offset_29 ? field_byte_29 : _GEN_9631; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9792 = 8'h1a == total_offset_29 ? field_byte_29 : _GEN_9632; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9793 = 8'h1b == total_offset_29 ? field_byte_29 : _GEN_9633; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9794 = 8'h1c == total_offset_29 ? field_byte_29 : _GEN_9634; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9795 = 8'h1d == total_offset_29 ? field_byte_29 : _GEN_9635; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9796 = 8'h1e == total_offset_29 ? field_byte_29 : _GEN_9636; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9797 = 8'h1f == total_offset_29 ? field_byte_29 : _GEN_9637; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9798 = 8'h20 == total_offset_29 ? field_byte_29 : _GEN_9638; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9799 = 8'h21 == total_offset_29 ? field_byte_29 : _GEN_9639; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9800 = 8'h22 == total_offset_29 ? field_byte_29 : _GEN_9640; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9801 = 8'h23 == total_offset_29 ? field_byte_29 : _GEN_9641; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9802 = 8'h24 == total_offset_29 ? field_byte_29 : _GEN_9642; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9803 = 8'h25 == total_offset_29 ? field_byte_29 : _GEN_9643; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9804 = 8'h26 == total_offset_29 ? field_byte_29 : _GEN_9644; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9805 = 8'h27 == total_offset_29 ? field_byte_29 : _GEN_9645; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9806 = 8'h28 == total_offset_29 ? field_byte_29 : _GEN_9646; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9807 = 8'h29 == total_offset_29 ? field_byte_29 : _GEN_9647; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9808 = 8'h2a == total_offset_29 ? field_byte_29 : _GEN_9648; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9809 = 8'h2b == total_offset_29 ? field_byte_29 : _GEN_9649; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9810 = 8'h2c == total_offset_29 ? field_byte_29 : _GEN_9650; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9811 = 8'h2d == total_offset_29 ? field_byte_29 : _GEN_9651; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9812 = 8'h2e == total_offset_29 ? field_byte_29 : _GEN_9652; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9813 = 8'h2f == total_offset_29 ? field_byte_29 : _GEN_9653; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9814 = 8'h30 == total_offset_29 ? field_byte_29 : _GEN_9654; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9815 = 8'h31 == total_offset_29 ? field_byte_29 : _GEN_9655; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9816 = 8'h32 == total_offset_29 ? field_byte_29 : _GEN_9656; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9817 = 8'h33 == total_offset_29 ? field_byte_29 : _GEN_9657; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9818 = 8'h34 == total_offset_29 ? field_byte_29 : _GEN_9658; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9819 = 8'h35 == total_offset_29 ? field_byte_29 : _GEN_9659; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9820 = 8'h36 == total_offset_29 ? field_byte_29 : _GEN_9660; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9821 = 8'h37 == total_offset_29 ? field_byte_29 : _GEN_9661; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9822 = 8'h38 == total_offset_29 ? field_byte_29 : _GEN_9662; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9823 = 8'h39 == total_offset_29 ? field_byte_29 : _GEN_9663; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9824 = 8'h3a == total_offset_29 ? field_byte_29 : _GEN_9664; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9825 = 8'h3b == total_offset_29 ? field_byte_29 : _GEN_9665; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9826 = 8'h3c == total_offset_29 ? field_byte_29 : _GEN_9666; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9827 = 8'h3d == total_offset_29 ? field_byte_29 : _GEN_9667; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9828 = 8'h3e == total_offset_29 ? field_byte_29 : _GEN_9668; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9829 = 8'h3f == total_offset_29 ? field_byte_29 : _GEN_9669; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9830 = 8'h40 == total_offset_29 ? field_byte_29 : _GEN_9670; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9831 = 8'h41 == total_offset_29 ? field_byte_29 : _GEN_9671; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9832 = 8'h42 == total_offset_29 ? field_byte_29 : _GEN_9672; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9833 = 8'h43 == total_offset_29 ? field_byte_29 : _GEN_9673; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9834 = 8'h44 == total_offset_29 ? field_byte_29 : _GEN_9674; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9835 = 8'h45 == total_offset_29 ? field_byte_29 : _GEN_9675; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9836 = 8'h46 == total_offset_29 ? field_byte_29 : _GEN_9676; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9837 = 8'h47 == total_offset_29 ? field_byte_29 : _GEN_9677; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9838 = 8'h48 == total_offset_29 ? field_byte_29 : _GEN_9678; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9839 = 8'h49 == total_offset_29 ? field_byte_29 : _GEN_9679; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9840 = 8'h4a == total_offset_29 ? field_byte_29 : _GEN_9680; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9841 = 8'h4b == total_offset_29 ? field_byte_29 : _GEN_9681; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9842 = 8'h4c == total_offset_29 ? field_byte_29 : _GEN_9682; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9843 = 8'h4d == total_offset_29 ? field_byte_29 : _GEN_9683; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9844 = 8'h4e == total_offset_29 ? field_byte_29 : _GEN_9684; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9845 = 8'h4f == total_offset_29 ? field_byte_29 : _GEN_9685; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9846 = 8'h50 == total_offset_29 ? field_byte_29 : _GEN_9686; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9847 = 8'h51 == total_offset_29 ? field_byte_29 : _GEN_9687; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9848 = 8'h52 == total_offset_29 ? field_byte_29 : _GEN_9688; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9849 = 8'h53 == total_offset_29 ? field_byte_29 : _GEN_9689; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9850 = 8'h54 == total_offset_29 ? field_byte_29 : _GEN_9690; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9851 = 8'h55 == total_offset_29 ? field_byte_29 : _GEN_9691; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9852 = 8'h56 == total_offset_29 ? field_byte_29 : _GEN_9692; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9853 = 8'h57 == total_offset_29 ? field_byte_29 : _GEN_9693; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9854 = 8'h58 == total_offset_29 ? field_byte_29 : _GEN_9694; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9855 = 8'h59 == total_offset_29 ? field_byte_29 : _GEN_9695; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9856 = 8'h5a == total_offset_29 ? field_byte_29 : _GEN_9696; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9857 = 8'h5b == total_offset_29 ? field_byte_29 : _GEN_9697; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9858 = 8'h5c == total_offset_29 ? field_byte_29 : _GEN_9698; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9859 = 8'h5d == total_offset_29 ? field_byte_29 : _GEN_9699; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9860 = 8'h5e == total_offset_29 ? field_byte_29 : _GEN_9700; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9861 = 8'h5f == total_offset_29 ? field_byte_29 : _GEN_9701; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9862 = 8'h60 == total_offset_29 ? field_byte_29 : _GEN_9702; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9863 = 8'h61 == total_offset_29 ? field_byte_29 : _GEN_9703; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9864 = 8'h62 == total_offset_29 ? field_byte_29 : _GEN_9704; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9865 = 8'h63 == total_offset_29 ? field_byte_29 : _GEN_9705; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9866 = 8'h64 == total_offset_29 ? field_byte_29 : _GEN_9706; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9867 = 8'h65 == total_offset_29 ? field_byte_29 : _GEN_9707; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9868 = 8'h66 == total_offset_29 ? field_byte_29 : _GEN_9708; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9869 = 8'h67 == total_offset_29 ? field_byte_29 : _GEN_9709; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9870 = 8'h68 == total_offset_29 ? field_byte_29 : _GEN_9710; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9871 = 8'h69 == total_offset_29 ? field_byte_29 : _GEN_9711; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9872 = 8'h6a == total_offset_29 ? field_byte_29 : _GEN_9712; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9873 = 8'h6b == total_offset_29 ? field_byte_29 : _GEN_9713; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9874 = 8'h6c == total_offset_29 ? field_byte_29 : _GEN_9714; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9875 = 8'h6d == total_offset_29 ? field_byte_29 : _GEN_9715; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9876 = 8'h6e == total_offset_29 ? field_byte_29 : _GEN_9716; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9877 = 8'h6f == total_offset_29 ? field_byte_29 : _GEN_9717; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9878 = 8'h70 == total_offset_29 ? field_byte_29 : _GEN_9718; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9879 = 8'h71 == total_offset_29 ? field_byte_29 : _GEN_9719; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9880 = 8'h72 == total_offset_29 ? field_byte_29 : _GEN_9720; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9881 = 8'h73 == total_offset_29 ? field_byte_29 : _GEN_9721; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9882 = 8'h74 == total_offset_29 ? field_byte_29 : _GEN_9722; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9883 = 8'h75 == total_offset_29 ? field_byte_29 : _GEN_9723; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9884 = 8'h76 == total_offset_29 ? field_byte_29 : _GEN_9724; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9885 = 8'h77 == total_offset_29 ? field_byte_29 : _GEN_9725; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9886 = 8'h78 == total_offset_29 ? field_byte_29 : _GEN_9726; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9887 = 8'h79 == total_offset_29 ? field_byte_29 : _GEN_9727; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9888 = 8'h7a == total_offset_29 ? field_byte_29 : _GEN_9728; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9889 = 8'h7b == total_offset_29 ? field_byte_29 : _GEN_9729; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9890 = 8'h7c == total_offset_29 ? field_byte_29 : _GEN_9730; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9891 = 8'h7d == total_offset_29 ? field_byte_29 : _GEN_9731; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9892 = 8'h7e == total_offset_29 ? field_byte_29 : _GEN_9732; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9893 = 8'h7f == total_offset_29 ? field_byte_29 : _GEN_9733; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9894 = 8'h80 == total_offset_29 ? field_byte_29 : _GEN_9734; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9895 = 8'h81 == total_offset_29 ? field_byte_29 : _GEN_9735; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9896 = 8'h82 == total_offset_29 ? field_byte_29 : _GEN_9736; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9897 = 8'h83 == total_offset_29 ? field_byte_29 : _GEN_9737; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9898 = 8'h84 == total_offset_29 ? field_byte_29 : _GEN_9738; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9899 = 8'h85 == total_offset_29 ? field_byte_29 : _GEN_9739; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9900 = 8'h86 == total_offset_29 ? field_byte_29 : _GEN_9740; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9901 = 8'h87 == total_offset_29 ? field_byte_29 : _GEN_9741; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9902 = 8'h88 == total_offset_29 ? field_byte_29 : _GEN_9742; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9903 = 8'h89 == total_offset_29 ? field_byte_29 : _GEN_9743; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9904 = 8'h8a == total_offset_29 ? field_byte_29 : _GEN_9744; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9905 = 8'h8b == total_offset_29 ? field_byte_29 : _GEN_9745; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9906 = 8'h8c == total_offset_29 ? field_byte_29 : _GEN_9746; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9907 = 8'h8d == total_offset_29 ? field_byte_29 : _GEN_9747; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9908 = 8'h8e == total_offset_29 ? field_byte_29 : _GEN_9748; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9909 = 8'h8f == total_offset_29 ? field_byte_29 : _GEN_9749; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9910 = 8'h90 == total_offset_29 ? field_byte_29 : _GEN_9750; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9911 = 8'h91 == total_offset_29 ? field_byte_29 : _GEN_9751; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9912 = 8'h92 == total_offset_29 ? field_byte_29 : _GEN_9752; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9913 = 8'h93 == total_offset_29 ? field_byte_29 : _GEN_9753; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9914 = 8'h94 == total_offset_29 ? field_byte_29 : _GEN_9754; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9915 = 8'h95 == total_offset_29 ? field_byte_29 : _GEN_9755; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9916 = 8'h96 == total_offset_29 ? field_byte_29 : _GEN_9756; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9917 = 8'h97 == total_offset_29 ? field_byte_29 : _GEN_9757; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9918 = 8'h98 == total_offset_29 ? field_byte_29 : _GEN_9758; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9919 = 8'h99 == total_offset_29 ? field_byte_29 : _GEN_9759; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9920 = 8'h9a == total_offset_29 ? field_byte_29 : _GEN_9760; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9921 = 8'h9b == total_offset_29 ? field_byte_29 : _GEN_9761; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9922 = 8'h9c == total_offset_29 ? field_byte_29 : _GEN_9762; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9923 = 8'h9d == total_offset_29 ? field_byte_29 : _GEN_9763; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9924 = 8'h9e == total_offset_29 ? field_byte_29 : _GEN_9764; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9925 = 8'h9f == total_offset_29 ? field_byte_29 : _GEN_9765; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_9926 = 8'h5 < length_3 ? _GEN_9766 : _GEN_9606; // @[executor.scala 308:60]
  wire [7:0] _GEN_9927 = 8'h5 < length_3 ? _GEN_9767 : _GEN_9607; // @[executor.scala 308:60]
  wire [7:0] _GEN_9928 = 8'h5 < length_3 ? _GEN_9768 : _GEN_9608; // @[executor.scala 308:60]
  wire [7:0] _GEN_9929 = 8'h5 < length_3 ? _GEN_9769 : _GEN_9609; // @[executor.scala 308:60]
  wire [7:0] _GEN_9930 = 8'h5 < length_3 ? _GEN_9770 : _GEN_9610; // @[executor.scala 308:60]
  wire [7:0] _GEN_9931 = 8'h5 < length_3 ? _GEN_9771 : _GEN_9611; // @[executor.scala 308:60]
  wire [7:0] _GEN_9932 = 8'h5 < length_3 ? _GEN_9772 : _GEN_9612; // @[executor.scala 308:60]
  wire [7:0] _GEN_9933 = 8'h5 < length_3 ? _GEN_9773 : _GEN_9613; // @[executor.scala 308:60]
  wire [7:0] _GEN_9934 = 8'h5 < length_3 ? _GEN_9774 : _GEN_9614; // @[executor.scala 308:60]
  wire [7:0] _GEN_9935 = 8'h5 < length_3 ? _GEN_9775 : _GEN_9615; // @[executor.scala 308:60]
  wire [7:0] _GEN_9936 = 8'h5 < length_3 ? _GEN_9776 : _GEN_9616; // @[executor.scala 308:60]
  wire [7:0] _GEN_9937 = 8'h5 < length_3 ? _GEN_9777 : _GEN_9617; // @[executor.scala 308:60]
  wire [7:0] _GEN_9938 = 8'h5 < length_3 ? _GEN_9778 : _GEN_9618; // @[executor.scala 308:60]
  wire [7:0] _GEN_9939 = 8'h5 < length_3 ? _GEN_9779 : _GEN_9619; // @[executor.scala 308:60]
  wire [7:0] _GEN_9940 = 8'h5 < length_3 ? _GEN_9780 : _GEN_9620; // @[executor.scala 308:60]
  wire [7:0] _GEN_9941 = 8'h5 < length_3 ? _GEN_9781 : _GEN_9621; // @[executor.scala 308:60]
  wire [7:0] _GEN_9942 = 8'h5 < length_3 ? _GEN_9782 : _GEN_9622; // @[executor.scala 308:60]
  wire [7:0] _GEN_9943 = 8'h5 < length_3 ? _GEN_9783 : _GEN_9623; // @[executor.scala 308:60]
  wire [7:0] _GEN_9944 = 8'h5 < length_3 ? _GEN_9784 : _GEN_9624; // @[executor.scala 308:60]
  wire [7:0] _GEN_9945 = 8'h5 < length_3 ? _GEN_9785 : _GEN_9625; // @[executor.scala 308:60]
  wire [7:0] _GEN_9946 = 8'h5 < length_3 ? _GEN_9786 : _GEN_9626; // @[executor.scala 308:60]
  wire [7:0] _GEN_9947 = 8'h5 < length_3 ? _GEN_9787 : _GEN_9627; // @[executor.scala 308:60]
  wire [7:0] _GEN_9948 = 8'h5 < length_3 ? _GEN_9788 : _GEN_9628; // @[executor.scala 308:60]
  wire [7:0] _GEN_9949 = 8'h5 < length_3 ? _GEN_9789 : _GEN_9629; // @[executor.scala 308:60]
  wire [7:0] _GEN_9950 = 8'h5 < length_3 ? _GEN_9790 : _GEN_9630; // @[executor.scala 308:60]
  wire [7:0] _GEN_9951 = 8'h5 < length_3 ? _GEN_9791 : _GEN_9631; // @[executor.scala 308:60]
  wire [7:0] _GEN_9952 = 8'h5 < length_3 ? _GEN_9792 : _GEN_9632; // @[executor.scala 308:60]
  wire [7:0] _GEN_9953 = 8'h5 < length_3 ? _GEN_9793 : _GEN_9633; // @[executor.scala 308:60]
  wire [7:0] _GEN_9954 = 8'h5 < length_3 ? _GEN_9794 : _GEN_9634; // @[executor.scala 308:60]
  wire [7:0] _GEN_9955 = 8'h5 < length_3 ? _GEN_9795 : _GEN_9635; // @[executor.scala 308:60]
  wire [7:0] _GEN_9956 = 8'h5 < length_3 ? _GEN_9796 : _GEN_9636; // @[executor.scala 308:60]
  wire [7:0] _GEN_9957 = 8'h5 < length_3 ? _GEN_9797 : _GEN_9637; // @[executor.scala 308:60]
  wire [7:0] _GEN_9958 = 8'h5 < length_3 ? _GEN_9798 : _GEN_9638; // @[executor.scala 308:60]
  wire [7:0] _GEN_9959 = 8'h5 < length_3 ? _GEN_9799 : _GEN_9639; // @[executor.scala 308:60]
  wire [7:0] _GEN_9960 = 8'h5 < length_3 ? _GEN_9800 : _GEN_9640; // @[executor.scala 308:60]
  wire [7:0] _GEN_9961 = 8'h5 < length_3 ? _GEN_9801 : _GEN_9641; // @[executor.scala 308:60]
  wire [7:0] _GEN_9962 = 8'h5 < length_3 ? _GEN_9802 : _GEN_9642; // @[executor.scala 308:60]
  wire [7:0] _GEN_9963 = 8'h5 < length_3 ? _GEN_9803 : _GEN_9643; // @[executor.scala 308:60]
  wire [7:0] _GEN_9964 = 8'h5 < length_3 ? _GEN_9804 : _GEN_9644; // @[executor.scala 308:60]
  wire [7:0] _GEN_9965 = 8'h5 < length_3 ? _GEN_9805 : _GEN_9645; // @[executor.scala 308:60]
  wire [7:0] _GEN_9966 = 8'h5 < length_3 ? _GEN_9806 : _GEN_9646; // @[executor.scala 308:60]
  wire [7:0] _GEN_9967 = 8'h5 < length_3 ? _GEN_9807 : _GEN_9647; // @[executor.scala 308:60]
  wire [7:0] _GEN_9968 = 8'h5 < length_3 ? _GEN_9808 : _GEN_9648; // @[executor.scala 308:60]
  wire [7:0] _GEN_9969 = 8'h5 < length_3 ? _GEN_9809 : _GEN_9649; // @[executor.scala 308:60]
  wire [7:0] _GEN_9970 = 8'h5 < length_3 ? _GEN_9810 : _GEN_9650; // @[executor.scala 308:60]
  wire [7:0] _GEN_9971 = 8'h5 < length_3 ? _GEN_9811 : _GEN_9651; // @[executor.scala 308:60]
  wire [7:0] _GEN_9972 = 8'h5 < length_3 ? _GEN_9812 : _GEN_9652; // @[executor.scala 308:60]
  wire [7:0] _GEN_9973 = 8'h5 < length_3 ? _GEN_9813 : _GEN_9653; // @[executor.scala 308:60]
  wire [7:0] _GEN_9974 = 8'h5 < length_3 ? _GEN_9814 : _GEN_9654; // @[executor.scala 308:60]
  wire [7:0] _GEN_9975 = 8'h5 < length_3 ? _GEN_9815 : _GEN_9655; // @[executor.scala 308:60]
  wire [7:0] _GEN_9976 = 8'h5 < length_3 ? _GEN_9816 : _GEN_9656; // @[executor.scala 308:60]
  wire [7:0] _GEN_9977 = 8'h5 < length_3 ? _GEN_9817 : _GEN_9657; // @[executor.scala 308:60]
  wire [7:0] _GEN_9978 = 8'h5 < length_3 ? _GEN_9818 : _GEN_9658; // @[executor.scala 308:60]
  wire [7:0] _GEN_9979 = 8'h5 < length_3 ? _GEN_9819 : _GEN_9659; // @[executor.scala 308:60]
  wire [7:0] _GEN_9980 = 8'h5 < length_3 ? _GEN_9820 : _GEN_9660; // @[executor.scala 308:60]
  wire [7:0] _GEN_9981 = 8'h5 < length_3 ? _GEN_9821 : _GEN_9661; // @[executor.scala 308:60]
  wire [7:0] _GEN_9982 = 8'h5 < length_3 ? _GEN_9822 : _GEN_9662; // @[executor.scala 308:60]
  wire [7:0] _GEN_9983 = 8'h5 < length_3 ? _GEN_9823 : _GEN_9663; // @[executor.scala 308:60]
  wire [7:0] _GEN_9984 = 8'h5 < length_3 ? _GEN_9824 : _GEN_9664; // @[executor.scala 308:60]
  wire [7:0] _GEN_9985 = 8'h5 < length_3 ? _GEN_9825 : _GEN_9665; // @[executor.scala 308:60]
  wire [7:0] _GEN_9986 = 8'h5 < length_3 ? _GEN_9826 : _GEN_9666; // @[executor.scala 308:60]
  wire [7:0] _GEN_9987 = 8'h5 < length_3 ? _GEN_9827 : _GEN_9667; // @[executor.scala 308:60]
  wire [7:0] _GEN_9988 = 8'h5 < length_3 ? _GEN_9828 : _GEN_9668; // @[executor.scala 308:60]
  wire [7:0] _GEN_9989 = 8'h5 < length_3 ? _GEN_9829 : _GEN_9669; // @[executor.scala 308:60]
  wire [7:0] _GEN_9990 = 8'h5 < length_3 ? _GEN_9830 : _GEN_9670; // @[executor.scala 308:60]
  wire [7:0] _GEN_9991 = 8'h5 < length_3 ? _GEN_9831 : _GEN_9671; // @[executor.scala 308:60]
  wire [7:0] _GEN_9992 = 8'h5 < length_3 ? _GEN_9832 : _GEN_9672; // @[executor.scala 308:60]
  wire [7:0] _GEN_9993 = 8'h5 < length_3 ? _GEN_9833 : _GEN_9673; // @[executor.scala 308:60]
  wire [7:0] _GEN_9994 = 8'h5 < length_3 ? _GEN_9834 : _GEN_9674; // @[executor.scala 308:60]
  wire [7:0] _GEN_9995 = 8'h5 < length_3 ? _GEN_9835 : _GEN_9675; // @[executor.scala 308:60]
  wire [7:0] _GEN_9996 = 8'h5 < length_3 ? _GEN_9836 : _GEN_9676; // @[executor.scala 308:60]
  wire [7:0] _GEN_9997 = 8'h5 < length_3 ? _GEN_9837 : _GEN_9677; // @[executor.scala 308:60]
  wire [7:0] _GEN_9998 = 8'h5 < length_3 ? _GEN_9838 : _GEN_9678; // @[executor.scala 308:60]
  wire [7:0] _GEN_9999 = 8'h5 < length_3 ? _GEN_9839 : _GEN_9679; // @[executor.scala 308:60]
  wire [7:0] _GEN_10000 = 8'h5 < length_3 ? _GEN_9840 : _GEN_9680; // @[executor.scala 308:60]
  wire [7:0] _GEN_10001 = 8'h5 < length_3 ? _GEN_9841 : _GEN_9681; // @[executor.scala 308:60]
  wire [7:0] _GEN_10002 = 8'h5 < length_3 ? _GEN_9842 : _GEN_9682; // @[executor.scala 308:60]
  wire [7:0] _GEN_10003 = 8'h5 < length_3 ? _GEN_9843 : _GEN_9683; // @[executor.scala 308:60]
  wire [7:0] _GEN_10004 = 8'h5 < length_3 ? _GEN_9844 : _GEN_9684; // @[executor.scala 308:60]
  wire [7:0] _GEN_10005 = 8'h5 < length_3 ? _GEN_9845 : _GEN_9685; // @[executor.scala 308:60]
  wire [7:0] _GEN_10006 = 8'h5 < length_3 ? _GEN_9846 : _GEN_9686; // @[executor.scala 308:60]
  wire [7:0] _GEN_10007 = 8'h5 < length_3 ? _GEN_9847 : _GEN_9687; // @[executor.scala 308:60]
  wire [7:0] _GEN_10008 = 8'h5 < length_3 ? _GEN_9848 : _GEN_9688; // @[executor.scala 308:60]
  wire [7:0] _GEN_10009 = 8'h5 < length_3 ? _GEN_9849 : _GEN_9689; // @[executor.scala 308:60]
  wire [7:0] _GEN_10010 = 8'h5 < length_3 ? _GEN_9850 : _GEN_9690; // @[executor.scala 308:60]
  wire [7:0] _GEN_10011 = 8'h5 < length_3 ? _GEN_9851 : _GEN_9691; // @[executor.scala 308:60]
  wire [7:0] _GEN_10012 = 8'h5 < length_3 ? _GEN_9852 : _GEN_9692; // @[executor.scala 308:60]
  wire [7:0] _GEN_10013 = 8'h5 < length_3 ? _GEN_9853 : _GEN_9693; // @[executor.scala 308:60]
  wire [7:0] _GEN_10014 = 8'h5 < length_3 ? _GEN_9854 : _GEN_9694; // @[executor.scala 308:60]
  wire [7:0] _GEN_10015 = 8'h5 < length_3 ? _GEN_9855 : _GEN_9695; // @[executor.scala 308:60]
  wire [7:0] _GEN_10016 = 8'h5 < length_3 ? _GEN_9856 : _GEN_9696; // @[executor.scala 308:60]
  wire [7:0] _GEN_10017 = 8'h5 < length_3 ? _GEN_9857 : _GEN_9697; // @[executor.scala 308:60]
  wire [7:0] _GEN_10018 = 8'h5 < length_3 ? _GEN_9858 : _GEN_9698; // @[executor.scala 308:60]
  wire [7:0] _GEN_10019 = 8'h5 < length_3 ? _GEN_9859 : _GEN_9699; // @[executor.scala 308:60]
  wire [7:0] _GEN_10020 = 8'h5 < length_3 ? _GEN_9860 : _GEN_9700; // @[executor.scala 308:60]
  wire [7:0] _GEN_10021 = 8'h5 < length_3 ? _GEN_9861 : _GEN_9701; // @[executor.scala 308:60]
  wire [7:0] _GEN_10022 = 8'h5 < length_3 ? _GEN_9862 : _GEN_9702; // @[executor.scala 308:60]
  wire [7:0] _GEN_10023 = 8'h5 < length_3 ? _GEN_9863 : _GEN_9703; // @[executor.scala 308:60]
  wire [7:0] _GEN_10024 = 8'h5 < length_3 ? _GEN_9864 : _GEN_9704; // @[executor.scala 308:60]
  wire [7:0] _GEN_10025 = 8'h5 < length_3 ? _GEN_9865 : _GEN_9705; // @[executor.scala 308:60]
  wire [7:0] _GEN_10026 = 8'h5 < length_3 ? _GEN_9866 : _GEN_9706; // @[executor.scala 308:60]
  wire [7:0] _GEN_10027 = 8'h5 < length_3 ? _GEN_9867 : _GEN_9707; // @[executor.scala 308:60]
  wire [7:0] _GEN_10028 = 8'h5 < length_3 ? _GEN_9868 : _GEN_9708; // @[executor.scala 308:60]
  wire [7:0] _GEN_10029 = 8'h5 < length_3 ? _GEN_9869 : _GEN_9709; // @[executor.scala 308:60]
  wire [7:0] _GEN_10030 = 8'h5 < length_3 ? _GEN_9870 : _GEN_9710; // @[executor.scala 308:60]
  wire [7:0] _GEN_10031 = 8'h5 < length_3 ? _GEN_9871 : _GEN_9711; // @[executor.scala 308:60]
  wire [7:0] _GEN_10032 = 8'h5 < length_3 ? _GEN_9872 : _GEN_9712; // @[executor.scala 308:60]
  wire [7:0] _GEN_10033 = 8'h5 < length_3 ? _GEN_9873 : _GEN_9713; // @[executor.scala 308:60]
  wire [7:0] _GEN_10034 = 8'h5 < length_3 ? _GEN_9874 : _GEN_9714; // @[executor.scala 308:60]
  wire [7:0] _GEN_10035 = 8'h5 < length_3 ? _GEN_9875 : _GEN_9715; // @[executor.scala 308:60]
  wire [7:0] _GEN_10036 = 8'h5 < length_3 ? _GEN_9876 : _GEN_9716; // @[executor.scala 308:60]
  wire [7:0] _GEN_10037 = 8'h5 < length_3 ? _GEN_9877 : _GEN_9717; // @[executor.scala 308:60]
  wire [7:0] _GEN_10038 = 8'h5 < length_3 ? _GEN_9878 : _GEN_9718; // @[executor.scala 308:60]
  wire [7:0] _GEN_10039 = 8'h5 < length_3 ? _GEN_9879 : _GEN_9719; // @[executor.scala 308:60]
  wire [7:0] _GEN_10040 = 8'h5 < length_3 ? _GEN_9880 : _GEN_9720; // @[executor.scala 308:60]
  wire [7:0] _GEN_10041 = 8'h5 < length_3 ? _GEN_9881 : _GEN_9721; // @[executor.scala 308:60]
  wire [7:0] _GEN_10042 = 8'h5 < length_3 ? _GEN_9882 : _GEN_9722; // @[executor.scala 308:60]
  wire [7:0] _GEN_10043 = 8'h5 < length_3 ? _GEN_9883 : _GEN_9723; // @[executor.scala 308:60]
  wire [7:0] _GEN_10044 = 8'h5 < length_3 ? _GEN_9884 : _GEN_9724; // @[executor.scala 308:60]
  wire [7:0] _GEN_10045 = 8'h5 < length_3 ? _GEN_9885 : _GEN_9725; // @[executor.scala 308:60]
  wire [7:0] _GEN_10046 = 8'h5 < length_3 ? _GEN_9886 : _GEN_9726; // @[executor.scala 308:60]
  wire [7:0] _GEN_10047 = 8'h5 < length_3 ? _GEN_9887 : _GEN_9727; // @[executor.scala 308:60]
  wire [7:0] _GEN_10048 = 8'h5 < length_3 ? _GEN_9888 : _GEN_9728; // @[executor.scala 308:60]
  wire [7:0] _GEN_10049 = 8'h5 < length_3 ? _GEN_9889 : _GEN_9729; // @[executor.scala 308:60]
  wire [7:0] _GEN_10050 = 8'h5 < length_3 ? _GEN_9890 : _GEN_9730; // @[executor.scala 308:60]
  wire [7:0] _GEN_10051 = 8'h5 < length_3 ? _GEN_9891 : _GEN_9731; // @[executor.scala 308:60]
  wire [7:0] _GEN_10052 = 8'h5 < length_3 ? _GEN_9892 : _GEN_9732; // @[executor.scala 308:60]
  wire [7:0] _GEN_10053 = 8'h5 < length_3 ? _GEN_9893 : _GEN_9733; // @[executor.scala 308:60]
  wire [7:0] _GEN_10054 = 8'h5 < length_3 ? _GEN_9894 : _GEN_9734; // @[executor.scala 308:60]
  wire [7:0] _GEN_10055 = 8'h5 < length_3 ? _GEN_9895 : _GEN_9735; // @[executor.scala 308:60]
  wire [7:0] _GEN_10056 = 8'h5 < length_3 ? _GEN_9896 : _GEN_9736; // @[executor.scala 308:60]
  wire [7:0] _GEN_10057 = 8'h5 < length_3 ? _GEN_9897 : _GEN_9737; // @[executor.scala 308:60]
  wire [7:0] _GEN_10058 = 8'h5 < length_3 ? _GEN_9898 : _GEN_9738; // @[executor.scala 308:60]
  wire [7:0] _GEN_10059 = 8'h5 < length_3 ? _GEN_9899 : _GEN_9739; // @[executor.scala 308:60]
  wire [7:0] _GEN_10060 = 8'h5 < length_3 ? _GEN_9900 : _GEN_9740; // @[executor.scala 308:60]
  wire [7:0] _GEN_10061 = 8'h5 < length_3 ? _GEN_9901 : _GEN_9741; // @[executor.scala 308:60]
  wire [7:0] _GEN_10062 = 8'h5 < length_3 ? _GEN_9902 : _GEN_9742; // @[executor.scala 308:60]
  wire [7:0] _GEN_10063 = 8'h5 < length_3 ? _GEN_9903 : _GEN_9743; // @[executor.scala 308:60]
  wire [7:0] _GEN_10064 = 8'h5 < length_3 ? _GEN_9904 : _GEN_9744; // @[executor.scala 308:60]
  wire [7:0] _GEN_10065 = 8'h5 < length_3 ? _GEN_9905 : _GEN_9745; // @[executor.scala 308:60]
  wire [7:0] _GEN_10066 = 8'h5 < length_3 ? _GEN_9906 : _GEN_9746; // @[executor.scala 308:60]
  wire [7:0] _GEN_10067 = 8'h5 < length_3 ? _GEN_9907 : _GEN_9747; // @[executor.scala 308:60]
  wire [7:0] _GEN_10068 = 8'h5 < length_3 ? _GEN_9908 : _GEN_9748; // @[executor.scala 308:60]
  wire [7:0] _GEN_10069 = 8'h5 < length_3 ? _GEN_9909 : _GEN_9749; // @[executor.scala 308:60]
  wire [7:0] _GEN_10070 = 8'h5 < length_3 ? _GEN_9910 : _GEN_9750; // @[executor.scala 308:60]
  wire [7:0] _GEN_10071 = 8'h5 < length_3 ? _GEN_9911 : _GEN_9751; // @[executor.scala 308:60]
  wire [7:0] _GEN_10072 = 8'h5 < length_3 ? _GEN_9912 : _GEN_9752; // @[executor.scala 308:60]
  wire [7:0] _GEN_10073 = 8'h5 < length_3 ? _GEN_9913 : _GEN_9753; // @[executor.scala 308:60]
  wire [7:0] _GEN_10074 = 8'h5 < length_3 ? _GEN_9914 : _GEN_9754; // @[executor.scala 308:60]
  wire [7:0] _GEN_10075 = 8'h5 < length_3 ? _GEN_9915 : _GEN_9755; // @[executor.scala 308:60]
  wire [7:0] _GEN_10076 = 8'h5 < length_3 ? _GEN_9916 : _GEN_9756; // @[executor.scala 308:60]
  wire [7:0] _GEN_10077 = 8'h5 < length_3 ? _GEN_9917 : _GEN_9757; // @[executor.scala 308:60]
  wire [7:0] _GEN_10078 = 8'h5 < length_3 ? _GEN_9918 : _GEN_9758; // @[executor.scala 308:60]
  wire [7:0] _GEN_10079 = 8'h5 < length_3 ? _GEN_9919 : _GEN_9759; // @[executor.scala 308:60]
  wire [7:0] _GEN_10080 = 8'h5 < length_3 ? _GEN_9920 : _GEN_9760; // @[executor.scala 308:60]
  wire [7:0] _GEN_10081 = 8'h5 < length_3 ? _GEN_9921 : _GEN_9761; // @[executor.scala 308:60]
  wire [7:0] _GEN_10082 = 8'h5 < length_3 ? _GEN_9922 : _GEN_9762; // @[executor.scala 308:60]
  wire [7:0] _GEN_10083 = 8'h5 < length_3 ? _GEN_9923 : _GEN_9763; // @[executor.scala 308:60]
  wire [7:0] _GEN_10084 = 8'h5 < length_3 ? _GEN_9924 : _GEN_9764; // @[executor.scala 308:60]
  wire [7:0] _GEN_10085 = 8'h5 < length_3 ? _GEN_9925 : _GEN_9765; // @[executor.scala 308:60]
  wire [7:0] field_byte_30 = field_3[15:8]; // @[executor.scala 305:57]
  wire [7:0] total_offset_30 = offset_3 + 8'h6; // @[executor.scala 307:57]
  wire [7:0] _GEN_10086 = 8'h0 == total_offset_30 ? field_byte_30 : _GEN_9926; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10087 = 8'h1 == total_offset_30 ? field_byte_30 : _GEN_9927; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10088 = 8'h2 == total_offset_30 ? field_byte_30 : _GEN_9928; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10089 = 8'h3 == total_offset_30 ? field_byte_30 : _GEN_9929; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10090 = 8'h4 == total_offset_30 ? field_byte_30 : _GEN_9930; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10091 = 8'h5 == total_offset_30 ? field_byte_30 : _GEN_9931; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10092 = 8'h6 == total_offset_30 ? field_byte_30 : _GEN_9932; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10093 = 8'h7 == total_offset_30 ? field_byte_30 : _GEN_9933; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10094 = 8'h8 == total_offset_30 ? field_byte_30 : _GEN_9934; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10095 = 8'h9 == total_offset_30 ? field_byte_30 : _GEN_9935; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10096 = 8'ha == total_offset_30 ? field_byte_30 : _GEN_9936; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10097 = 8'hb == total_offset_30 ? field_byte_30 : _GEN_9937; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10098 = 8'hc == total_offset_30 ? field_byte_30 : _GEN_9938; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10099 = 8'hd == total_offset_30 ? field_byte_30 : _GEN_9939; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10100 = 8'he == total_offset_30 ? field_byte_30 : _GEN_9940; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10101 = 8'hf == total_offset_30 ? field_byte_30 : _GEN_9941; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10102 = 8'h10 == total_offset_30 ? field_byte_30 : _GEN_9942; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10103 = 8'h11 == total_offset_30 ? field_byte_30 : _GEN_9943; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10104 = 8'h12 == total_offset_30 ? field_byte_30 : _GEN_9944; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10105 = 8'h13 == total_offset_30 ? field_byte_30 : _GEN_9945; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10106 = 8'h14 == total_offset_30 ? field_byte_30 : _GEN_9946; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10107 = 8'h15 == total_offset_30 ? field_byte_30 : _GEN_9947; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10108 = 8'h16 == total_offset_30 ? field_byte_30 : _GEN_9948; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10109 = 8'h17 == total_offset_30 ? field_byte_30 : _GEN_9949; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10110 = 8'h18 == total_offset_30 ? field_byte_30 : _GEN_9950; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10111 = 8'h19 == total_offset_30 ? field_byte_30 : _GEN_9951; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10112 = 8'h1a == total_offset_30 ? field_byte_30 : _GEN_9952; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10113 = 8'h1b == total_offset_30 ? field_byte_30 : _GEN_9953; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10114 = 8'h1c == total_offset_30 ? field_byte_30 : _GEN_9954; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10115 = 8'h1d == total_offset_30 ? field_byte_30 : _GEN_9955; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10116 = 8'h1e == total_offset_30 ? field_byte_30 : _GEN_9956; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10117 = 8'h1f == total_offset_30 ? field_byte_30 : _GEN_9957; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10118 = 8'h20 == total_offset_30 ? field_byte_30 : _GEN_9958; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10119 = 8'h21 == total_offset_30 ? field_byte_30 : _GEN_9959; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10120 = 8'h22 == total_offset_30 ? field_byte_30 : _GEN_9960; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10121 = 8'h23 == total_offset_30 ? field_byte_30 : _GEN_9961; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10122 = 8'h24 == total_offset_30 ? field_byte_30 : _GEN_9962; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10123 = 8'h25 == total_offset_30 ? field_byte_30 : _GEN_9963; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10124 = 8'h26 == total_offset_30 ? field_byte_30 : _GEN_9964; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10125 = 8'h27 == total_offset_30 ? field_byte_30 : _GEN_9965; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10126 = 8'h28 == total_offset_30 ? field_byte_30 : _GEN_9966; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10127 = 8'h29 == total_offset_30 ? field_byte_30 : _GEN_9967; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10128 = 8'h2a == total_offset_30 ? field_byte_30 : _GEN_9968; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10129 = 8'h2b == total_offset_30 ? field_byte_30 : _GEN_9969; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10130 = 8'h2c == total_offset_30 ? field_byte_30 : _GEN_9970; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10131 = 8'h2d == total_offset_30 ? field_byte_30 : _GEN_9971; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10132 = 8'h2e == total_offset_30 ? field_byte_30 : _GEN_9972; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10133 = 8'h2f == total_offset_30 ? field_byte_30 : _GEN_9973; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10134 = 8'h30 == total_offset_30 ? field_byte_30 : _GEN_9974; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10135 = 8'h31 == total_offset_30 ? field_byte_30 : _GEN_9975; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10136 = 8'h32 == total_offset_30 ? field_byte_30 : _GEN_9976; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10137 = 8'h33 == total_offset_30 ? field_byte_30 : _GEN_9977; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10138 = 8'h34 == total_offset_30 ? field_byte_30 : _GEN_9978; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10139 = 8'h35 == total_offset_30 ? field_byte_30 : _GEN_9979; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10140 = 8'h36 == total_offset_30 ? field_byte_30 : _GEN_9980; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10141 = 8'h37 == total_offset_30 ? field_byte_30 : _GEN_9981; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10142 = 8'h38 == total_offset_30 ? field_byte_30 : _GEN_9982; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10143 = 8'h39 == total_offset_30 ? field_byte_30 : _GEN_9983; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10144 = 8'h3a == total_offset_30 ? field_byte_30 : _GEN_9984; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10145 = 8'h3b == total_offset_30 ? field_byte_30 : _GEN_9985; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10146 = 8'h3c == total_offset_30 ? field_byte_30 : _GEN_9986; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10147 = 8'h3d == total_offset_30 ? field_byte_30 : _GEN_9987; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10148 = 8'h3e == total_offset_30 ? field_byte_30 : _GEN_9988; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10149 = 8'h3f == total_offset_30 ? field_byte_30 : _GEN_9989; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10150 = 8'h40 == total_offset_30 ? field_byte_30 : _GEN_9990; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10151 = 8'h41 == total_offset_30 ? field_byte_30 : _GEN_9991; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10152 = 8'h42 == total_offset_30 ? field_byte_30 : _GEN_9992; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10153 = 8'h43 == total_offset_30 ? field_byte_30 : _GEN_9993; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10154 = 8'h44 == total_offset_30 ? field_byte_30 : _GEN_9994; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10155 = 8'h45 == total_offset_30 ? field_byte_30 : _GEN_9995; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10156 = 8'h46 == total_offset_30 ? field_byte_30 : _GEN_9996; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10157 = 8'h47 == total_offset_30 ? field_byte_30 : _GEN_9997; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10158 = 8'h48 == total_offset_30 ? field_byte_30 : _GEN_9998; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10159 = 8'h49 == total_offset_30 ? field_byte_30 : _GEN_9999; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10160 = 8'h4a == total_offset_30 ? field_byte_30 : _GEN_10000; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10161 = 8'h4b == total_offset_30 ? field_byte_30 : _GEN_10001; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10162 = 8'h4c == total_offset_30 ? field_byte_30 : _GEN_10002; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10163 = 8'h4d == total_offset_30 ? field_byte_30 : _GEN_10003; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10164 = 8'h4e == total_offset_30 ? field_byte_30 : _GEN_10004; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10165 = 8'h4f == total_offset_30 ? field_byte_30 : _GEN_10005; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10166 = 8'h50 == total_offset_30 ? field_byte_30 : _GEN_10006; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10167 = 8'h51 == total_offset_30 ? field_byte_30 : _GEN_10007; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10168 = 8'h52 == total_offset_30 ? field_byte_30 : _GEN_10008; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10169 = 8'h53 == total_offset_30 ? field_byte_30 : _GEN_10009; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10170 = 8'h54 == total_offset_30 ? field_byte_30 : _GEN_10010; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10171 = 8'h55 == total_offset_30 ? field_byte_30 : _GEN_10011; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10172 = 8'h56 == total_offset_30 ? field_byte_30 : _GEN_10012; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10173 = 8'h57 == total_offset_30 ? field_byte_30 : _GEN_10013; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10174 = 8'h58 == total_offset_30 ? field_byte_30 : _GEN_10014; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10175 = 8'h59 == total_offset_30 ? field_byte_30 : _GEN_10015; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10176 = 8'h5a == total_offset_30 ? field_byte_30 : _GEN_10016; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10177 = 8'h5b == total_offset_30 ? field_byte_30 : _GEN_10017; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10178 = 8'h5c == total_offset_30 ? field_byte_30 : _GEN_10018; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10179 = 8'h5d == total_offset_30 ? field_byte_30 : _GEN_10019; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10180 = 8'h5e == total_offset_30 ? field_byte_30 : _GEN_10020; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10181 = 8'h5f == total_offset_30 ? field_byte_30 : _GEN_10021; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10182 = 8'h60 == total_offset_30 ? field_byte_30 : _GEN_10022; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10183 = 8'h61 == total_offset_30 ? field_byte_30 : _GEN_10023; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10184 = 8'h62 == total_offset_30 ? field_byte_30 : _GEN_10024; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10185 = 8'h63 == total_offset_30 ? field_byte_30 : _GEN_10025; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10186 = 8'h64 == total_offset_30 ? field_byte_30 : _GEN_10026; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10187 = 8'h65 == total_offset_30 ? field_byte_30 : _GEN_10027; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10188 = 8'h66 == total_offset_30 ? field_byte_30 : _GEN_10028; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10189 = 8'h67 == total_offset_30 ? field_byte_30 : _GEN_10029; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10190 = 8'h68 == total_offset_30 ? field_byte_30 : _GEN_10030; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10191 = 8'h69 == total_offset_30 ? field_byte_30 : _GEN_10031; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10192 = 8'h6a == total_offset_30 ? field_byte_30 : _GEN_10032; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10193 = 8'h6b == total_offset_30 ? field_byte_30 : _GEN_10033; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10194 = 8'h6c == total_offset_30 ? field_byte_30 : _GEN_10034; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10195 = 8'h6d == total_offset_30 ? field_byte_30 : _GEN_10035; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10196 = 8'h6e == total_offset_30 ? field_byte_30 : _GEN_10036; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10197 = 8'h6f == total_offset_30 ? field_byte_30 : _GEN_10037; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10198 = 8'h70 == total_offset_30 ? field_byte_30 : _GEN_10038; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10199 = 8'h71 == total_offset_30 ? field_byte_30 : _GEN_10039; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10200 = 8'h72 == total_offset_30 ? field_byte_30 : _GEN_10040; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10201 = 8'h73 == total_offset_30 ? field_byte_30 : _GEN_10041; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10202 = 8'h74 == total_offset_30 ? field_byte_30 : _GEN_10042; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10203 = 8'h75 == total_offset_30 ? field_byte_30 : _GEN_10043; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10204 = 8'h76 == total_offset_30 ? field_byte_30 : _GEN_10044; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10205 = 8'h77 == total_offset_30 ? field_byte_30 : _GEN_10045; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10206 = 8'h78 == total_offset_30 ? field_byte_30 : _GEN_10046; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10207 = 8'h79 == total_offset_30 ? field_byte_30 : _GEN_10047; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10208 = 8'h7a == total_offset_30 ? field_byte_30 : _GEN_10048; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10209 = 8'h7b == total_offset_30 ? field_byte_30 : _GEN_10049; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10210 = 8'h7c == total_offset_30 ? field_byte_30 : _GEN_10050; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10211 = 8'h7d == total_offset_30 ? field_byte_30 : _GEN_10051; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10212 = 8'h7e == total_offset_30 ? field_byte_30 : _GEN_10052; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10213 = 8'h7f == total_offset_30 ? field_byte_30 : _GEN_10053; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10214 = 8'h80 == total_offset_30 ? field_byte_30 : _GEN_10054; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10215 = 8'h81 == total_offset_30 ? field_byte_30 : _GEN_10055; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10216 = 8'h82 == total_offset_30 ? field_byte_30 : _GEN_10056; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10217 = 8'h83 == total_offset_30 ? field_byte_30 : _GEN_10057; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10218 = 8'h84 == total_offset_30 ? field_byte_30 : _GEN_10058; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10219 = 8'h85 == total_offset_30 ? field_byte_30 : _GEN_10059; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10220 = 8'h86 == total_offset_30 ? field_byte_30 : _GEN_10060; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10221 = 8'h87 == total_offset_30 ? field_byte_30 : _GEN_10061; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10222 = 8'h88 == total_offset_30 ? field_byte_30 : _GEN_10062; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10223 = 8'h89 == total_offset_30 ? field_byte_30 : _GEN_10063; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10224 = 8'h8a == total_offset_30 ? field_byte_30 : _GEN_10064; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10225 = 8'h8b == total_offset_30 ? field_byte_30 : _GEN_10065; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10226 = 8'h8c == total_offset_30 ? field_byte_30 : _GEN_10066; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10227 = 8'h8d == total_offset_30 ? field_byte_30 : _GEN_10067; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10228 = 8'h8e == total_offset_30 ? field_byte_30 : _GEN_10068; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10229 = 8'h8f == total_offset_30 ? field_byte_30 : _GEN_10069; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10230 = 8'h90 == total_offset_30 ? field_byte_30 : _GEN_10070; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10231 = 8'h91 == total_offset_30 ? field_byte_30 : _GEN_10071; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10232 = 8'h92 == total_offset_30 ? field_byte_30 : _GEN_10072; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10233 = 8'h93 == total_offset_30 ? field_byte_30 : _GEN_10073; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10234 = 8'h94 == total_offset_30 ? field_byte_30 : _GEN_10074; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10235 = 8'h95 == total_offset_30 ? field_byte_30 : _GEN_10075; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10236 = 8'h96 == total_offset_30 ? field_byte_30 : _GEN_10076; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10237 = 8'h97 == total_offset_30 ? field_byte_30 : _GEN_10077; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10238 = 8'h98 == total_offset_30 ? field_byte_30 : _GEN_10078; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10239 = 8'h99 == total_offset_30 ? field_byte_30 : _GEN_10079; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10240 = 8'h9a == total_offset_30 ? field_byte_30 : _GEN_10080; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10241 = 8'h9b == total_offset_30 ? field_byte_30 : _GEN_10081; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10242 = 8'h9c == total_offset_30 ? field_byte_30 : _GEN_10082; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10243 = 8'h9d == total_offset_30 ? field_byte_30 : _GEN_10083; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10244 = 8'h9e == total_offset_30 ? field_byte_30 : _GEN_10084; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10245 = 8'h9f == total_offset_30 ? field_byte_30 : _GEN_10085; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10246 = 8'h6 < length_3 ? _GEN_10086 : _GEN_9926; // @[executor.scala 308:60]
  wire [7:0] _GEN_10247 = 8'h6 < length_3 ? _GEN_10087 : _GEN_9927; // @[executor.scala 308:60]
  wire [7:0] _GEN_10248 = 8'h6 < length_3 ? _GEN_10088 : _GEN_9928; // @[executor.scala 308:60]
  wire [7:0] _GEN_10249 = 8'h6 < length_3 ? _GEN_10089 : _GEN_9929; // @[executor.scala 308:60]
  wire [7:0] _GEN_10250 = 8'h6 < length_3 ? _GEN_10090 : _GEN_9930; // @[executor.scala 308:60]
  wire [7:0] _GEN_10251 = 8'h6 < length_3 ? _GEN_10091 : _GEN_9931; // @[executor.scala 308:60]
  wire [7:0] _GEN_10252 = 8'h6 < length_3 ? _GEN_10092 : _GEN_9932; // @[executor.scala 308:60]
  wire [7:0] _GEN_10253 = 8'h6 < length_3 ? _GEN_10093 : _GEN_9933; // @[executor.scala 308:60]
  wire [7:0] _GEN_10254 = 8'h6 < length_3 ? _GEN_10094 : _GEN_9934; // @[executor.scala 308:60]
  wire [7:0] _GEN_10255 = 8'h6 < length_3 ? _GEN_10095 : _GEN_9935; // @[executor.scala 308:60]
  wire [7:0] _GEN_10256 = 8'h6 < length_3 ? _GEN_10096 : _GEN_9936; // @[executor.scala 308:60]
  wire [7:0] _GEN_10257 = 8'h6 < length_3 ? _GEN_10097 : _GEN_9937; // @[executor.scala 308:60]
  wire [7:0] _GEN_10258 = 8'h6 < length_3 ? _GEN_10098 : _GEN_9938; // @[executor.scala 308:60]
  wire [7:0] _GEN_10259 = 8'h6 < length_3 ? _GEN_10099 : _GEN_9939; // @[executor.scala 308:60]
  wire [7:0] _GEN_10260 = 8'h6 < length_3 ? _GEN_10100 : _GEN_9940; // @[executor.scala 308:60]
  wire [7:0] _GEN_10261 = 8'h6 < length_3 ? _GEN_10101 : _GEN_9941; // @[executor.scala 308:60]
  wire [7:0] _GEN_10262 = 8'h6 < length_3 ? _GEN_10102 : _GEN_9942; // @[executor.scala 308:60]
  wire [7:0] _GEN_10263 = 8'h6 < length_3 ? _GEN_10103 : _GEN_9943; // @[executor.scala 308:60]
  wire [7:0] _GEN_10264 = 8'h6 < length_3 ? _GEN_10104 : _GEN_9944; // @[executor.scala 308:60]
  wire [7:0] _GEN_10265 = 8'h6 < length_3 ? _GEN_10105 : _GEN_9945; // @[executor.scala 308:60]
  wire [7:0] _GEN_10266 = 8'h6 < length_3 ? _GEN_10106 : _GEN_9946; // @[executor.scala 308:60]
  wire [7:0] _GEN_10267 = 8'h6 < length_3 ? _GEN_10107 : _GEN_9947; // @[executor.scala 308:60]
  wire [7:0] _GEN_10268 = 8'h6 < length_3 ? _GEN_10108 : _GEN_9948; // @[executor.scala 308:60]
  wire [7:0] _GEN_10269 = 8'h6 < length_3 ? _GEN_10109 : _GEN_9949; // @[executor.scala 308:60]
  wire [7:0] _GEN_10270 = 8'h6 < length_3 ? _GEN_10110 : _GEN_9950; // @[executor.scala 308:60]
  wire [7:0] _GEN_10271 = 8'h6 < length_3 ? _GEN_10111 : _GEN_9951; // @[executor.scala 308:60]
  wire [7:0] _GEN_10272 = 8'h6 < length_3 ? _GEN_10112 : _GEN_9952; // @[executor.scala 308:60]
  wire [7:0] _GEN_10273 = 8'h6 < length_3 ? _GEN_10113 : _GEN_9953; // @[executor.scala 308:60]
  wire [7:0] _GEN_10274 = 8'h6 < length_3 ? _GEN_10114 : _GEN_9954; // @[executor.scala 308:60]
  wire [7:0] _GEN_10275 = 8'h6 < length_3 ? _GEN_10115 : _GEN_9955; // @[executor.scala 308:60]
  wire [7:0] _GEN_10276 = 8'h6 < length_3 ? _GEN_10116 : _GEN_9956; // @[executor.scala 308:60]
  wire [7:0] _GEN_10277 = 8'h6 < length_3 ? _GEN_10117 : _GEN_9957; // @[executor.scala 308:60]
  wire [7:0] _GEN_10278 = 8'h6 < length_3 ? _GEN_10118 : _GEN_9958; // @[executor.scala 308:60]
  wire [7:0] _GEN_10279 = 8'h6 < length_3 ? _GEN_10119 : _GEN_9959; // @[executor.scala 308:60]
  wire [7:0] _GEN_10280 = 8'h6 < length_3 ? _GEN_10120 : _GEN_9960; // @[executor.scala 308:60]
  wire [7:0] _GEN_10281 = 8'h6 < length_3 ? _GEN_10121 : _GEN_9961; // @[executor.scala 308:60]
  wire [7:0] _GEN_10282 = 8'h6 < length_3 ? _GEN_10122 : _GEN_9962; // @[executor.scala 308:60]
  wire [7:0] _GEN_10283 = 8'h6 < length_3 ? _GEN_10123 : _GEN_9963; // @[executor.scala 308:60]
  wire [7:0] _GEN_10284 = 8'h6 < length_3 ? _GEN_10124 : _GEN_9964; // @[executor.scala 308:60]
  wire [7:0] _GEN_10285 = 8'h6 < length_3 ? _GEN_10125 : _GEN_9965; // @[executor.scala 308:60]
  wire [7:0] _GEN_10286 = 8'h6 < length_3 ? _GEN_10126 : _GEN_9966; // @[executor.scala 308:60]
  wire [7:0] _GEN_10287 = 8'h6 < length_3 ? _GEN_10127 : _GEN_9967; // @[executor.scala 308:60]
  wire [7:0] _GEN_10288 = 8'h6 < length_3 ? _GEN_10128 : _GEN_9968; // @[executor.scala 308:60]
  wire [7:0] _GEN_10289 = 8'h6 < length_3 ? _GEN_10129 : _GEN_9969; // @[executor.scala 308:60]
  wire [7:0] _GEN_10290 = 8'h6 < length_3 ? _GEN_10130 : _GEN_9970; // @[executor.scala 308:60]
  wire [7:0] _GEN_10291 = 8'h6 < length_3 ? _GEN_10131 : _GEN_9971; // @[executor.scala 308:60]
  wire [7:0] _GEN_10292 = 8'h6 < length_3 ? _GEN_10132 : _GEN_9972; // @[executor.scala 308:60]
  wire [7:0] _GEN_10293 = 8'h6 < length_3 ? _GEN_10133 : _GEN_9973; // @[executor.scala 308:60]
  wire [7:0] _GEN_10294 = 8'h6 < length_3 ? _GEN_10134 : _GEN_9974; // @[executor.scala 308:60]
  wire [7:0] _GEN_10295 = 8'h6 < length_3 ? _GEN_10135 : _GEN_9975; // @[executor.scala 308:60]
  wire [7:0] _GEN_10296 = 8'h6 < length_3 ? _GEN_10136 : _GEN_9976; // @[executor.scala 308:60]
  wire [7:0] _GEN_10297 = 8'h6 < length_3 ? _GEN_10137 : _GEN_9977; // @[executor.scala 308:60]
  wire [7:0] _GEN_10298 = 8'h6 < length_3 ? _GEN_10138 : _GEN_9978; // @[executor.scala 308:60]
  wire [7:0] _GEN_10299 = 8'h6 < length_3 ? _GEN_10139 : _GEN_9979; // @[executor.scala 308:60]
  wire [7:0] _GEN_10300 = 8'h6 < length_3 ? _GEN_10140 : _GEN_9980; // @[executor.scala 308:60]
  wire [7:0] _GEN_10301 = 8'h6 < length_3 ? _GEN_10141 : _GEN_9981; // @[executor.scala 308:60]
  wire [7:0] _GEN_10302 = 8'h6 < length_3 ? _GEN_10142 : _GEN_9982; // @[executor.scala 308:60]
  wire [7:0] _GEN_10303 = 8'h6 < length_3 ? _GEN_10143 : _GEN_9983; // @[executor.scala 308:60]
  wire [7:0] _GEN_10304 = 8'h6 < length_3 ? _GEN_10144 : _GEN_9984; // @[executor.scala 308:60]
  wire [7:0] _GEN_10305 = 8'h6 < length_3 ? _GEN_10145 : _GEN_9985; // @[executor.scala 308:60]
  wire [7:0] _GEN_10306 = 8'h6 < length_3 ? _GEN_10146 : _GEN_9986; // @[executor.scala 308:60]
  wire [7:0] _GEN_10307 = 8'h6 < length_3 ? _GEN_10147 : _GEN_9987; // @[executor.scala 308:60]
  wire [7:0] _GEN_10308 = 8'h6 < length_3 ? _GEN_10148 : _GEN_9988; // @[executor.scala 308:60]
  wire [7:0] _GEN_10309 = 8'h6 < length_3 ? _GEN_10149 : _GEN_9989; // @[executor.scala 308:60]
  wire [7:0] _GEN_10310 = 8'h6 < length_3 ? _GEN_10150 : _GEN_9990; // @[executor.scala 308:60]
  wire [7:0] _GEN_10311 = 8'h6 < length_3 ? _GEN_10151 : _GEN_9991; // @[executor.scala 308:60]
  wire [7:0] _GEN_10312 = 8'h6 < length_3 ? _GEN_10152 : _GEN_9992; // @[executor.scala 308:60]
  wire [7:0] _GEN_10313 = 8'h6 < length_3 ? _GEN_10153 : _GEN_9993; // @[executor.scala 308:60]
  wire [7:0] _GEN_10314 = 8'h6 < length_3 ? _GEN_10154 : _GEN_9994; // @[executor.scala 308:60]
  wire [7:0] _GEN_10315 = 8'h6 < length_3 ? _GEN_10155 : _GEN_9995; // @[executor.scala 308:60]
  wire [7:0] _GEN_10316 = 8'h6 < length_3 ? _GEN_10156 : _GEN_9996; // @[executor.scala 308:60]
  wire [7:0] _GEN_10317 = 8'h6 < length_3 ? _GEN_10157 : _GEN_9997; // @[executor.scala 308:60]
  wire [7:0] _GEN_10318 = 8'h6 < length_3 ? _GEN_10158 : _GEN_9998; // @[executor.scala 308:60]
  wire [7:0] _GEN_10319 = 8'h6 < length_3 ? _GEN_10159 : _GEN_9999; // @[executor.scala 308:60]
  wire [7:0] _GEN_10320 = 8'h6 < length_3 ? _GEN_10160 : _GEN_10000; // @[executor.scala 308:60]
  wire [7:0] _GEN_10321 = 8'h6 < length_3 ? _GEN_10161 : _GEN_10001; // @[executor.scala 308:60]
  wire [7:0] _GEN_10322 = 8'h6 < length_3 ? _GEN_10162 : _GEN_10002; // @[executor.scala 308:60]
  wire [7:0] _GEN_10323 = 8'h6 < length_3 ? _GEN_10163 : _GEN_10003; // @[executor.scala 308:60]
  wire [7:0] _GEN_10324 = 8'h6 < length_3 ? _GEN_10164 : _GEN_10004; // @[executor.scala 308:60]
  wire [7:0] _GEN_10325 = 8'h6 < length_3 ? _GEN_10165 : _GEN_10005; // @[executor.scala 308:60]
  wire [7:0] _GEN_10326 = 8'h6 < length_3 ? _GEN_10166 : _GEN_10006; // @[executor.scala 308:60]
  wire [7:0] _GEN_10327 = 8'h6 < length_3 ? _GEN_10167 : _GEN_10007; // @[executor.scala 308:60]
  wire [7:0] _GEN_10328 = 8'h6 < length_3 ? _GEN_10168 : _GEN_10008; // @[executor.scala 308:60]
  wire [7:0] _GEN_10329 = 8'h6 < length_3 ? _GEN_10169 : _GEN_10009; // @[executor.scala 308:60]
  wire [7:0] _GEN_10330 = 8'h6 < length_3 ? _GEN_10170 : _GEN_10010; // @[executor.scala 308:60]
  wire [7:0] _GEN_10331 = 8'h6 < length_3 ? _GEN_10171 : _GEN_10011; // @[executor.scala 308:60]
  wire [7:0] _GEN_10332 = 8'h6 < length_3 ? _GEN_10172 : _GEN_10012; // @[executor.scala 308:60]
  wire [7:0] _GEN_10333 = 8'h6 < length_3 ? _GEN_10173 : _GEN_10013; // @[executor.scala 308:60]
  wire [7:0] _GEN_10334 = 8'h6 < length_3 ? _GEN_10174 : _GEN_10014; // @[executor.scala 308:60]
  wire [7:0] _GEN_10335 = 8'h6 < length_3 ? _GEN_10175 : _GEN_10015; // @[executor.scala 308:60]
  wire [7:0] _GEN_10336 = 8'h6 < length_3 ? _GEN_10176 : _GEN_10016; // @[executor.scala 308:60]
  wire [7:0] _GEN_10337 = 8'h6 < length_3 ? _GEN_10177 : _GEN_10017; // @[executor.scala 308:60]
  wire [7:0] _GEN_10338 = 8'h6 < length_3 ? _GEN_10178 : _GEN_10018; // @[executor.scala 308:60]
  wire [7:0] _GEN_10339 = 8'h6 < length_3 ? _GEN_10179 : _GEN_10019; // @[executor.scala 308:60]
  wire [7:0] _GEN_10340 = 8'h6 < length_3 ? _GEN_10180 : _GEN_10020; // @[executor.scala 308:60]
  wire [7:0] _GEN_10341 = 8'h6 < length_3 ? _GEN_10181 : _GEN_10021; // @[executor.scala 308:60]
  wire [7:0] _GEN_10342 = 8'h6 < length_3 ? _GEN_10182 : _GEN_10022; // @[executor.scala 308:60]
  wire [7:0] _GEN_10343 = 8'h6 < length_3 ? _GEN_10183 : _GEN_10023; // @[executor.scala 308:60]
  wire [7:0] _GEN_10344 = 8'h6 < length_3 ? _GEN_10184 : _GEN_10024; // @[executor.scala 308:60]
  wire [7:0] _GEN_10345 = 8'h6 < length_3 ? _GEN_10185 : _GEN_10025; // @[executor.scala 308:60]
  wire [7:0] _GEN_10346 = 8'h6 < length_3 ? _GEN_10186 : _GEN_10026; // @[executor.scala 308:60]
  wire [7:0] _GEN_10347 = 8'h6 < length_3 ? _GEN_10187 : _GEN_10027; // @[executor.scala 308:60]
  wire [7:0] _GEN_10348 = 8'h6 < length_3 ? _GEN_10188 : _GEN_10028; // @[executor.scala 308:60]
  wire [7:0] _GEN_10349 = 8'h6 < length_3 ? _GEN_10189 : _GEN_10029; // @[executor.scala 308:60]
  wire [7:0] _GEN_10350 = 8'h6 < length_3 ? _GEN_10190 : _GEN_10030; // @[executor.scala 308:60]
  wire [7:0] _GEN_10351 = 8'h6 < length_3 ? _GEN_10191 : _GEN_10031; // @[executor.scala 308:60]
  wire [7:0] _GEN_10352 = 8'h6 < length_3 ? _GEN_10192 : _GEN_10032; // @[executor.scala 308:60]
  wire [7:0] _GEN_10353 = 8'h6 < length_3 ? _GEN_10193 : _GEN_10033; // @[executor.scala 308:60]
  wire [7:0] _GEN_10354 = 8'h6 < length_3 ? _GEN_10194 : _GEN_10034; // @[executor.scala 308:60]
  wire [7:0] _GEN_10355 = 8'h6 < length_3 ? _GEN_10195 : _GEN_10035; // @[executor.scala 308:60]
  wire [7:0] _GEN_10356 = 8'h6 < length_3 ? _GEN_10196 : _GEN_10036; // @[executor.scala 308:60]
  wire [7:0] _GEN_10357 = 8'h6 < length_3 ? _GEN_10197 : _GEN_10037; // @[executor.scala 308:60]
  wire [7:0] _GEN_10358 = 8'h6 < length_3 ? _GEN_10198 : _GEN_10038; // @[executor.scala 308:60]
  wire [7:0] _GEN_10359 = 8'h6 < length_3 ? _GEN_10199 : _GEN_10039; // @[executor.scala 308:60]
  wire [7:0] _GEN_10360 = 8'h6 < length_3 ? _GEN_10200 : _GEN_10040; // @[executor.scala 308:60]
  wire [7:0] _GEN_10361 = 8'h6 < length_3 ? _GEN_10201 : _GEN_10041; // @[executor.scala 308:60]
  wire [7:0] _GEN_10362 = 8'h6 < length_3 ? _GEN_10202 : _GEN_10042; // @[executor.scala 308:60]
  wire [7:0] _GEN_10363 = 8'h6 < length_3 ? _GEN_10203 : _GEN_10043; // @[executor.scala 308:60]
  wire [7:0] _GEN_10364 = 8'h6 < length_3 ? _GEN_10204 : _GEN_10044; // @[executor.scala 308:60]
  wire [7:0] _GEN_10365 = 8'h6 < length_3 ? _GEN_10205 : _GEN_10045; // @[executor.scala 308:60]
  wire [7:0] _GEN_10366 = 8'h6 < length_3 ? _GEN_10206 : _GEN_10046; // @[executor.scala 308:60]
  wire [7:0] _GEN_10367 = 8'h6 < length_3 ? _GEN_10207 : _GEN_10047; // @[executor.scala 308:60]
  wire [7:0] _GEN_10368 = 8'h6 < length_3 ? _GEN_10208 : _GEN_10048; // @[executor.scala 308:60]
  wire [7:0] _GEN_10369 = 8'h6 < length_3 ? _GEN_10209 : _GEN_10049; // @[executor.scala 308:60]
  wire [7:0] _GEN_10370 = 8'h6 < length_3 ? _GEN_10210 : _GEN_10050; // @[executor.scala 308:60]
  wire [7:0] _GEN_10371 = 8'h6 < length_3 ? _GEN_10211 : _GEN_10051; // @[executor.scala 308:60]
  wire [7:0] _GEN_10372 = 8'h6 < length_3 ? _GEN_10212 : _GEN_10052; // @[executor.scala 308:60]
  wire [7:0] _GEN_10373 = 8'h6 < length_3 ? _GEN_10213 : _GEN_10053; // @[executor.scala 308:60]
  wire [7:0] _GEN_10374 = 8'h6 < length_3 ? _GEN_10214 : _GEN_10054; // @[executor.scala 308:60]
  wire [7:0] _GEN_10375 = 8'h6 < length_3 ? _GEN_10215 : _GEN_10055; // @[executor.scala 308:60]
  wire [7:0] _GEN_10376 = 8'h6 < length_3 ? _GEN_10216 : _GEN_10056; // @[executor.scala 308:60]
  wire [7:0] _GEN_10377 = 8'h6 < length_3 ? _GEN_10217 : _GEN_10057; // @[executor.scala 308:60]
  wire [7:0] _GEN_10378 = 8'h6 < length_3 ? _GEN_10218 : _GEN_10058; // @[executor.scala 308:60]
  wire [7:0] _GEN_10379 = 8'h6 < length_3 ? _GEN_10219 : _GEN_10059; // @[executor.scala 308:60]
  wire [7:0] _GEN_10380 = 8'h6 < length_3 ? _GEN_10220 : _GEN_10060; // @[executor.scala 308:60]
  wire [7:0] _GEN_10381 = 8'h6 < length_3 ? _GEN_10221 : _GEN_10061; // @[executor.scala 308:60]
  wire [7:0] _GEN_10382 = 8'h6 < length_3 ? _GEN_10222 : _GEN_10062; // @[executor.scala 308:60]
  wire [7:0] _GEN_10383 = 8'h6 < length_3 ? _GEN_10223 : _GEN_10063; // @[executor.scala 308:60]
  wire [7:0] _GEN_10384 = 8'h6 < length_3 ? _GEN_10224 : _GEN_10064; // @[executor.scala 308:60]
  wire [7:0] _GEN_10385 = 8'h6 < length_3 ? _GEN_10225 : _GEN_10065; // @[executor.scala 308:60]
  wire [7:0] _GEN_10386 = 8'h6 < length_3 ? _GEN_10226 : _GEN_10066; // @[executor.scala 308:60]
  wire [7:0] _GEN_10387 = 8'h6 < length_3 ? _GEN_10227 : _GEN_10067; // @[executor.scala 308:60]
  wire [7:0] _GEN_10388 = 8'h6 < length_3 ? _GEN_10228 : _GEN_10068; // @[executor.scala 308:60]
  wire [7:0] _GEN_10389 = 8'h6 < length_3 ? _GEN_10229 : _GEN_10069; // @[executor.scala 308:60]
  wire [7:0] _GEN_10390 = 8'h6 < length_3 ? _GEN_10230 : _GEN_10070; // @[executor.scala 308:60]
  wire [7:0] _GEN_10391 = 8'h6 < length_3 ? _GEN_10231 : _GEN_10071; // @[executor.scala 308:60]
  wire [7:0] _GEN_10392 = 8'h6 < length_3 ? _GEN_10232 : _GEN_10072; // @[executor.scala 308:60]
  wire [7:0] _GEN_10393 = 8'h6 < length_3 ? _GEN_10233 : _GEN_10073; // @[executor.scala 308:60]
  wire [7:0] _GEN_10394 = 8'h6 < length_3 ? _GEN_10234 : _GEN_10074; // @[executor.scala 308:60]
  wire [7:0] _GEN_10395 = 8'h6 < length_3 ? _GEN_10235 : _GEN_10075; // @[executor.scala 308:60]
  wire [7:0] _GEN_10396 = 8'h6 < length_3 ? _GEN_10236 : _GEN_10076; // @[executor.scala 308:60]
  wire [7:0] _GEN_10397 = 8'h6 < length_3 ? _GEN_10237 : _GEN_10077; // @[executor.scala 308:60]
  wire [7:0] _GEN_10398 = 8'h6 < length_3 ? _GEN_10238 : _GEN_10078; // @[executor.scala 308:60]
  wire [7:0] _GEN_10399 = 8'h6 < length_3 ? _GEN_10239 : _GEN_10079; // @[executor.scala 308:60]
  wire [7:0] _GEN_10400 = 8'h6 < length_3 ? _GEN_10240 : _GEN_10080; // @[executor.scala 308:60]
  wire [7:0] _GEN_10401 = 8'h6 < length_3 ? _GEN_10241 : _GEN_10081; // @[executor.scala 308:60]
  wire [7:0] _GEN_10402 = 8'h6 < length_3 ? _GEN_10242 : _GEN_10082; // @[executor.scala 308:60]
  wire [7:0] _GEN_10403 = 8'h6 < length_3 ? _GEN_10243 : _GEN_10083; // @[executor.scala 308:60]
  wire [7:0] _GEN_10404 = 8'h6 < length_3 ? _GEN_10244 : _GEN_10084; // @[executor.scala 308:60]
  wire [7:0] _GEN_10405 = 8'h6 < length_3 ? _GEN_10245 : _GEN_10085; // @[executor.scala 308:60]
  wire [7:0] field_byte_31 = field_3[7:0]; // @[executor.scala 305:57]
  wire [7:0] total_offset_31 = offset_3 + 8'h7; // @[executor.scala 307:57]
  wire [7:0] _GEN_10406 = 8'h0 == total_offset_31 ? field_byte_31 : _GEN_10246; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10407 = 8'h1 == total_offset_31 ? field_byte_31 : _GEN_10247; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10408 = 8'h2 == total_offset_31 ? field_byte_31 : _GEN_10248; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10409 = 8'h3 == total_offset_31 ? field_byte_31 : _GEN_10249; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10410 = 8'h4 == total_offset_31 ? field_byte_31 : _GEN_10250; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10411 = 8'h5 == total_offset_31 ? field_byte_31 : _GEN_10251; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10412 = 8'h6 == total_offset_31 ? field_byte_31 : _GEN_10252; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10413 = 8'h7 == total_offset_31 ? field_byte_31 : _GEN_10253; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10414 = 8'h8 == total_offset_31 ? field_byte_31 : _GEN_10254; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10415 = 8'h9 == total_offset_31 ? field_byte_31 : _GEN_10255; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10416 = 8'ha == total_offset_31 ? field_byte_31 : _GEN_10256; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10417 = 8'hb == total_offset_31 ? field_byte_31 : _GEN_10257; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10418 = 8'hc == total_offset_31 ? field_byte_31 : _GEN_10258; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10419 = 8'hd == total_offset_31 ? field_byte_31 : _GEN_10259; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10420 = 8'he == total_offset_31 ? field_byte_31 : _GEN_10260; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10421 = 8'hf == total_offset_31 ? field_byte_31 : _GEN_10261; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10422 = 8'h10 == total_offset_31 ? field_byte_31 : _GEN_10262; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10423 = 8'h11 == total_offset_31 ? field_byte_31 : _GEN_10263; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10424 = 8'h12 == total_offset_31 ? field_byte_31 : _GEN_10264; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10425 = 8'h13 == total_offset_31 ? field_byte_31 : _GEN_10265; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10426 = 8'h14 == total_offset_31 ? field_byte_31 : _GEN_10266; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10427 = 8'h15 == total_offset_31 ? field_byte_31 : _GEN_10267; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10428 = 8'h16 == total_offset_31 ? field_byte_31 : _GEN_10268; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10429 = 8'h17 == total_offset_31 ? field_byte_31 : _GEN_10269; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10430 = 8'h18 == total_offset_31 ? field_byte_31 : _GEN_10270; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10431 = 8'h19 == total_offset_31 ? field_byte_31 : _GEN_10271; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10432 = 8'h1a == total_offset_31 ? field_byte_31 : _GEN_10272; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10433 = 8'h1b == total_offset_31 ? field_byte_31 : _GEN_10273; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10434 = 8'h1c == total_offset_31 ? field_byte_31 : _GEN_10274; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10435 = 8'h1d == total_offset_31 ? field_byte_31 : _GEN_10275; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10436 = 8'h1e == total_offset_31 ? field_byte_31 : _GEN_10276; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10437 = 8'h1f == total_offset_31 ? field_byte_31 : _GEN_10277; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10438 = 8'h20 == total_offset_31 ? field_byte_31 : _GEN_10278; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10439 = 8'h21 == total_offset_31 ? field_byte_31 : _GEN_10279; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10440 = 8'h22 == total_offset_31 ? field_byte_31 : _GEN_10280; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10441 = 8'h23 == total_offset_31 ? field_byte_31 : _GEN_10281; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10442 = 8'h24 == total_offset_31 ? field_byte_31 : _GEN_10282; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10443 = 8'h25 == total_offset_31 ? field_byte_31 : _GEN_10283; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10444 = 8'h26 == total_offset_31 ? field_byte_31 : _GEN_10284; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10445 = 8'h27 == total_offset_31 ? field_byte_31 : _GEN_10285; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10446 = 8'h28 == total_offset_31 ? field_byte_31 : _GEN_10286; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10447 = 8'h29 == total_offset_31 ? field_byte_31 : _GEN_10287; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10448 = 8'h2a == total_offset_31 ? field_byte_31 : _GEN_10288; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10449 = 8'h2b == total_offset_31 ? field_byte_31 : _GEN_10289; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10450 = 8'h2c == total_offset_31 ? field_byte_31 : _GEN_10290; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10451 = 8'h2d == total_offset_31 ? field_byte_31 : _GEN_10291; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10452 = 8'h2e == total_offset_31 ? field_byte_31 : _GEN_10292; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10453 = 8'h2f == total_offset_31 ? field_byte_31 : _GEN_10293; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10454 = 8'h30 == total_offset_31 ? field_byte_31 : _GEN_10294; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10455 = 8'h31 == total_offset_31 ? field_byte_31 : _GEN_10295; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10456 = 8'h32 == total_offset_31 ? field_byte_31 : _GEN_10296; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10457 = 8'h33 == total_offset_31 ? field_byte_31 : _GEN_10297; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10458 = 8'h34 == total_offset_31 ? field_byte_31 : _GEN_10298; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10459 = 8'h35 == total_offset_31 ? field_byte_31 : _GEN_10299; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10460 = 8'h36 == total_offset_31 ? field_byte_31 : _GEN_10300; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10461 = 8'h37 == total_offset_31 ? field_byte_31 : _GEN_10301; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10462 = 8'h38 == total_offset_31 ? field_byte_31 : _GEN_10302; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10463 = 8'h39 == total_offset_31 ? field_byte_31 : _GEN_10303; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10464 = 8'h3a == total_offset_31 ? field_byte_31 : _GEN_10304; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10465 = 8'h3b == total_offset_31 ? field_byte_31 : _GEN_10305; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10466 = 8'h3c == total_offset_31 ? field_byte_31 : _GEN_10306; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10467 = 8'h3d == total_offset_31 ? field_byte_31 : _GEN_10307; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10468 = 8'h3e == total_offset_31 ? field_byte_31 : _GEN_10308; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10469 = 8'h3f == total_offset_31 ? field_byte_31 : _GEN_10309; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10470 = 8'h40 == total_offset_31 ? field_byte_31 : _GEN_10310; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10471 = 8'h41 == total_offset_31 ? field_byte_31 : _GEN_10311; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10472 = 8'h42 == total_offset_31 ? field_byte_31 : _GEN_10312; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10473 = 8'h43 == total_offset_31 ? field_byte_31 : _GEN_10313; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10474 = 8'h44 == total_offset_31 ? field_byte_31 : _GEN_10314; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10475 = 8'h45 == total_offset_31 ? field_byte_31 : _GEN_10315; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10476 = 8'h46 == total_offset_31 ? field_byte_31 : _GEN_10316; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10477 = 8'h47 == total_offset_31 ? field_byte_31 : _GEN_10317; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10478 = 8'h48 == total_offset_31 ? field_byte_31 : _GEN_10318; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10479 = 8'h49 == total_offset_31 ? field_byte_31 : _GEN_10319; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10480 = 8'h4a == total_offset_31 ? field_byte_31 : _GEN_10320; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10481 = 8'h4b == total_offset_31 ? field_byte_31 : _GEN_10321; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10482 = 8'h4c == total_offset_31 ? field_byte_31 : _GEN_10322; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10483 = 8'h4d == total_offset_31 ? field_byte_31 : _GEN_10323; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10484 = 8'h4e == total_offset_31 ? field_byte_31 : _GEN_10324; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10485 = 8'h4f == total_offset_31 ? field_byte_31 : _GEN_10325; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10486 = 8'h50 == total_offset_31 ? field_byte_31 : _GEN_10326; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10487 = 8'h51 == total_offset_31 ? field_byte_31 : _GEN_10327; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10488 = 8'h52 == total_offset_31 ? field_byte_31 : _GEN_10328; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10489 = 8'h53 == total_offset_31 ? field_byte_31 : _GEN_10329; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10490 = 8'h54 == total_offset_31 ? field_byte_31 : _GEN_10330; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10491 = 8'h55 == total_offset_31 ? field_byte_31 : _GEN_10331; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10492 = 8'h56 == total_offset_31 ? field_byte_31 : _GEN_10332; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10493 = 8'h57 == total_offset_31 ? field_byte_31 : _GEN_10333; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10494 = 8'h58 == total_offset_31 ? field_byte_31 : _GEN_10334; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10495 = 8'h59 == total_offset_31 ? field_byte_31 : _GEN_10335; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10496 = 8'h5a == total_offset_31 ? field_byte_31 : _GEN_10336; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10497 = 8'h5b == total_offset_31 ? field_byte_31 : _GEN_10337; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10498 = 8'h5c == total_offset_31 ? field_byte_31 : _GEN_10338; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10499 = 8'h5d == total_offset_31 ? field_byte_31 : _GEN_10339; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10500 = 8'h5e == total_offset_31 ? field_byte_31 : _GEN_10340; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10501 = 8'h5f == total_offset_31 ? field_byte_31 : _GEN_10341; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10502 = 8'h60 == total_offset_31 ? field_byte_31 : _GEN_10342; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10503 = 8'h61 == total_offset_31 ? field_byte_31 : _GEN_10343; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10504 = 8'h62 == total_offset_31 ? field_byte_31 : _GEN_10344; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10505 = 8'h63 == total_offset_31 ? field_byte_31 : _GEN_10345; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10506 = 8'h64 == total_offset_31 ? field_byte_31 : _GEN_10346; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10507 = 8'h65 == total_offset_31 ? field_byte_31 : _GEN_10347; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10508 = 8'h66 == total_offset_31 ? field_byte_31 : _GEN_10348; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10509 = 8'h67 == total_offset_31 ? field_byte_31 : _GEN_10349; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10510 = 8'h68 == total_offset_31 ? field_byte_31 : _GEN_10350; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10511 = 8'h69 == total_offset_31 ? field_byte_31 : _GEN_10351; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10512 = 8'h6a == total_offset_31 ? field_byte_31 : _GEN_10352; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10513 = 8'h6b == total_offset_31 ? field_byte_31 : _GEN_10353; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10514 = 8'h6c == total_offset_31 ? field_byte_31 : _GEN_10354; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10515 = 8'h6d == total_offset_31 ? field_byte_31 : _GEN_10355; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10516 = 8'h6e == total_offset_31 ? field_byte_31 : _GEN_10356; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10517 = 8'h6f == total_offset_31 ? field_byte_31 : _GEN_10357; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10518 = 8'h70 == total_offset_31 ? field_byte_31 : _GEN_10358; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10519 = 8'h71 == total_offset_31 ? field_byte_31 : _GEN_10359; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10520 = 8'h72 == total_offset_31 ? field_byte_31 : _GEN_10360; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10521 = 8'h73 == total_offset_31 ? field_byte_31 : _GEN_10361; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10522 = 8'h74 == total_offset_31 ? field_byte_31 : _GEN_10362; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10523 = 8'h75 == total_offset_31 ? field_byte_31 : _GEN_10363; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10524 = 8'h76 == total_offset_31 ? field_byte_31 : _GEN_10364; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10525 = 8'h77 == total_offset_31 ? field_byte_31 : _GEN_10365; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10526 = 8'h78 == total_offset_31 ? field_byte_31 : _GEN_10366; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10527 = 8'h79 == total_offset_31 ? field_byte_31 : _GEN_10367; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10528 = 8'h7a == total_offset_31 ? field_byte_31 : _GEN_10368; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10529 = 8'h7b == total_offset_31 ? field_byte_31 : _GEN_10369; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10530 = 8'h7c == total_offset_31 ? field_byte_31 : _GEN_10370; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10531 = 8'h7d == total_offset_31 ? field_byte_31 : _GEN_10371; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10532 = 8'h7e == total_offset_31 ? field_byte_31 : _GEN_10372; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10533 = 8'h7f == total_offset_31 ? field_byte_31 : _GEN_10373; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10534 = 8'h80 == total_offset_31 ? field_byte_31 : _GEN_10374; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10535 = 8'h81 == total_offset_31 ? field_byte_31 : _GEN_10375; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10536 = 8'h82 == total_offset_31 ? field_byte_31 : _GEN_10376; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10537 = 8'h83 == total_offset_31 ? field_byte_31 : _GEN_10377; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10538 = 8'h84 == total_offset_31 ? field_byte_31 : _GEN_10378; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10539 = 8'h85 == total_offset_31 ? field_byte_31 : _GEN_10379; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10540 = 8'h86 == total_offset_31 ? field_byte_31 : _GEN_10380; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10541 = 8'h87 == total_offset_31 ? field_byte_31 : _GEN_10381; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10542 = 8'h88 == total_offset_31 ? field_byte_31 : _GEN_10382; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10543 = 8'h89 == total_offset_31 ? field_byte_31 : _GEN_10383; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10544 = 8'h8a == total_offset_31 ? field_byte_31 : _GEN_10384; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10545 = 8'h8b == total_offset_31 ? field_byte_31 : _GEN_10385; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10546 = 8'h8c == total_offset_31 ? field_byte_31 : _GEN_10386; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10547 = 8'h8d == total_offset_31 ? field_byte_31 : _GEN_10387; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10548 = 8'h8e == total_offset_31 ? field_byte_31 : _GEN_10388; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10549 = 8'h8f == total_offset_31 ? field_byte_31 : _GEN_10389; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10550 = 8'h90 == total_offset_31 ? field_byte_31 : _GEN_10390; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10551 = 8'h91 == total_offset_31 ? field_byte_31 : _GEN_10391; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10552 = 8'h92 == total_offset_31 ? field_byte_31 : _GEN_10392; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10553 = 8'h93 == total_offset_31 ? field_byte_31 : _GEN_10393; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10554 = 8'h94 == total_offset_31 ? field_byte_31 : _GEN_10394; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10555 = 8'h95 == total_offset_31 ? field_byte_31 : _GEN_10395; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10556 = 8'h96 == total_offset_31 ? field_byte_31 : _GEN_10396; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10557 = 8'h97 == total_offset_31 ? field_byte_31 : _GEN_10397; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10558 = 8'h98 == total_offset_31 ? field_byte_31 : _GEN_10398; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10559 = 8'h99 == total_offset_31 ? field_byte_31 : _GEN_10399; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10560 = 8'h9a == total_offset_31 ? field_byte_31 : _GEN_10400; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10561 = 8'h9b == total_offset_31 ? field_byte_31 : _GEN_10401; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10562 = 8'h9c == total_offset_31 ? field_byte_31 : _GEN_10402; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10563 = 8'h9d == total_offset_31 ? field_byte_31 : _GEN_10403; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10564 = 8'h9e == total_offset_31 ? field_byte_31 : _GEN_10404; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10565 = 8'h9f == total_offset_31 ? field_byte_31 : _GEN_10405; // @[executor.scala 309:64 executor.scala 309:64]
  wire [7:0] _GEN_10566 = 8'h7 < length_3 ? _GEN_10406 : _GEN_10246; // @[executor.scala 308:60]
  wire [7:0] _GEN_10567 = 8'h7 < length_3 ? _GEN_10407 : _GEN_10247; // @[executor.scala 308:60]
  wire [7:0] _GEN_10568 = 8'h7 < length_3 ? _GEN_10408 : _GEN_10248; // @[executor.scala 308:60]
  wire [7:0] _GEN_10569 = 8'h7 < length_3 ? _GEN_10409 : _GEN_10249; // @[executor.scala 308:60]
  wire [7:0] _GEN_10570 = 8'h7 < length_3 ? _GEN_10410 : _GEN_10250; // @[executor.scala 308:60]
  wire [7:0] _GEN_10571 = 8'h7 < length_3 ? _GEN_10411 : _GEN_10251; // @[executor.scala 308:60]
  wire [7:0] _GEN_10572 = 8'h7 < length_3 ? _GEN_10412 : _GEN_10252; // @[executor.scala 308:60]
  wire [7:0] _GEN_10573 = 8'h7 < length_3 ? _GEN_10413 : _GEN_10253; // @[executor.scala 308:60]
  wire [7:0] _GEN_10574 = 8'h7 < length_3 ? _GEN_10414 : _GEN_10254; // @[executor.scala 308:60]
  wire [7:0] _GEN_10575 = 8'h7 < length_3 ? _GEN_10415 : _GEN_10255; // @[executor.scala 308:60]
  wire [7:0] _GEN_10576 = 8'h7 < length_3 ? _GEN_10416 : _GEN_10256; // @[executor.scala 308:60]
  wire [7:0] _GEN_10577 = 8'h7 < length_3 ? _GEN_10417 : _GEN_10257; // @[executor.scala 308:60]
  wire [7:0] _GEN_10578 = 8'h7 < length_3 ? _GEN_10418 : _GEN_10258; // @[executor.scala 308:60]
  wire [7:0] _GEN_10579 = 8'h7 < length_3 ? _GEN_10419 : _GEN_10259; // @[executor.scala 308:60]
  wire [7:0] _GEN_10580 = 8'h7 < length_3 ? _GEN_10420 : _GEN_10260; // @[executor.scala 308:60]
  wire [7:0] _GEN_10581 = 8'h7 < length_3 ? _GEN_10421 : _GEN_10261; // @[executor.scala 308:60]
  wire [7:0] _GEN_10582 = 8'h7 < length_3 ? _GEN_10422 : _GEN_10262; // @[executor.scala 308:60]
  wire [7:0] _GEN_10583 = 8'h7 < length_3 ? _GEN_10423 : _GEN_10263; // @[executor.scala 308:60]
  wire [7:0] _GEN_10584 = 8'h7 < length_3 ? _GEN_10424 : _GEN_10264; // @[executor.scala 308:60]
  wire [7:0] _GEN_10585 = 8'h7 < length_3 ? _GEN_10425 : _GEN_10265; // @[executor.scala 308:60]
  wire [7:0] _GEN_10586 = 8'h7 < length_3 ? _GEN_10426 : _GEN_10266; // @[executor.scala 308:60]
  wire [7:0] _GEN_10587 = 8'h7 < length_3 ? _GEN_10427 : _GEN_10267; // @[executor.scala 308:60]
  wire [7:0] _GEN_10588 = 8'h7 < length_3 ? _GEN_10428 : _GEN_10268; // @[executor.scala 308:60]
  wire [7:0] _GEN_10589 = 8'h7 < length_3 ? _GEN_10429 : _GEN_10269; // @[executor.scala 308:60]
  wire [7:0] _GEN_10590 = 8'h7 < length_3 ? _GEN_10430 : _GEN_10270; // @[executor.scala 308:60]
  wire [7:0] _GEN_10591 = 8'h7 < length_3 ? _GEN_10431 : _GEN_10271; // @[executor.scala 308:60]
  wire [7:0] _GEN_10592 = 8'h7 < length_3 ? _GEN_10432 : _GEN_10272; // @[executor.scala 308:60]
  wire [7:0] _GEN_10593 = 8'h7 < length_3 ? _GEN_10433 : _GEN_10273; // @[executor.scala 308:60]
  wire [7:0] _GEN_10594 = 8'h7 < length_3 ? _GEN_10434 : _GEN_10274; // @[executor.scala 308:60]
  wire [7:0] _GEN_10595 = 8'h7 < length_3 ? _GEN_10435 : _GEN_10275; // @[executor.scala 308:60]
  wire [7:0] _GEN_10596 = 8'h7 < length_3 ? _GEN_10436 : _GEN_10276; // @[executor.scala 308:60]
  wire [7:0] _GEN_10597 = 8'h7 < length_3 ? _GEN_10437 : _GEN_10277; // @[executor.scala 308:60]
  wire [7:0] _GEN_10598 = 8'h7 < length_3 ? _GEN_10438 : _GEN_10278; // @[executor.scala 308:60]
  wire [7:0] _GEN_10599 = 8'h7 < length_3 ? _GEN_10439 : _GEN_10279; // @[executor.scala 308:60]
  wire [7:0] _GEN_10600 = 8'h7 < length_3 ? _GEN_10440 : _GEN_10280; // @[executor.scala 308:60]
  wire [7:0] _GEN_10601 = 8'h7 < length_3 ? _GEN_10441 : _GEN_10281; // @[executor.scala 308:60]
  wire [7:0] _GEN_10602 = 8'h7 < length_3 ? _GEN_10442 : _GEN_10282; // @[executor.scala 308:60]
  wire [7:0] _GEN_10603 = 8'h7 < length_3 ? _GEN_10443 : _GEN_10283; // @[executor.scala 308:60]
  wire [7:0] _GEN_10604 = 8'h7 < length_3 ? _GEN_10444 : _GEN_10284; // @[executor.scala 308:60]
  wire [7:0] _GEN_10605 = 8'h7 < length_3 ? _GEN_10445 : _GEN_10285; // @[executor.scala 308:60]
  wire [7:0] _GEN_10606 = 8'h7 < length_3 ? _GEN_10446 : _GEN_10286; // @[executor.scala 308:60]
  wire [7:0] _GEN_10607 = 8'h7 < length_3 ? _GEN_10447 : _GEN_10287; // @[executor.scala 308:60]
  wire [7:0] _GEN_10608 = 8'h7 < length_3 ? _GEN_10448 : _GEN_10288; // @[executor.scala 308:60]
  wire [7:0] _GEN_10609 = 8'h7 < length_3 ? _GEN_10449 : _GEN_10289; // @[executor.scala 308:60]
  wire [7:0] _GEN_10610 = 8'h7 < length_3 ? _GEN_10450 : _GEN_10290; // @[executor.scala 308:60]
  wire [7:0] _GEN_10611 = 8'h7 < length_3 ? _GEN_10451 : _GEN_10291; // @[executor.scala 308:60]
  wire [7:0] _GEN_10612 = 8'h7 < length_3 ? _GEN_10452 : _GEN_10292; // @[executor.scala 308:60]
  wire [7:0] _GEN_10613 = 8'h7 < length_3 ? _GEN_10453 : _GEN_10293; // @[executor.scala 308:60]
  wire [7:0] _GEN_10614 = 8'h7 < length_3 ? _GEN_10454 : _GEN_10294; // @[executor.scala 308:60]
  wire [7:0] _GEN_10615 = 8'h7 < length_3 ? _GEN_10455 : _GEN_10295; // @[executor.scala 308:60]
  wire [7:0] _GEN_10616 = 8'h7 < length_3 ? _GEN_10456 : _GEN_10296; // @[executor.scala 308:60]
  wire [7:0] _GEN_10617 = 8'h7 < length_3 ? _GEN_10457 : _GEN_10297; // @[executor.scala 308:60]
  wire [7:0] _GEN_10618 = 8'h7 < length_3 ? _GEN_10458 : _GEN_10298; // @[executor.scala 308:60]
  wire [7:0] _GEN_10619 = 8'h7 < length_3 ? _GEN_10459 : _GEN_10299; // @[executor.scala 308:60]
  wire [7:0] _GEN_10620 = 8'h7 < length_3 ? _GEN_10460 : _GEN_10300; // @[executor.scala 308:60]
  wire [7:0] _GEN_10621 = 8'h7 < length_3 ? _GEN_10461 : _GEN_10301; // @[executor.scala 308:60]
  wire [7:0] _GEN_10622 = 8'h7 < length_3 ? _GEN_10462 : _GEN_10302; // @[executor.scala 308:60]
  wire [7:0] _GEN_10623 = 8'h7 < length_3 ? _GEN_10463 : _GEN_10303; // @[executor.scala 308:60]
  wire [7:0] _GEN_10624 = 8'h7 < length_3 ? _GEN_10464 : _GEN_10304; // @[executor.scala 308:60]
  wire [7:0] _GEN_10625 = 8'h7 < length_3 ? _GEN_10465 : _GEN_10305; // @[executor.scala 308:60]
  wire [7:0] _GEN_10626 = 8'h7 < length_3 ? _GEN_10466 : _GEN_10306; // @[executor.scala 308:60]
  wire [7:0] _GEN_10627 = 8'h7 < length_3 ? _GEN_10467 : _GEN_10307; // @[executor.scala 308:60]
  wire [7:0] _GEN_10628 = 8'h7 < length_3 ? _GEN_10468 : _GEN_10308; // @[executor.scala 308:60]
  wire [7:0] _GEN_10629 = 8'h7 < length_3 ? _GEN_10469 : _GEN_10309; // @[executor.scala 308:60]
  wire [7:0] _GEN_10630 = 8'h7 < length_3 ? _GEN_10470 : _GEN_10310; // @[executor.scala 308:60]
  wire [7:0] _GEN_10631 = 8'h7 < length_3 ? _GEN_10471 : _GEN_10311; // @[executor.scala 308:60]
  wire [7:0] _GEN_10632 = 8'h7 < length_3 ? _GEN_10472 : _GEN_10312; // @[executor.scala 308:60]
  wire [7:0] _GEN_10633 = 8'h7 < length_3 ? _GEN_10473 : _GEN_10313; // @[executor.scala 308:60]
  wire [7:0] _GEN_10634 = 8'h7 < length_3 ? _GEN_10474 : _GEN_10314; // @[executor.scala 308:60]
  wire [7:0] _GEN_10635 = 8'h7 < length_3 ? _GEN_10475 : _GEN_10315; // @[executor.scala 308:60]
  wire [7:0] _GEN_10636 = 8'h7 < length_3 ? _GEN_10476 : _GEN_10316; // @[executor.scala 308:60]
  wire [7:0] _GEN_10637 = 8'h7 < length_3 ? _GEN_10477 : _GEN_10317; // @[executor.scala 308:60]
  wire [7:0] _GEN_10638 = 8'h7 < length_3 ? _GEN_10478 : _GEN_10318; // @[executor.scala 308:60]
  wire [7:0] _GEN_10639 = 8'h7 < length_3 ? _GEN_10479 : _GEN_10319; // @[executor.scala 308:60]
  wire [7:0] _GEN_10640 = 8'h7 < length_3 ? _GEN_10480 : _GEN_10320; // @[executor.scala 308:60]
  wire [7:0] _GEN_10641 = 8'h7 < length_3 ? _GEN_10481 : _GEN_10321; // @[executor.scala 308:60]
  wire [7:0] _GEN_10642 = 8'h7 < length_3 ? _GEN_10482 : _GEN_10322; // @[executor.scala 308:60]
  wire [7:0] _GEN_10643 = 8'h7 < length_3 ? _GEN_10483 : _GEN_10323; // @[executor.scala 308:60]
  wire [7:0] _GEN_10644 = 8'h7 < length_3 ? _GEN_10484 : _GEN_10324; // @[executor.scala 308:60]
  wire [7:0] _GEN_10645 = 8'h7 < length_3 ? _GEN_10485 : _GEN_10325; // @[executor.scala 308:60]
  wire [7:0] _GEN_10646 = 8'h7 < length_3 ? _GEN_10486 : _GEN_10326; // @[executor.scala 308:60]
  wire [7:0] _GEN_10647 = 8'h7 < length_3 ? _GEN_10487 : _GEN_10327; // @[executor.scala 308:60]
  wire [7:0] _GEN_10648 = 8'h7 < length_3 ? _GEN_10488 : _GEN_10328; // @[executor.scala 308:60]
  wire [7:0] _GEN_10649 = 8'h7 < length_3 ? _GEN_10489 : _GEN_10329; // @[executor.scala 308:60]
  wire [7:0] _GEN_10650 = 8'h7 < length_3 ? _GEN_10490 : _GEN_10330; // @[executor.scala 308:60]
  wire [7:0] _GEN_10651 = 8'h7 < length_3 ? _GEN_10491 : _GEN_10331; // @[executor.scala 308:60]
  wire [7:0] _GEN_10652 = 8'h7 < length_3 ? _GEN_10492 : _GEN_10332; // @[executor.scala 308:60]
  wire [7:0] _GEN_10653 = 8'h7 < length_3 ? _GEN_10493 : _GEN_10333; // @[executor.scala 308:60]
  wire [7:0] _GEN_10654 = 8'h7 < length_3 ? _GEN_10494 : _GEN_10334; // @[executor.scala 308:60]
  wire [7:0] _GEN_10655 = 8'h7 < length_3 ? _GEN_10495 : _GEN_10335; // @[executor.scala 308:60]
  wire [7:0] _GEN_10656 = 8'h7 < length_3 ? _GEN_10496 : _GEN_10336; // @[executor.scala 308:60]
  wire [7:0] _GEN_10657 = 8'h7 < length_3 ? _GEN_10497 : _GEN_10337; // @[executor.scala 308:60]
  wire [7:0] _GEN_10658 = 8'h7 < length_3 ? _GEN_10498 : _GEN_10338; // @[executor.scala 308:60]
  wire [7:0] _GEN_10659 = 8'h7 < length_3 ? _GEN_10499 : _GEN_10339; // @[executor.scala 308:60]
  wire [7:0] _GEN_10660 = 8'h7 < length_3 ? _GEN_10500 : _GEN_10340; // @[executor.scala 308:60]
  wire [7:0] _GEN_10661 = 8'h7 < length_3 ? _GEN_10501 : _GEN_10341; // @[executor.scala 308:60]
  wire [7:0] _GEN_10662 = 8'h7 < length_3 ? _GEN_10502 : _GEN_10342; // @[executor.scala 308:60]
  wire [7:0] _GEN_10663 = 8'h7 < length_3 ? _GEN_10503 : _GEN_10343; // @[executor.scala 308:60]
  wire [7:0] _GEN_10664 = 8'h7 < length_3 ? _GEN_10504 : _GEN_10344; // @[executor.scala 308:60]
  wire [7:0] _GEN_10665 = 8'h7 < length_3 ? _GEN_10505 : _GEN_10345; // @[executor.scala 308:60]
  wire [7:0] _GEN_10666 = 8'h7 < length_3 ? _GEN_10506 : _GEN_10346; // @[executor.scala 308:60]
  wire [7:0] _GEN_10667 = 8'h7 < length_3 ? _GEN_10507 : _GEN_10347; // @[executor.scala 308:60]
  wire [7:0] _GEN_10668 = 8'h7 < length_3 ? _GEN_10508 : _GEN_10348; // @[executor.scala 308:60]
  wire [7:0] _GEN_10669 = 8'h7 < length_3 ? _GEN_10509 : _GEN_10349; // @[executor.scala 308:60]
  wire [7:0] _GEN_10670 = 8'h7 < length_3 ? _GEN_10510 : _GEN_10350; // @[executor.scala 308:60]
  wire [7:0] _GEN_10671 = 8'h7 < length_3 ? _GEN_10511 : _GEN_10351; // @[executor.scala 308:60]
  wire [7:0] _GEN_10672 = 8'h7 < length_3 ? _GEN_10512 : _GEN_10352; // @[executor.scala 308:60]
  wire [7:0] _GEN_10673 = 8'h7 < length_3 ? _GEN_10513 : _GEN_10353; // @[executor.scala 308:60]
  wire [7:0] _GEN_10674 = 8'h7 < length_3 ? _GEN_10514 : _GEN_10354; // @[executor.scala 308:60]
  wire [7:0] _GEN_10675 = 8'h7 < length_3 ? _GEN_10515 : _GEN_10355; // @[executor.scala 308:60]
  wire [7:0] _GEN_10676 = 8'h7 < length_3 ? _GEN_10516 : _GEN_10356; // @[executor.scala 308:60]
  wire [7:0] _GEN_10677 = 8'h7 < length_3 ? _GEN_10517 : _GEN_10357; // @[executor.scala 308:60]
  wire [7:0] _GEN_10678 = 8'h7 < length_3 ? _GEN_10518 : _GEN_10358; // @[executor.scala 308:60]
  wire [7:0] _GEN_10679 = 8'h7 < length_3 ? _GEN_10519 : _GEN_10359; // @[executor.scala 308:60]
  wire [7:0] _GEN_10680 = 8'h7 < length_3 ? _GEN_10520 : _GEN_10360; // @[executor.scala 308:60]
  wire [7:0] _GEN_10681 = 8'h7 < length_3 ? _GEN_10521 : _GEN_10361; // @[executor.scala 308:60]
  wire [7:0] _GEN_10682 = 8'h7 < length_3 ? _GEN_10522 : _GEN_10362; // @[executor.scala 308:60]
  wire [7:0] _GEN_10683 = 8'h7 < length_3 ? _GEN_10523 : _GEN_10363; // @[executor.scala 308:60]
  wire [7:0] _GEN_10684 = 8'h7 < length_3 ? _GEN_10524 : _GEN_10364; // @[executor.scala 308:60]
  wire [7:0] _GEN_10685 = 8'h7 < length_3 ? _GEN_10525 : _GEN_10365; // @[executor.scala 308:60]
  wire [7:0] _GEN_10686 = 8'h7 < length_3 ? _GEN_10526 : _GEN_10366; // @[executor.scala 308:60]
  wire [7:0] _GEN_10687 = 8'h7 < length_3 ? _GEN_10527 : _GEN_10367; // @[executor.scala 308:60]
  wire [7:0] _GEN_10688 = 8'h7 < length_3 ? _GEN_10528 : _GEN_10368; // @[executor.scala 308:60]
  wire [7:0] _GEN_10689 = 8'h7 < length_3 ? _GEN_10529 : _GEN_10369; // @[executor.scala 308:60]
  wire [7:0] _GEN_10690 = 8'h7 < length_3 ? _GEN_10530 : _GEN_10370; // @[executor.scala 308:60]
  wire [7:0] _GEN_10691 = 8'h7 < length_3 ? _GEN_10531 : _GEN_10371; // @[executor.scala 308:60]
  wire [7:0] _GEN_10692 = 8'h7 < length_3 ? _GEN_10532 : _GEN_10372; // @[executor.scala 308:60]
  wire [7:0] _GEN_10693 = 8'h7 < length_3 ? _GEN_10533 : _GEN_10373; // @[executor.scala 308:60]
  wire [7:0] _GEN_10694 = 8'h7 < length_3 ? _GEN_10534 : _GEN_10374; // @[executor.scala 308:60]
  wire [7:0] _GEN_10695 = 8'h7 < length_3 ? _GEN_10535 : _GEN_10375; // @[executor.scala 308:60]
  wire [7:0] _GEN_10696 = 8'h7 < length_3 ? _GEN_10536 : _GEN_10376; // @[executor.scala 308:60]
  wire [7:0] _GEN_10697 = 8'h7 < length_3 ? _GEN_10537 : _GEN_10377; // @[executor.scala 308:60]
  wire [7:0] _GEN_10698 = 8'h7 < length_3 ? _GEN_10538 : _GEN_10378; // @[executor.scala 308:60]
  wire [7:0] _GEN_10699 = 8'h7 < length_3 ? _GEN_10539 : _GEN_10379; // @[executor.scala 308:60]
  wire [7:0] _GEN_10700 = 8'h7 < length_3 ? _GEN_10540 : _GEN_10380; // @[executor.scala 308:60]
  wire [7:0] _GEN_10701 = 8'h7 < length_3 ? _GEN_10541 : _GEN_10381; // @[executor.scala 308:60]
  wire [7:0] _GEN_10702 = 8'h7 < length_3 ? _GEN_10542 : _GEN_10382; // @[executor.scala 308:60]
  wire [7:0] _GEN_10703 = 8'h7 < length_3 ? _GEN_10543 : _GEN_10383; // @[executor.scala 308:60]
  wire [7:0] _GEN_10704 = 8'h7 < length_3 ? _GEN_10544 : _GEN_10384; // @[executor.scala 308:60]
  wire [7:0] _GEN_10705 = 8'h7 < length_3 ? _GEN_10545 : _GEN_10385; // @[executor.scala 308:60]
  wire [7:0] _GEN_10706 = 8'h7 < length_3 ? _GEN_10546 : _GEN_10386; // @[executor.scala 308:60]
  wire [7:0] _GEN_10707 = 8'h7 < length_3 ? _GEN_10547 : _GEN_10387; // @[executor.scala 308:60]
  wire [7:0] _GEN_10708 = 8'h7 < length_3 ? _GEN_10548 : _GEN_10388; // @[executor.scala 308:60]
  wire [7:0] _GEN_10709 = 8'h7 < length_3 ? _GEN_10549 : _GEN_10389; // @[executor.scala 308:60]
  wire [7:0] _GEN_10710 = 8'h7 < length_3 ? _GEN_10550 : _GEN_10390; // @[executor.scala 308:60]
  wire [7:0] _GEN_10711 = 8'h7 < length_3 ? _GEN_10551 : _GEN_10391; // @[executor.scala 308:60]
  wire [7:0] _GEN_10712 = 8'h7 < length_3 ? _GEN_10552 : _GEN_10392; // @[executor.scala 308:60]
  wire [7:0] _GEN_10713 = 8'h7 < length_3 ? _GEN_10553 : _GEN_10393; // @[executor.scala 308:60]
  wire [7:0] _GEN_10714 = 8'h7 < length_3 ? _GEN_10554 : _GEN_10394; // @[executor.scala 308:60]
  wire [7:0] _GEN_10715 = 8'h7 < length_3 ? _GEN_10555 : _GEN_10395; // @[executor.scala 308:60]
  wire [7:0] _GEN_10716 = 8'h7 < length_3 ? _GEN_10556 : _GEN_10396; // @[executor.scala 308:60]
  wire [7:0] _GEN_10717 = 8'h7 < length_3 ? _GEN_10557 : _GEN_10397; // @[executor.scala 308:60]
  wire [7:0] _GEN_10718 = 8'h7 < length_3 ? _GEN_10558 : _GEN_10398; // @[executor.scala 308:60]
  wire [7:0] _GEN_10719 = 8'h7 < length_3 ? _GEN_10559 : _GEN_10399; // @[executor.scala 308:60]
  wire [7:0] _GEN_10720 = 8'h7 < length_3 ? _GEN_10560 : _GEN_10400; // @[executor.scala 308:60]
  wire [7:0] _GEN_10721 = 8'h7 < length_3 ? _GEN_10561 : _GEN_10401; // @[executor.scala 308:60]
  wire [7:0] _GEN_10722 = 8'h7 < length_3 ? _GEN_10562 : _GEN_10402; // @[executor.scala 308:60]
  wire [7:0] _GEN_10723 = 8'h7 < length_3 ? _GEN_10563 : _GEN_10403; // @[executor.scala 308:60]
  wire [7:0] _GEN_10724 = 8'h7 < length_3 ? _GEN_10564 : _GEN_10404; // @[executor.scala 308:60]
  wire [7:0] _GEN_10725 = 8'h7 < length_3 ? _GEN_10565 : _GEN_10405; // @[executor.scala 308:60]
  wire [3:0] _GEN_10726 = length_3 == 8'h0 ? field_3[13:10] : _GEN_8004; // @[executor.scala 300:71 executor.scala 301:55]
  wire  _GEN_10727 = length_3 == 8'h0 ? field_3[0] : _GEN_8005; // @[executor.scala 300:71 executor.scala 302:55]
  wire [7:0] _GEN_10728 = length_3 == 8'h0 ? _GEN_8006 : _GEN_10566; // @[executor.scala 300:71]
  wire [7:0] _GEN_10729 = length_3 == 8'h0 ? _GEN_8007 : _GEN_10567; // @[executor.scala 300:71]
  wire [7:0] _GEN_10730 = length_3 == 8'h0 ? _GEN_8008 : _GEN_10568; // @[executor.scala 300:71]
  wire [7:0] _GEN_10731 = length_3 == 8'h0 ? _GEN_8009 : _GEN_10569; // @[executor.scala 300:71]
  wire [7:0] _GEN_10732 = length_3 == 8'h0 ? _GEN_8010 : _GEN_10570; // @[executor.scala 300:71]
  wire [7:0] _GEN_10733 = length_3 == 8'h0 ? _GEN_8011 : _GEN_10571; // @[executor.scala 300:71]
  wire [7:0] _GEN_10734 = length_3 == 8'h0 ? _GEN_8012 : _GEN_10572; // @[executor.scala 300:71]
  wire [7:0] _GEN_10735 = length_3 == 8'h0 ? _GEN_8013 : _GEN_10573; // @[executor.scala 300:71]
  wire [7:0] _GEN_10736 = length_3 == 8'h0 ? _GEN_8014 : _GEN_10574; // @[executor.scala 300:71]
  wire [7:0] _GEN_10737 = length_3 == 8'h0 ? _GEN_8015 : _GEN_10575; // @[executor.scala 300:71]
  wire [7:0] _GEN_10738 = length_3 == 8'h0 ? _GEN_8016 : _GEN_10576; // @[executor.scala 300:71]
  wire [7:0] _GEN_10739 = length_3 == 8'h0 ? _GEN_8017 : _GEN_10577; // @[executor.scala 300:71]
  wire [7:0] _GEN_10740 = length_3 == 8'h0 ? _GEN_8018 : _GEN_10578; // @[executor.scala 300:71]
  wire [7:0] _GEN_10741 = length_3 == 8'h0 ? _GEN_8019 : _GEN_10579; // @[executor.scala 300:71]
  wire [7:0] _GEN_10742 = length_3 == 8'h0 ? _GEN_8020 : _GEN_10580; // @[executor.scala 300:71]
  wire [7:0] _GEN_10743 = length_3 == 8'h0 ? _GEN_8021 : _GEN_10581; // @[executor.scala 300:71]
  wire [7:0] _GEN_10744 = length_3 == 8'h0 ? _GEN_8022 : _GEN_10582; // @[executor.scala 300:71]
  wire [7:0] _GEN_10745 = length_3 == 8'h0 ? _GEN_8023 : _GEN_10583; // @[executor.scala 300:71]
  wire [7:0] _GEN_10746 = length_3 == 8'h0 ? _GEN_8024 : _GEN_10584; // @[executor.scala 300:71]
  wire [7:0] _GEN_10747 = length_3 == 8'h0 ? _GEN_8025 : _GEN_10585; // @[executor.scala 300:71]
  wire [7:0] _GEN_10748 = length_3 == 8'h0 ? _GEN_8026 : _GEN_10586; // @[executor.scala 300:71]
  wire [7:0] _GEN_10749 = length_3 == 8'h0 ? _GEN_8027 : _GEN_10587; // @[executor.scala 300:71]
  wire [7:0] _GEN_10750 = length_3 == 8'h0 ? _GEN_8028 : _GEN_10588; // @[executor.scala 300:71]
  wire [7:0] _GEN_10751 = length_3 == 8'h0 ? _GEN_8029 : _GEN_10589; // @[executor.scala 300:71]
  wire [7:0] _GEN_10752 = length_3 == 8'h0 ? _GEN_8030 : _GEN_10590; // @[executor.scala 300:71]
  wire [7:0] _GEN_10753 = length_3 == 8'h0 ? _GEN_8031 : _GEN_10591; // @[executor.scala 300:71]
  wire [7:0] _GEN_10754 = length_3 == 8'h0 ? _GEN_8032 : _GEN_10592; // @[executor.scala 300:71]
  wire [7:0] _GEN_10755 = length_3 == 8'h0 ? _GEN_8033 : _GEN_10593; // @[executor.scala 300:71]
  wire [7:0] _GEN_10756 = length_3 == 8'h0 ? _GEN_8034 : _GEN_10594; // @[executor.scala 300:71]
  wire [7:0] _GEN_10757 = length_3 == 8'h0 ? _GEN_8035 : _GEN_10595; // @[executor.scala 300:71]
  wire [7:0] _GEN_10758 = length_3 == 8'h0 ? _GEN_8036 : _GEN_10596; // @[executor.scala 300:71]
  wire [7:0] _GEN_10759 = length_3 == 8'h0 ? _GEN_8037 : _GEN_10597; // @[executor.scala 300:71]
  wire [7:0] _GEN_10760 = length_3 == 8'h0 ? _GEN_8038 : _GEN_10598; // @[executor.scala 300:71]
  wire [7:0] _GEN_10761 = length_3 == 8'h0 ? _GEN_8039 : _GEN_10599; // @[executor.scala 300:71]
  wire [7:0] _GEN_10762 = length_3 == 8'h0 ? _GEN_8040 : _GEN_10600; // @[executor.scala 300:71]
  wire [7:0] _GEN_10763 = length_3 == 8'h0 ? _GEN_8041 : _GEN_10601; // @[executor.scala 300:71]
  wire [7:0] _GEN_10764 = length_3 == 8'h0 ? _GEN_8042 : _GEN_10602; // @[executor.scala 300:71]
  wire [7:0] _GEN_10765 = length_3 == 8'h0 ? _GEN_8043 : _GEN_10603; // @[executor.scala 300:71]
  wire [7:0] _GEN_10766 = length_3 == 8'h0 ? _GEN_8044 : _GEN_10604; // @[executor.scala 300:71]
  wire [7:0] _GEN_10767 = length_3 == 8'h0 ? _GEN_8045 : _GEN_10605; // @[executor.scala 300:71]
  wire [7:0] _GEN_10768 = length_3 == 8'h0 ? _GEN_8046 : _GEN_10606; // @[executor.scala 300:71]
  wire [7:0] _GEN_10769 = length_3 == 8'h0 ? _GEN_8047 : _GEN_10607; // @[executor.scala 300:71]
  wire [7:0] _GEN_10770 = length_3 == 8'h0 ? _GEN_8048 : _GEN_10608; // @[executor.scala 300:71]
  wire [7:0] _GEN_10771 = length_3 == 8'h0 ? _GEN_8049 : _GEN_10609; // @[executor.scala 300:71]
  wire [7:0] _GEN_10772 = length_3 == 8'h0 ? _GEN_8050 : _GEN_10610; // @[executor.scala 300:71]
  wire [7:0] _GEN_10773 = length_3 == 8'h0 ? _GEN_8051 : _GEN_10611; // @[executor.scala 300:71]
  wire [7:0] _GEN_10774 = length_3 == 8'h0 ? _GEN_8052 : _GEN_10612; // @[executor.scala 300:71]
  wire [7:0] _GEN_10775 = length_3 == 8'h0 ? _GEN_8053 : _GEN_10613; // @[executor.scala 300:71]
  wire [7:0] _GEN_10776 = length_3 == 8'h0 ? _GEN_8054 : _GEN_10614; // @[executor.scala 300:71]
  wire [7:0] _GEN_10777 = length_3 == 8'h0 ? _GEN_8055 : _GEN_10615; // @[executor.scala 300:71]
  wire [7:0] _GEN_10778 = length_3 == 8'h0 ? _GEN_8056 : _GEN_10616; // @[executor.scala 300:71]
  wire [7:0] _GEN_10779 = length_3 == 8'h0 ? _GEN_8057 : _GEN_10617; // @[executor.scala 300:71]
  wire [7:0] _GEN_10780 = length_3 == 8'h0 ? _GEN_8058 : _GEN_10618; // @[executor.scala 300:71]
  wire [7:0] _GEN_10781 = length_3 == 8'h0 ? _GEN_8059 : _GEN_10619; // @[executor.scala 300:71]
  wire [7:0] _GEN_10782 = length_3 == 8'h0 ? _GEN_8060 : _GEN_10620; // @[executor.scala 300:71]
  wire [7:0] _GEN_10783 = length_3 == 8'h0 ? _GEN_8061 : _GEN_10621; // @[executor.scala 300:71]
  wire [7:0] _GEN_10784 = length_3 == 8'h0 ? _GEN_8062 : _GEN_10622; // @[executor.scala 300:71]
  wire [7:0] _GEN_10785 = length_3 == 8'h0 ? _GEN_8063 : _GEN_10623; // @[executor.scala 300:71]
  wire [7:0] _GEN_10786 = length_3 == 8'h0 ? _GEN_8064 : _GEN_10624; // @[executor.scala 300:71]
  wire [7:0] _GEN_10787 = length_3 == 8'h0 ? _GEN_8065 : _GEN_10625; // @[executor.scala 300:71]
  wire [7:0] _GEN_10788 = length_3 == 8'h0 ? _GEN_8066 : _GEN_10626; // @[executor.scala 300:71]
  wire [7:0] _GEN_10789 = length_3 == 8'h0 ? _GEN_8067 : _GEN_10627; // @[executor.scala 300:71]
  wire [7:0] _GEN_10790 = length_3 == 8'h0 ? _GEN_8068 : _GEN_10628; // @[executor.scala 300:71]
  wire [7:0] _GEN_10791 = length_3 == 8'h0 ? _GEN_8069 : _GEN_10629; // @[executor.scala 300:71]
  wire [7:0] _GEN_10792 = length_3 == 8'h0 ? _GEN_8070 : _GEN_10630; // @[executor.scala 300:71]
  wire [7:0] _GEN_10793 = length_3 == 8'h0 ? _GEN_8071 : _GEN_10631; // @[executor.scala 300:71]
  wire [7:0] _GEN_10794 = length_3 == 8'h0 ? _GEN_8072 : _GEN_10632; // @[executor.scala 300:71]
  wire [7:0] _GEN_10795 = length_3 == 8'h0 ? _GEN_8073 : _GEN_10633; // @[executor.scala 300:71]
  wire [7:0] _GEN_10796 = length_3 == 8'h0 ? _GEN_8074 : _GEN_10634; // @[executor.scala 300:71]
  wire [7:0] _GEN_10797 = length_3 == 8'h0 ? _GEN_8075 : _GEN_10635; // @[executor.scala 300:71]
  wire [7:0] _GEN_10798 = length_3 == 8'h0 ? _GEN_8076 : _GEN_10636; // @[executor.scala 300:71]
  wire [7:0] _GEN_10799 = length_3 == 8'h0 ? _GEN_8077 : _GEN_10637; // @[executor.scala 300:71]
  wire [7:0] _GEN_10800 = length_3 == 8'h0 ? _GEN_8078 : _GEN_10638; // @[executor.scala 300:71]
  wire [7:0] _GEN_10801 = length_3 == 8'h0 ? _GEN_8079 : _GEN_10639; // @[executor.scala 300:71]
  wire [7:0] _GEN_10802 = length_3 == 8'h0 ? _GEN_8080 : _GEN_10640; // @[executor.scala 300:71]
  wire [7:0] _GEN_10803 = length_3 == 8'h0 ? _GEN_8081 : _GEN_10641; // @[executor.scala 300:71]
  wire [7:0] _GEN_10804 = length_3 == 8'h0 ? _GEN_8082 : _GEN_10642; // @[executor.scala 300:71]
  wire [7:0] _GEN_10805 = length_3 == 8'h0 ? _GEN_8083 : _GEN_10643; // @[executor.scala 300:71]
  wire [7:0] _GEN_10806 = length_3 == 8'h0 ? _GEN_8084 : _GEN_10644; // @[executor.scala 300:71]
  wire [7:0] _GEN_10807 = length_3 == 8'h0 ? _GEN_8085 : _GEN_10645; // @[executor.scala 300:71]
  wire [7:0] _GEN_10808 = length_3 == 8'h0 ? _GEN_8086 : _GEN_10646; // @[executor.scala 300:71]
  wire [7:0] _GEN_10809 = length_3 == 8'h0 ? _GEN_8087 : _GEN_10647; // @[executor.scala 300:71]
  wire [7:0] _GEN_10810 = length_3 == 8'h0 ? _GEN_8088 : _GEN_10648; // @[executor.scala 300:71]
  wire [7:0] _GEN_10811 = length_3 == 8'h0 ? _GEN_8089 : _GEN_10649; // @[executor.scala 300:71]
  wire [7:0] _GEN_10812 = length_3 == 8'h0 ? _GEN_8090 : _GEN_10650; // @[executor.scala 300:71]
  wire [7:0] _GEN_10813 = length_3 == 8'h0 ? _GEN_8091 : _GEN_10651; // @[executor.scala 300:71]
  wire [7:0] _GEN_10814 = length_3 == 8'h0 ? _GEN_8092 : _GEN_10652; // @[executor.scala 300:71]
  wire [7:0] _GEN_10815 = length_3 == 8'h0 ? _GEN_8093 : _GEN_10653; // @[executor.scala 300:71]
  wire [7:0] _GEN_10816 = length_3 == 8'h0 ? _GEN_8094 : _GEN_10654; // @[executor.scala 300:71]
  wire [7:0] _GEN_10817 = length_3 == 8'h0 ? _GEN_8095 : _GEN_10655; // @[executor.scala 300:71]
  wire [7:0] _GEN_10818 = length_3 == 8'h0 ? _GEN_8096 : _GEN_10656; // @[executor.scala 300:71]
  wire [7:0] _GEN_10819 = length_3 == 8'h0 ? _GEN_8097 : _GEN_10657; // @[executor.scala 300:71]
  wire [7:0] _GEN_10820 = length_3 == 8'h0 ? _GEN_8098 : _GEN_10658; // @[executor.scala 300:71]
  wire [7:0] _GEN_10821 = length_3 == 8'h0 ? _GEN_8099 : _GEN_10659; // @[executor.scala 300:71]
  wire [7:0] _GEN_10822 = length_3 == 8'h0 ? _GEN_8100 : _GEN_10660; // @[executor.scala 300:71]
  wire [7:0] _GEN_10823 = length_3 == 8'h0 ? _GEN_8101 : _GEN_10661; // @[executor.scala 300:71]
  wire [7:0] _GEN_10824 = length_3 == 8'h0 ? _GEN_8102 : _GEN_10662; // @[executor.scala 300:71]
  wire [7:0] _GEN_10825 = length_3 == 8'h0 ? _GEN_8103 : _GEN_10663; // @[executor.scala 300:71]
  wire [7:0] _GEN_10826 = length_3 == 8'h0 ? _GEN_8104 : _GEN_10664; // @[executor.scala 300:71]
  wire [7:0] _GEN_10827 = length_3 == 8'h0 ? _GEN_8105 : _GEN_10665; // @[executor.scala 300:71]
  wire [7:0] _GEN_10828 = length_3 == 8'h0 ? _GEN_8106 : _GEN_10666; // @[executor.scala 300:71]
  wire [7:0] _GEN_10829 = length_3 == 8'h0 ? _GEN_8107 : _GEN_10667; // @[executor.scala 300:71]
  wire [7:0] _GEN_10830 = length_3 == 8'h0 ? _GEN_8108 : _GEN_10668; // @[executor.scala 300:71]
  wire [7:0] _GEN_10831 = length_3 == 8'h0 ? _GEN_8109 : _GEN_10669; // @[executor.scala 300:71]
  wire [7:0] _GEN_10832 = length_3 == 8'h0 ? _GEN_8110 : _GEN_10670; // @[executor.scala 300:71]
  wire [7:0] _GEN_10833 = length_3 == 8'h0 ? _GEN_8111 : _GEN_10671; // @[executor.scala 300:71]
  wire [7:0] _GEN_10834 = length_3 == 8'h0 ? _GEN_8112 : _GEN_10672; // @[executor.scala 300:71]
  wire [7:0] _GEN_10835 = length_3 == 8'h0 ? _GEN_8113 : _GEN_10673; // @[executor.scala 300:71]
  wire [7:0] _GEN_10836 = length_3 == 8'h0 ? _GEN_8114 : _GEN_10674; // @[executor.scala 300:71]
  wire [7:0] _GEN_10837 = length_3 == 8'h0 ? _GEN_8115 : _GEN_10675; // @[executor.scala 300:71]
  wire [7:0] _GEN_10838 = length_3 == 8'h0 ? _GEN_8116 : _GEN_10676; // @[executor.scala 300:71]
  wire [7:0] _GEN_10839 = length_3 == 8'h0 ? _GEN_8117 : _GEN_10677; // @[executor.scala 300:71]
  wire [7:0] _GEN_10840 = length_3 == 8'h0 ? _GEN_8118 : _GEN_10678; // @[executor.scala 300:71]
  wire [7:0] _GEN_10841 = length_3 == 8'h0 ? _GEN_8119 : _GEN_10679; // @[executor.scala 300:71]
  wire [7:0] _GEN_10842 = length_3 == 8'h0 ? _GEN_8120 : _GEN_10680; // @[executor.scala 300:71]
  wire [7:0] _GEN_10843 = length_3 == 8'h0 ? _GEN_8121 : _GEN_10681; // @[executor.scala 300:71]
  wire [7:0] _GEN_10844 = length_3 == 8'h0 ? _GEN_8122 : _GEN_10682; // @[executor.scala 300:71]
  wire [7:0] _GEN_10845 = length_3 == 8'h0 ? _GEN_8123 : _GEN_10683; // @[executor.scala 300:71]
  wire [7:0] _GEN_10846 = length_3 == 8'h0 ? _GEN_8124 : _GEN_10684; // @[executor.scala 300:71]
  wire [7:0] _GEN_10847 = length_3 == 8'h0 ? _GEN_8125 : _GEN_10685; // @[executor.scala 300:71]
  wire [7:0] _GEN_10848 = length_3 == 8'h0 ? _GEN_8126 : _GEN_10686; // @[executor.scala 300:71]
  wire [7:0] _GEN_10849 = length_3 == 8'h0 ? _GEN_8127 : _GEN_10687; // @[executor.scala 300:71]
  wire [7:0] _GEN_10850 = length_3 == 8'h0 ? _GEN_8128 : _GEN_10688; // @[executor.scala 300:71]
  wire [7:0] _GEN_10851 = length_3 == 8'h0 ? _GEN_8129 : _GEN_10689; // @[executor.scala 300:71]
  wire [7:0] _GEN_10852 = length_3 == 8'h0 ? _GEN_8130 : _GEN_10690; // @[executor.scala 300:71]
  wire [7:0] _GEN_10853 = length_3 == 8'h0 ? _GEN_8131 : _GEN_10691; // @[executor.scala 300:71]
  wire [7:0] _GEN_10854 = length_3 == 8'h0 ? _GEN_8132 : _GEN_10692; // @[executor.scala 300:71]
  wire [7:0] _GEN_10855 = length_3 == 8'h0 ? _GEN_8133 : _GEN_10693; // @[executor.scala 300:71]
  wire [7:0] _GEN_10856 = length_3 == 8'h0 ? _GEN_8134 : _GEN_10694; // @[executor.scala 300:71]
  wire [7:0] _GEN_10857 = length_3 == 8'h0 ? _GEN_8135 : _GEN_10695; // @[executor.scala 300:71]
  wire [7:0] _GEN_10858 = length_3 == 8'h0 ? _GEN_8136 : _GEN_10696; // @[executor.scala 300:71]
  wire [7:0] _GEN_10859 = length_3 == 8'h0 ? _GEN_8137 : _GEN_10697; // @[executor.scala 300:71]
  wire [7:0] _GEN_10860 = length_3 == 8'h0 ? _GEN_8138 : _GEN_10698; // @[executor.scala 300:71]
  wire [7:0] _GEN_10861 = length_3 == 8'h0 ? _GEN_8139 : _GEN_10699; // @[executor.scala 300:71]
  wire [7:0] _GEN_10862 = length_3 == 8'h0 ? _GEN_8140 : _GEN_10700; // @[executor.scala 300:71]
  wire [7:0] _GEN_10863 = length_3 == 8'h0 ? _GEN_8141 : _GEN_10701; // @[executor.scala 300:71]
  wire [7:0] _GEN_10864 = length_3 == 8'h0 ? _GEN_8142 : _GEN_10702; // @[executor.scala 300:71]
  wire [7:0] _GEN_10865 = length_3 == 8'h0 ? _GEN_8143 : _GEN_10703; // @[executor.scala 300:71]
  wire [7:0] _GEN_10866 = length_3 == 8'h0 ? _GEN_8144 : _GEN_10704; // @[executor.scala 300:71]
  wire [7:0] _GEN_10867 = length_3 == 8'h0 ? _GEN_8145 : _GEN_10705; // @[executor.scala 300:71]
  wire [7:0] _GEN_10868 = length_3 == 8'h0 ? _GEN_8146 : _GEN_10706; // @[executor.scala 300:71]
  wire [7:0] _GEN_10869 = length_3 == 8'h0 ? _GEN_8147 : _GEN_10707; // @[executor.scala 300:71]
  wire [7:0] _GEN_10870 = length_3 == 8'h0 ? _GEN_8148 : _GEN_10708; // @[executor.scala 300:71]
  wire [7:0] _GEN_10871 = length_3 == 8'h0 ? _GEN_8149 : _GEN_10709; // @[executor.scala 300:71]
  wire [7:0] _GEN_10872 = length_3 == 8'h0 ? _GEN_8150 : _GEN_10710; // @[executor.scala 300:71]
  wire [7:0] _GEN_10873 = length_3 == 8'h0 ? _GEN_8151 : _GEN_10711; // @[executor.scala 300:71]
  wire [7:0] _GEN_10874 = length_3 == 8'h0 ? _GEN_8152 : _GEN_10712; // @[executor.scala 300:71]
  wire [7:0] _GEN_10875 = length_3 == 8'h0 ? _GEN_8153 : _GEN_10713; // @[executor.scala 300:71]
  wire [7:0] _GEN_10876 = length_3 == 8'h0 ? _GEN_8154 : _GEN_10714; // @[executor.scala 300:71]
  wire [7:0] _GEN_10877 = length_3 == 8'h0 ? _GEN_8155 : _GEN_10715; // @[executor.scala 300:71]
  wire [7:0] _GEN_10878 = length_3 == 8'h0 ? _GEN_8156 : _GEN_10716; // @[executor.scala 300:71]
  wire [7:0] _GEN_10879 = length_3 == 8'h0 ? _GEN_8157 : _GEN_10717; // @[executor.scala 300:71]
  wire [7:0] _GEN_10880 = length_3 == 8'h0 ? _GEN_8158 : _GEN_10718; // @[executor.scala 300:71]
  wire [7:0] _GEN_10881 = length_3 == 8'h0 ? _GEN_8159 : _GEN_10719; // @[executor.scala 300:71]
  wire [7:0] _GEN_10882 = length_3 == 8'h0 ? _GEN_8160 : _GEN_10720; // @[executor.scala 300:71]
  wire [7:0] _GEN_10883 = length_3 == 8'h0 ? _GEN_8161 : _GEN_10721; // @[executor.scala 300:71]
  wire [7:0] _GEN_10884 = length_3 == 8'h0 ? _GEN_8162 : _GEN_10722; // @[executor.scala 300:71]
  wire [7:0] _GEN_10885 = length_3 == 8'h0 ? _GEN_8163 : _GEN_10723; // @[executor.scala 300:71]
  wire [7:0] _GEN_10886 = length_3 == 8'h0 ? _GEN_8164 : _GEN_10724; // @[executor.scala 300:71]
  wire [7:0] _GEN_10887 = length_3 == 8'h0 ? _GEN_8165 : _GEN_10725; // @[executor.scala 300:71]
  assign io_pipe_phv_out_data_0 = phv_is_valid_processor ? _GEN_10728 : phv_data_0; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_1 = phv_is_valid_processor ? _GEN_10729 : phv_data_1; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_2 = phv_is_valid_processor ? _GEN_10730 : phv_data_2; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_3 = phv_is_valid_processor ? _GEN_10731 : phv_data_3; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_4 = phv_is_valid_processor ? _GEN_10732 : phv_data_4; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_5 = phv_is_valid_processor ? _GEN_10733 : phv_data_5; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_6 = phv_is_valid_processor ? _GEN_10734 : phv_data_6; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_7 = phv_is_valid_processor ? _GEN_10735 : phv_data_7; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_8 = phv_is_valid_processor ? _GEN_10736 : phv_data_8; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_9 = phv_is_valid_processor ? _GEN_10737 : phv_data_9; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_10 = phv_is_valid_processor ? _GEN_10738 : phv_data_10; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_11 = phv_is_valid_processor ? _GEN_10739 : phv_data_11; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_12 = phv_is_valid_processor ? _GEN_10740 : phv_data_12; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_13 = phv_is_valid_processor ? _GEN_10741 : phv_data_13; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_14 = phv_is_valid_processor ? _GEN_10742 : phv_data_14; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_15 = phv_is_valid_processor ? _GEN_10743 : phv_data_15; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_16 = phv_is_valid_processor ? _GEN_10744 : phv_data_16; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_17 = phv_is_valid_processor ? _GEN_10745 : phv_data_17; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_18 = phv_is_valid_processor ? _GEN_10746 : phv_data_18; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_19 = phv_is_valid_processor ? _GEN_10747 : phv_data_19; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_20 = phv_is_valid_processor ? _GEN_10748 : phv_data_20; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_21 = phv_is_valid_processor ? _GEN_10749 : phv_data_21; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_22 = phv_is_valid_processor ? _GEN_10750 : phv_data_22; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_23 = phv_is_valid_processor ? _GEN_10751 : phv_data_23; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_24 = phv_is_valid_processor ? _GEN_10752 : phv_data_24; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_25 = phv_is_valid_processor ? _GEN_10753 : phv_data_25; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_26 = phv_is_valid_processor ? _GEN_10754 : phv_data_26; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_27 = phv_is_valid_processor ? _GEN_10755 : phv_data_27; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_28 = phv_is_valid_processor ? _GEN_10756 : phv_data_28; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_29 = phv_is_valid_processor ? _GEN_10757 : phv_data_29; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_30 = phv_is_valid_processor ? _GEN_10758 : phv_data_30; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_31 = phv_is_valid_processor ? _GEN_10759 : phv_data_31; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_32 = phv_is_valid_processor ? _GEN_10760 : phv_data_32; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_33 = phv_is_valid_processor ? _GEN_10761 : phv_data_33; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_34 = phv_is_valid_processor ? _GEN_10762 : phv_data_34; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_35 = phv_is_valid_processor ? _GEN_10763 : phv_data_35; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_36 = phv_is_valid_processor ? _GEN_10764 : phv_data_36; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_37 = phv_is_valid_processor ? _GEN_10765 : phv_data_37; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_38 = phv_is_valid_processor ? _GEN_10766 : phv_data_38; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_39 = phv_is_valid_processor ? _GEN_10767 : phv_data_39; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_40 = phv_is_valid_processor ? _GEN_10768 : phv_data_40; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_41 = phv_is_valid_processor ? _GEN_10769 : phv_data_41; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_42 = phv_is_valid_processor ? _GEN_10770 : phv_data_42; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_43 = phv_is_valid_processor ? _GEN_10771 : phv_data_43; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_44 = phv_is_valid_processor ? _GEN_10772 : phv_data_44; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_45 = phv_is_valid_processor ? _GEN_10773 : phv_data_45; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_46 = phv_is_valid_processor ? _GEN_10774 : phv_data_46; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_47 = phv_is_valid_processor ? _GEN_10775 : phv_data_47; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_48 = phv_is_valid_processor ? _GEN_10776 : phv_data_48; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_49 = phv_is_valid_processor ? _GEN_10777 : phv_data_49; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_50 = phv_is_valid_processor ? _GEN_10778 : phv_data_50; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_51 = phv_is_valid_processor ? _GEN_10779 : phv_data_51; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_52 = phv_is_valid_processor ? _GEN_10780 : phv_data_52; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_53 = phv_is_valid_processor ? _GEN_10781 : phv_data_53; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_54 = phv_is_valid_processor ? _GEN_10782 : phv_data_54; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_55 = phv_is_valid_processor ? _GEN_10783 : phv_data_55; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_56 = phv_is_valid_processor ? _GEN_10784 : phv_data_56; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_57 = phv_is_valid_processor ? _GEN_10785 : phv_data_57; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_58 = phv_is_valid_processor ? _GEN_10786 : phv_data_58; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_59 = phv_is_valid_processor ? _GEN_10787 : phv_data_59; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_60 = phv_is_valid_processor ? _GEN_10788 : phv_data_60; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_61 = phv_is_valid_processor ? _GEN_10789 : phv_data_61; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_62 = phv_is_valid_processor ? _GEN_10790 : phv_data_62; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_63 = phv_is_valid_processor ? _GEN_10791 : phv_data_63; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_64 = phv_is_valid_processor ? _GEN_10792 : phv_data_64; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_65 = phv_is_valid_processor ? _GEN_10793 : phv_data_65; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_66 = phv_is_valid_processor ? _GEN_10794 : phv_data_66; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_67 = phv_is_valid_processor ? _GEN_10795 : phv_data_67; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_68 = phv_is_valid_processor ? _GEN_10796 : phv_data_68; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_69 = phv_is_valid_processor ? _GEN_10797 : phv_data_69; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_70 = phv_is_valid_processor ? _GEN_10798 : phv_data_70; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_71 = phv_is_valid_processor ? _GEN_10799 : phv_data_71; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_72 = phv_is_valid_processor ? _GEN_10800 : phv_data_72; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_73 = phv_is_valid_processor ? _GEN_10801 : phv_data_73; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_74 = phv_is_valid_processor ? _GEN_10802 : phv_data_74; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_75 = phv_is_valid_processor ? _GEN_10803 : phv_data_75; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_76 = phv_is_valid_processor ? _GEN_10804 : phv_data_76; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_77 = phv_is_valid_processor ? _GEN_10805 : phv_data_77; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_78 = phv_is_valid_processor ? _GEN_10806 : phv_data_78; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_79 = phv_is_valid_processor ? _GEN_10807 : phv_data_79; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_80 = phv_is_valid_processor ? _GEN_10808 : phv_data_80; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_81 = phv_is_valid_processor ? _GEN_10809 : phv_data_81; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_82 = phv_is_valid_processor ? _GEN_10810 : phv_data_82; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_83 = phv_is_valid_processor ? _GEN_10811 : phv_data_83; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_84 = phv_is_valid_processor ? _GEN_10812 : phv_data_84; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_85 = phv_is_valid_processor ? _GEN_10813 : phv_data_85; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_86 = phv_is_valid_processor ? _GEN_10814 : phv_data_86; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_87 = phv_is_valid_processor ? _GEN_10815 : phv_data_87; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_88 = phv_is_valid_processor ? _GEN_10816 : phv_data_88; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_89 = phv_is_valid_processor ? _GEN_10817 : phv_data_89; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_90 = phv_is_valid_processor ? _GEN_10818 : phv_data_90; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_91 = phv_is_valid_processor ? _GEN_10819 : phv_data_91; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_92 = phv_is_valid_processor ? _GEN_10820 : phv_data_92; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_93 = phv_is_valid_processor ? _GEN_10821 : phv_data_93; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_94 = phv_is_valid_processor ? _GEN_10822 : phv_data_94; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_95 = phv_is_valid_processor ? _GEN_10823 : phv_data_95; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_96 = phv_is_valid_processor ? _GEN_10824 : phv_data_96; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_97 = phv_is_valid_processor ? _GEN_10825 : phv_data_97; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_98 = phv_is_valid_processor ? _GEN_10826 : phv_data_98; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_99 = phv_is_valid_processor ? _GEN_10827 : phv_data_99; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_100 = phv_is_valid_processor ? _GEN_10828 : phv_data_100; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_101 = phv_is_valid_processor ? _GEN_10829 : phv_data_101; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_102 = phv_is_valid_processor ? _GEN_10830 : phv_data_102; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_103 = phv_is_valid_processor ? _GEN_10831 : phv_data_103; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_104 = phv_is_valid_processor ? _GEN_10832 : phv_data_104; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_105 = phv_is_valid_processor ? _GEN_10833 : phv_data_105; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_106 = phv_is_valid_processor ? _GEN_10834 : phv_data_106; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_107 = phv_is_valid_processor ? _GEN_10835 : phv_data_107; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_108 = phv_is_valid_processor ? _GEN_10836 : phv_data_108; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_109 = phv_is_valid_processor ? _GEN_10837 : phv_data_109; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_110 = phv_is_valid_processor ? _GEN_10838 : phv_data_110; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_111 = phv_is_valid_processor ? _GEN_10839 : phv_data_111; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_112 = phv_is_valid_processor ? _GEN_10840 : phv_data_112; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_113 = phv_is_valid_processor ? _GEN_10841 : phv_data_113; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_114 = phv_is_valid_processor ? _GEN_10842 : phv_data_114; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_115 = phv_is_valid_processor ? _GEN_10843 : phv_data_115; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_116 = phv_is_valid_processor ? _GEN_10844 : phv_data_116; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_117 = phv_is_valid_processor ? _GEN_10845 : phv_data_117; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_118 = phv_is_valid_processor ? _GEN_10846 : phv_data_118; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_119 = phv_is_valid_processor ? _GEN_10847 : phv_data_119; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_120 = phv_is_valid_processor ? _GEN_10848 : phv_data_120; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_121 = phv_is_valid_processor ? _GEN_10849 : phv_data_121; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_122 = phv_is_valid_processor ? _GEN_10850 : phv_data_122; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_123 = phv_is_valid_processor ? _GEN_10851 : phv_data_123; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_124 = phv_is_valid_processor ? _GEN_10852 : phv_data_124; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_125 = phv_is_valid_processor ? _GEN_10853 : phv_data_125; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_126 = phv_is_valid_processor ? _GEN_10854 : phv_data_126; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_127 = phv_is_valid_processor ? _GEN_10855 : phv_data_127; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_128 = phv_is_valid_processor ? _GEN_10856 : phv_data_128; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_129 = phv_is_valid_processor ? _GEN_10857 : phv_data_129; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_130 = phv_is_valid_processor ? _GEN_10858 : phv_data_130; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_131 = phv_is_valid_processor ? _GEN_10859 : phv_data_131; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_132 = phv_is_valid_processor ? _GEN_10860 : phv_data_132; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_133 = phv_is_valid_processor ? _GEN_10861 : phv_data_133; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_134 = phv_is_valid_processor ? _GEN_10862 : phv_data_134; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_135 = phv_is_valid_processor ? _GEN_10863 : phv_data_135; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_136 = phv_is_valid_processor ? _GEN_10864 : phv_data_136; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_137 = phv_is_valid_processor ? _GEN_10865 : phv_data_137; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_138 = phv_is_valid_processor ? _GEN_10866 : phv_data_138; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_139 = phv_is_valid_processor ? _GEN_10867 : phv_data_139; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_140 = phv_is_valid_processor ? _GEN_10868 : phv_data_140; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_141 = phv_is_valid_processor ? _GEN_10869 : phv_data_141; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_142 = phv_is_valid_processor ? _GEN_10870 : phv_data_142; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_143 = phv_is_valid_processor ? _GEN_10871 : phv_data_143; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_144 = phv_is_valid_processor ? _GEN_10872 : phv_data_144; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_145 = phv_is_valid_processor ? _GEN_10873 : phv_data_145; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_146 = phv_is_valid_processor ? _GEN_10874 : phv_data_146; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_147 = phv_is_valid_processor ? _GEN_10875 : phv_data_147; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_148 = phv_is_valid_processor ? _GEN_10876 : phv_data_148; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_149 = phv_is_valid_processor ? _GEN_10877 : phv_data_149; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_150 = phv_is_valid_processor ? _GEN_10878 : phv_data_150; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_151 = phv_is_valid_processor ? _GEN_10879 : phv_data_151; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_152 = phv_is_valid_processor ? _GEN_10880 : phv_data_152; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_153 = phv_is_valid_processor ? _GEN_10881 : phv_data_153; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_154 = phv_is_valid_processor ? _GEN_10882 : phv_data_154; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_155 = phv_is_valid_processor ? _GEN_10883 : phv_data_155; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_156 = phv_is_valid_processor ? _GEN_10884 : phv_data_156; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_157 = phv_is_valid_processor ? _GEN_10885 : phv_data_157; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_158 = phv_is_valid_processor ? _GEN_10886 : phv_data_158; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_data_159 = phv_is_valid_processor ? _GEN_10887 : phv_data_159; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_header_0 = phv_header_0; // @[executor.scala 286:25]
  assign io_pipe_phv_out_header_1 = phv_header_1; // @[executor.scala 286:25]
  assign io_pipe_phv_out_header_2 = phv_header_2; // @[executor.scala 286:25]
  assign io_pipe_phv_out_header_3 = phv_header_3; // @[executor.scala 286:25]
  assign io_pipe_phv_out_header_4 = phv_header_4; // @[executor.scala 286:25]
  assign io_pipe_phv_out_header_5 = phv_header_5; // @[executor.scala 286:25]
  assign io_pipe_phv_out_header_6 = phv_header_6; // @[executor.scala 286:25]
  assign io_pipe_phv_out_header_7 = phv_header_7; // @[executor.scala 286:25]
  assign io_pipe_phv_out_header_8 = phv_header_8; // @[executor.scala 286:25]
  assign io_pipe_phv_out_header_9 = phv_header_9; // @[executor.scala 286:25]
  assign io_pipe_phv_out_header_10 = phv_header_10; // @[executor.scala 286:25]
  assign io_pipe_phv_out_header_11 = phv_header_11; // @[executor.scala 286:25]
  assign io_pipe_phv_out_header_12 = phv_header_12; // @[executor.scala 286:25]
  assign io_pipe_phv_out_header_13 = phv_header_13; // @[executor.scala 286:25]
  assign io_pipe_phv_out_header_14 = phv_header_14; // @[executor.scala 286:25]
  assign io_pipe_phv_out_header_15 = phv_header_15; // @[executor.scala 286:25]
  assign io_pipe_phv_out_parse_current_state = phv_parse_current_state; // @[executor.scala 286:25]
  assign io_pipe_phv_out_parse_current_offset = phv_parse_current_offset; // @[executor.scala 286:25]
  assign io_pipe_phv_out_parse_transition_field = phv_parse_transition_field; // @[executor.scala 286:25]
  assign io_pipe_phv_out_next_processor_id = phv_is_valid_processor ? _GEN_10726 : phv_next_processor_id; // @[executor.scala 295:39 executor.scala 286:25]
  assign io_pipe_phv_out_next_config_id = phv_is_valid_processor ? _GEN_10727 : phv_next_config_id; // @[executor.scala 295:39 executor.scala 286:25]
  always @(posedge clock) begin
    phv_data_0 <= io_pipe_phv_in_data_0; // @[executor.scala 285:13]
    phv_data_1 <= io_pipe_phv_in_data_1; // @[executor.scala 285:13]
    phv_data_2 <= io_pipe_phv_in_data_2; // @[executor.scala 285:13]
    phv_data_3 <= io_pipe_phv_in_data_3; // @[executor.scala 285:13]
    phv_data_4 <= io_pipe_phv_in_data_4; // @[executor.scala 285:13]
    phv_data_5 <= io_pipe_phv_in_data_5; // @[executor.scala 285:13]
    phv_data_6 <= io_pipe_phv_in_data_6; // @[executor.scala 285:13]
    phv_data_7 <= io_pipe_phv_in_data_7; // @[executor.scala 285:13]
    phv_data_8 <= io_pipe_phv_in_data_8; // @[executor.scala 285:13]
    phv_data_9 <= io_pipe_phv_in_data_9; // @[executor.scala 285:13]
    phv_data_10 <= io_pipe_phv_in_data_10; // @[executor.scala 285:13]
    phv_data_11 <= io_pipe_phv_in_data_11; // @[executor.scala 285:13]
    phv_data_12 <= io_pipe_phv_in_data_12; // @[executor.scala 285:13]
    phv_data_13 <= io_pipe_phv_in_data_13; // @[executor.scala 285:13]
    phv_data_14 <= io_pipe_phv_in_data_14; // @[executor.scala 285:13]
    phv_data_15 <= io_pipe_phv_in_data_15; // @[executor.scala 285:13]
    phv_data_16 <= io_pipe_phv_in_data_16; // @[executor.scala 285:13]
    phv_data_17 <= io_pipe_phv_in_data_17; // @[executor.scala 285:13]
    phv_data_18 <= io_pipe_phv_in_data_18; // @[executor.scala 285:13]
    phv_data_19 <= io_pipe_phv_in_data_19; // @[executor.scala 285:13]
    phv_data_20 <= io_pipe_phv_in_data_20; // @[executor.scala 285:13]
    phv_data_21 <= io_pipe_phv_in_data_21; // @[executor.scala 285:13]
    phv_data_22 <= io_pipe_phv_in_data_22; // @[executor.scala 285:13]
    phv_data_23 <= io_pipe_phv_in_data_23; // @[executor.scala 285:13]
    phv_data_24 <= io_pipe_phv_in_data_24; // @[executor.scala 285:13]
    phv_data_25 <= io_pipe_phv_in_data_25; // @[executor.scala 285:13]
    phv_data_26 <= io_pipe_phv_in_data_26; // @[executor.scala 285:13]
    phv_data_27 <= io_pipe_phv_in_data_27; // @[executor.scala 285:13]
    phv_data_28 <= io_pipe_phv_in_data_28; // @[executor.scala 285:13]
    phv_data_29 <= io_pipe_phv_in_data_29; // @[executor.scala 285:13]
    phv_data_30 <= io_pipe_phv_in_data_30; // @[executor.scala 285:13]
    phv_data_31 <= io_pipe_phv_in_data_31; // @[executor.scala 285:13]
    phv_data_32 <= io_pipe_phv_in_data_32; // @[executor.scala 285:13]
    phv_data_33 <= io_pipe_phv_in_data_33; // @[executor.scala 285:13]
    phv_data_34 <= io_pipe_phv_in_data_34; // @[executor.scala 285:13]
    phv_data_35 <= io_pipe_phv_in_data_35; // @[executor.scala 285:13]
    phv_data_36 <= io_pipe_phv_in_data_36; // @[executor.scala 285:13]
    phv_data_37 <= io_pipe_phv_in_data_37; // @[executor.scala 285:13]
    phv_data_38 <= io_pipe_phv_in_data_38; // @[executor.scala 285:13]
    phv_data_39 <= io_pipe_phv_in_data_39; // @[executor.scala 285:13]
    phv_data_40 <= io_pipe_phv_in_data_40; // @[executor.scala 285:13]
    phv_data_41 <= io_pipe_phv_in_data_41; // @[executor.scala 285:13]
    phv_data_42 <= io_pipe_phv_in_data_42; // @[executor.scala 285:13]
    phv_data_43 <= io_pipe_phv_in_data_43; // @[executor.scala 285:13]
    phv_data_44 <= io_pipe_phv_in_data_44; // @[executor.scala 285:13]
    phv_data_45 <= io_pipe_phv_in_data_45; // @[executor.scala 285:13]
    phv_data_46 <= io_pipe_phv_in_data_46; // @[executor.scala 285:13]
    phv_data_47 <= io_pipe_phv_in_data_47; // @[executor.scala 285:13]
    phv_data_48 <= io_pipe_phv_in_data_48; // @[executor.scala 285:13]
    phv_data_49 <= io_pipe_phv_in_data_49; // @[executor.scala 285:13]
    phv_data_50 <= io_pipe_phv_in_data_50; // @[executor.scala 285:13]
    phv_data_51 <= io_pipe_phv_in_data_51; // @[executor.scala 285:13]
    phv_data_52 <= io_pipe_phv_in_data_52; // @[executor.scala 285:13]
    phv_data_53 <= io_pipe_phv_in_data_53; // @[executor.scala 285:13]
    phv_data_54 <= io_pipe_phv_in_data_54; // @[executor.scala 285:13]
    phv_data_55 <= io_pipe_phv_in_data_55; // @[executor.scala 285:13]
    phv_data_56 <= io_pipe_phv_in_data_56; // @[executor.scala 285:13]
    phv_data_57 <= io_pipe_phv_in_data_57; // @[executor.scala 285:13]
    phv_data_58 <= io_pipe_phv_in_data_58; // @[executor.scala 285:13]
    phv_data_59 <= io_pipe_phv_in_data_59; // @[executor.scala 285:13]
    phv_data_60 <= io_pipe_phv_in_data_60; // @[executor.scala 285:13]
    phv_data_61 <= io_pipe_phv_in_data_61; // @[executor.scala 285:13]
    phv_data_62 <= io_pipe_phv_in_data_62; // @[executor.scala 285:13]
    phv_data_63 <= io_pipe_phv_in_data_63; // @[executor.scala 285:13]
    phv_data_64 <= io_pipe_phv_in_data_64; // @[executor.scala 285:13]
    phv_data_65 <= io_pipe_phv_in_data_65; // @[executor.scala 285:13]
    phv_data_66 <= io_pipe_phv_in_data_66; // @[executor.scala 285:13]
    phv_data_67 <= io_pipe_phv_in_data_67; // @[executor.scala 285:13]
    phv_data_68 <= io_pipe_phv_in_data_68; // @[executor.scala 285:13]
    phv_data_69 <= io_pipe_phv_in_data_69; // @[executor.scala 285:13]
    phv_data_70 <= io_pipe_phv_in_data_70; // @[executor.scala 285:13]
    phv_data_71 <= io_pipe_phv_in_data_71; // @[executor.scala 285:13]
    phv_data_72 <= io_pipe_phv_in_data_72; // @[executor.scala 285:13]
    phv_data_73 <= io_pipe_phv_in_data_73; // @[executor.scala 285:13]
    phv_data_74 <= io_pipe_phv_in_data_74; // @[executor.scala 285:13]
    phv_data_75 <= io_pipe_phv_in_data_75; // @[executor.scala 285:13]
    phv_data_76 <= io_pipe_phv_in_data_76; // @[executor.scala 285:13]
    phv_data_77 <= io_pipe_phv_in_data_77; // @[executor.scala 285:13]
    phv_data_78 <= io_pipe_phv_in_data_78; // @[executor.scala 285:13]
    phv_data_79 <= io_pipe_phv_in_data_79; // @[executor.scala 285:13]
    phv_data_80 <= io_pipe_phv_in_data_80; // @[executor.scala 285:13]
    phv_data_81 <= io_pipe_phv_in_data_81; // @[executor.scala 285:13]
    phv_data_82 <= io_pipe_phv_in_data_82; // @[executor.scala 285:13]
    phv_data_83 <= io_pipe_phv_in_data_83; // @[executor.scala 285:13]
    phv_data_84 <= io_pipe_phv_in_data_84; // @[executor.scala 285:13]
    phv_data_85 <= io_pipe_phv_in_data_85; // @[executor.scala 285:13]
    phv_data_86 <= io_pipe_phv_in_data_86; // @[executor.scala 285:13]
    phv_data_87 <= io_pipe_phv_in_data_87; // @[executor.scala 285:13]
    phv_data_88 <= io_pipe_phv_in_data_88; // @[executor.scala 285:13]
    phv_data_89 <= io_pipe_phv_in_data_89; // @[executor.scala 285:13]
    phv_data_90 <= io_pipe_phv_in_data_90; // @[executor.scala 285:13]
    phv_data_91 <= io_pipe_phv_in_data_91; // @[executor.scala 285:13]
    phv_data_92 <= io_pipe_phv_in_data_92; // @[executor.scala 285:13]
    phv_data_93 <= io_pipe_phv_in_data_93; // @[executor.scala 285:13]
    phv_data_94 <= io_pipe_phv_in_data_94; // @[executor.scala 285:13]
    phv_data_95 <= io_pipe_phv_in_data_95; // @[executor.scala 285:13]
    phv_data_96 <= io_pipe_phv_in_data_96; // @[executor.scala 285:13]
    phv_data_97 <= io_pipe_phv_in_data_97; // @[executor.scala 285:13]
    phv_data_98 <= io_pipe_phv_in_data_98; // @[executor.scala 285:13]
    phv_data_99 <= io_pipe_phv_in_data_99; // @[executor.scala 285:13]
    phv_data_100 <= io_pipe_phv_in_data_100; // @[executor.scala 285:13]
    phv_data_101 <= io_pipe_phv_in_data_101; // @[executor.scala 285:13]
    phv_data_102 <= io_pipe_phv_in_data_102; // @[executor.scala 285:13]
    phv_data_103 <= io_pipe_phv_in_data_103; // @[executor.scala 285:13]
    phv_data_104 <= io_pipe_phv_in_data_104; // @[executor.scala 285:13]
    phv_data_105 <= io_pipe_phv_in_data_105; // @[executor.scala 285:13]
    phv_data_106 <= io_pipe_phv_in_data_106; // @[executor.scala 285:13]
    phv_data_107 <= io_pipe_phv_in_data_107; // @[executor.scala 285:13]
    phv_data_108 <= io_pipe_phv_in_data_108; // @[executor.scala 285:13]
    phv_data_109 <= io_pipe_phv_in_data_109; // @[executor.scala 285:13]
    phv_data_110 <= io_pipe_phv_in_data_110; // @[executor.scala 285:13]
    phv_data_111 <= io_pipe_phv_in_data_111; // @[executor.scala 285:13]
    phv_data_112 <= io_pipe_phv_in_data_112; // @[executor.scala 285:13]
    phv_data_113 <= io_pipe_phv_in_data_113; // @[executor.scala 285:13]
    phv_data_114 <= io_pipe_phv_in_data_114; // @[executor.scala 285:13]
    phv_data_115 <= io_pipe_phv_in_data_115; // @[executor.scala 285:13]
    phv_data_116 <= io_pipe_phv_in_data_116; // @[executor.scala 285:13]
    phv_data_117 <= io_pipe_phv_in_data_117; // @[executor.scala 285:13]
    phv_data_118 <= io_pipe_phv_in_data_118; // @[executor.scala 285:13]
    phv_data_119 <= io_pipe_phv_in_data_119; // @[executor.scala 285:13]
    phv_data_120 <= io_pipe_phv_in_data_120; // @[executor.scala 285:13]
    phv_data_121 <= io_pipe_phv_in_data_121; // @[executor.scala 285:13]
    phv_data_122 <= io_pipe_phv_in_data_122; // @[executor.scala 285:13]
    phv_data_123 <= io_pipe_phv_in_data_123; // @[executor.scala 285:13]
    phv_data_124 <= io_pipe_phv_in_data_124; // @[executor.scala 285:13]
    phv_data_125 <= io_pipe_phv_in_data_125; // @[executor.scala 285:13]
    phv_data_126 <= io_pipe_phv_in_data_126; // @[executor.scala 285:13]
    phv_data_127 <= io_pipe_phv_in_data_127; // @[executor.scala 285:13]
    phv_data_128 <= io_pipe_phv_in_data_128; // @[executor.scala 285:13]
    phv_data_129 <= io_pipe_phv_in_data_129; // @[executor.scala 285:13]
    phv_data_130 <= io_pipe_phv_in_data_130; // @[executor.scala 285:13]
    phv_data_131 <= io_pipe_phv_in_data_131; // @[executor.scala 285:13]
    phv_data_132 <= io_pipe_phv_in_data_132; // @[executor.scala 285:13]
    phv_data_133 <= io_pipe_phv_in_data_133; // @[executor.scala 285:13]
    phv_data_134 <= io_pipe_phv_in_data_134; // @[executor.scala 285:13]
    phv_data_135 <= io_pipe_phv_in_data_135; // @[executor.scala 285:13]
    phv_data_136 <= io_pipe_phv_in_data_136; // @[executor.scala 285:13]
    phv_data_137 <= io_pipe_phv_in_data_137; // @[executor.scala 285:13]
    phv_data_138 <= io_pipe_phv_in_data_138; // @[executor.scala 285:13]
    phv_data_139 <= io_pipe_phv_in_data_139; // @[executor.scala 285:13]
    phv_data_140 <= io_pipe_phv_in_data_140; // @[executor.scala 285:13]
    phv_data_141 <= io_pipe_phv_in_data_141; // @[executor.scala 285:13]
    phv_data_142 <= io_pipe_phv_in_data_142; // @[executor.scala 285:13]
    phv_data_143 <= io_pipe_phv_in_data_143; // @[executor.scala 285:13]
    phv_data_144 <= io_pipe_phv_in_data_144; // @[executor.scala 285:13]
    phv_data_145 <= io_pipe_phv_in_data_145; // @[executor.scala 285:13]
    phv_data_146 <= io_pipe_phv_in_data_146; // @[executor.scala 285:13]
    phv_data_147 <= io_pipe_phv_in_data_147; // @[executor.scala 285:13]
    phv_data_148 <= io_pipe_phv_in_data_148; // @[executor.scala 285:13]
    phv_data_149 <= io_pipe_phv_in_data_149; // @[executor.scala 285:13]
    phv_data_150 <= io_pipe_phv_in_data_150; // @[executor.scala 285:13]
    phv_data_151 <= io_pipe_phv_in_data_151; // @[executor.scala 285:13]
    phv_data_152 <= io_pipe_phv_in_data_152; // @[executor.scala 285:13]
    phv_data_153 <= io_pipe_phv_in_data_153; // @[executor.scala 285:13]
    phv_data_154 <= io_pipe_phv_in_data_154; // @[executor.scala 285:13]
    phv_data_155 <= io_pipe_phv_in_data_155; // @[executor.scala 285:13]
    phv_data_156 <= io_pipe_phv_in_data_156; // @[executor.scala 285:13]
    phv_data_157 <= io_pipe_phv_in_data_157; // @[executor.scala 285:13]
    phv_data_158 <= io_pipe_phv_in_data_158; // @[executor.scala 285:13]
    phv_data_159 <= io_pipe_phv_in_data_159; // @[executor.scala 285:13]
    phv_header_0 <= io_pipe_phv_in_header_0; // @[executor.scala 285:13]
    phv_header_1 <= io_pipe_phv_in_header_1; // @[executor.scala 285:13]
    phv_header_2 <= io_pipe_phv_in_header_2; // @[executor.scala 285:13]
    phv_header_3 <= io_pipe_phv_in_header_3; // @[executor.scala 285:13]
    phv_header_4 <= io_pipe_phv_in_header_4; // @[executor.scala 285:13]
    phv_header_5 <= io_pipe_phv_in_header_5; // @[executor.scala 285:13]
    phv_header_6 <= io_pipe_phv_in_header_6; // @[executor.scala 285:13]
    phv_header_7 <= io_pipe_phv_in_header_7; // @[executor.scala 285:13]
    phv_header_8 <= io_pipe_phv_in_header_8; // @[executor.scala 285:13]
    phv_header_9 <= io_pipe_phv_in_header_9; // @[executor.scala 285:13]
    phv_header_10 <= io_pipe_phv_in_header_10; // @[executor.scala 285:13]
    phv_header_11 <= io_pipe_phv_in_header_11; // @[executor.scala 285:13]
    phv_header_12 <= io_pipe_phv_in_header_12; // @[executor.scala 285:13]
    phv_header_13 <= io_pipe_phv_in_header_13; // @[executor.scala 285:13]
    phv_header_14 <= io_pipe_phv_in_header_14; // @[executor.scala 285:13]
    phv_header_15 <= io_pipe_phv_in_header_15; // @[executor.scala 285:13]
    phv_parse_current_state <= io_pipe_phv_in_parse_current_state; // @[executor.scala 285:13]
    phv_parse_current_offset <= io_pipe_phv_in_parse_current_offset; // @[executor.scala 285:13]
    phv_parse_transition_field <= io_pipe_phv_in_parse_transition_field; // @[executor.scala 285:13]
    phv_next_processor_id <= io_pipe_phv_in_next_processor_id; // @[executor.scala 285:13]
    phv_next_config_id <= io_pipe_phv_in_next_config_id; // @[executor.scala 285:13]
    phv_is_valid_processor <= io_pipe_phv_in_is_valid_processor; // @[executor.scala 285:13]
    offset_0 <= io_offset_in_0; // @[executor.scala 291:16]
    offset_1 <= io_offset_in_1; // @[executor.scala 291:16]
    offset_2 <= io_offset_in_2; // @[executor.scala 291:16]
    offset_3 <= io_offset_in_3; // @[executor.scala 291:16]
    length_0 <= io_length_in_0; // @[executor.scala 292:16]
    length_1 <= io_length_in_1; // @[executor.scala 292:16]
    length_2 <= io_length_in_2; // @[executor.scala 292:16]
    length_3 <= io_length_in_3; // @[executor.scala 292:16]
    field_0 <= io_field_in_0; // @[executor.scala 293:16]
    field_1 <= io_field_in_1; // @[executor.scala 293:16]
    field_2 <= io_field_in_2; // @[executor.scala 293:16]
    field_3 <= io_field_in_3; // @[executor.scala 293:16]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  phv_data_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  phv_data_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  phv_data_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  phv_data_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  phv_data_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  phv_data_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  phv_data_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  phv_data_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  phv_data_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  phv_data_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  phv_data_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  phv_data_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  phv_data_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  phv_data_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  phv_data_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  phv_data_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  phv_data_16 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  phv_data_17 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  phv_data_18 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  phv_data_19 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  phv_data_20 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  phv_data_21 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  phv_data_22 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  phv_data_23 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  phv_data_24 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  phv_data_25 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  phv_data_26 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  phv_data_27 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  phv_data_28 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  phv_data_29 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  phv_data_30 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  phv_data_31 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  phv_data_32 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  phv_data_33 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  phv_data_34 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  phv_data_35 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  phv_data_36 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  phv_data_37 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  phv_data_38 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  phv_data_39 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  phv_data_40 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  phv_data_41 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  phv_data_42 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  phv_data_43 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  phv_data_44 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  phv_data_45 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  phv_data_46 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  phv_data_47 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  phv_data_48 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  phv_data_49 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  phv_data_50 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  phv_data_51 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  phv_data_52 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  phv_data_53 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  phv_data_54 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  phv_data_55 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  phv_data_56 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  phv_data_57 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  phv_data_58 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  phv_data_59 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  phv_data_60 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  phv_data_61 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  phv_data_62 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  phv_data_63 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  phv_data_64 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  phv_data_65 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  phv_data_66 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  phv_data_67 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  phv_data_68 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  phv_data_69 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  phv_data_70 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  phv_data_71 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  phv_data_72 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  phv_data_73 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  phv_data_74 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  phv_data_75 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  phv_data_76 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  phv_data_77 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  phv_data_78 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  phv_data_79 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  phv_data_80 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  phv_data_81 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  phv_data_82 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  phv_data_83 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  phv_data_84 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  phv_data_85 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  phv_data_86 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  phv_data_87 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  phv_data_88 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  phv_data_89 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  phv_data_90 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  phv_data_91 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  phv_data_92 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  phv_data_93 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  phv_data_94 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  phv_data_95 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  phv_data_96 = _RAND_96[7:0];
  _RAND_97 = {1{`RANDOM}};
  phv_data_97 = _RAND_97[7:0];
  _RAND_98 = {1{`RANDOM}};
  phv_data_98 = _RAND_98[7:0];
  _RAND_99 = {1{`RANDOM}};
  phv_data_99 = _RAND_99[7:0];
  _RAND_100 = {1{`RANDOM}};
  phv_data_100 = _RAND_100[7:0];
  _RAND_101 = {1{`RANDOM}};
  phv_data_101 = _RAND_101[7:0];
  _RAND_102 = {1{`RANDOM}};
  phv_data_102 = _RAND_102[7:0];
  _RAND_103 = {1{`RANDOM}};
  phv_data_103 = _RAND_103[7:0];
  _RAND_104 = {1{`RANDOM}};
  phv_data_104 = _RAND_104[7:0];
  _RAND_105 = {1{`RANDOM}};
  phv_data_105 = _RAND_105[7:0];
  _RAND_106 = {1{`RANDOM}};
  phv_data_106 = _RAND_106[7:0];
  _RAND_107 = {1{`RANDOM}};
  phv_data_107 = _RAND_107[7:0];
  _RAND_108 = {1{`RANDOM}};
  phv_data_108 = _RAND_108[7:0];
  _RAND_109 = {1{`RANDOM}};
  phv_data_109 = _RAND_109[7:0];
  _RAND_110 = {1{`RANDOM}};
  phv_data_110 = _RAND_110[7:0];
  _RAND_111 = {1{`RANDOM}};
  phv_data_111 = _RAND_111[7:0];
  _RAND_112 = {1{`RANDOM}};
  phv_data_112 = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  phv_data_113 = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  phv_data_114 = _RAND_114[7:0];
  _RAND_115 = {1{`RANDOM}};
  phv_data_115 = _RAND_115[7:0];
  _RAND_116 = {1{`RANDOM}};
  phv_data_116 = _RAND_116[7:0];
  _RAND_117 = {1{`RANDOM}};
  phv_data_117 = _RAND_117[7:0];
  _RAND_118 = {1{`RANDOM}};
  phv_data_118 = _RAND_118[7:0];
  _RAND_119 = {1{`RANDOM}};
  phv_data_119 = _RAND_119[7:0];
  _RAND_120 = {1{`RANDOM}};
  phv_data_120 = _RAND_120[7:0];
  _RAND_121 = {1{`RANDOM}};
  phv_data_121 = _RAND_121[7:0];
  _RAND_122 = {1{`RANDOM}};
  phv_data_122 = _RAND_122[7:0];
  _RAND_123 = {1{`RANDOM}};
  phv_data_123 = _RAND_123[7:0];
  _RAND_124 = {1{`RANDOM}};
  phv_data_124 = _RAND_124[7:0];
  _RAND_125 = {1{`RANDOM}};
  phv_data_125 = _RAND_125[7:0];
  _RAND_126 = {1{`RANDOM}};
  phv_data_126 = _RAND_126[7:0];
  _RAND_127 = {1{`RANDOM}};
  phv_data_127 = _RAND_127[7:0];
  _RAND_128 = {1{`RANDOM}};
  phv_data_128 = _RAND_128[7:0];
  _RAND_129 = {1{`RANDOM}};
  phv_data_129 = _RAND_129[7:0];
  _RAND_130 = {1{`RANDOM}};
  phv_data_130 = _RAND_130[7:0];
  _RAND_131 = {1{`RANDOM}};
  phv_data_131 = _RAND_131[7:0];
  _RAND_132 = {1{`RANDOM}};
  phv_data_132 = _RAND_132[7:0];
  _RAND_133 = {1{`RANDOM}};
  phv_data_133 = _RAND_133[7:0];
  _RAND_134 = {1{`RANDOM}};
  phv_data_134 = _RAND_134[7:0];
  _RAND_135 = {1{`RANDOM}};
  phv_data_135 = _RAND_135[7:0];
  _RAND_136 = {1{`RANDOM}};
  phv_data_136 = _RAND_136[7:0];
  _RAND_137 = {1{`RANDOM}};
  phv_data_137 = _RAND_137[7:0];
  _RAND_138 = {1{`RANDOM}};
  phv_data_138 = _RAND_138[7:0];
  _RAND_139 = {1{`RANDOM}};
  phv_data_139 = _RAND_139[7:0];
  _RAND_140 = {1{`RANDOM}};
  phv_data_140 = _RAND_140[7:0];
  _RAND_141 = {1{`RANDOM}};
  phv_data_141 = _RAND_141[7:0];
  _RAND_142 = {1{`RANDOM}};
  phv_data_142 = _RAND_142[7:0];
  _RAND_143 = {1{`RANDOM}};
  phv_data_143 = _RAND_143[7:0];
  _RAND_144 = {1{`RANDOM}};
  phv_data_144 = _RAND_144[7:0];
  _RAND_145 = {1{`RANDOM}};
  phv_data_145 = _RAND_145[7:0];
  _RAND_146 = {1{`RANDOM}};
  phv_data_146 = _RAND_146[7:0];
  _RAND_147 = {1{`RANDOM}};
  phv_data_147 = _RAND_147[7:0];
  _RAND_148 = {1{`RANDOM}};
  phv_data_148 = _RAND_148[7:0];
  _RAND_149 = {1{`RANDOM}};
  phv_data_149 = _RAND_149[7:0];
  _RAND_150 = {1{`RANDOM}};
  phv_data_150 = _RAND_150[7:0];
  _RAND_151 = {1{`RANDOM}};
  phv_data_151 = _RAND_151[7:0];
  _RAND_152 = {1{`RANDOM}};
  phv_data_152 = _RAND_152[7:0];
  _RAND_153 = {1{`RANDOM}};
  phv_data_153 = _RAND_153[7:0];
  _RAND_154 = {1{`RANDOM}};
  phv_data_154 = _RAND_154[7:0];
  _RAND_155 = {1{`RANDOM}};
  phv_data_155 = _RAND_155[7:0];
  _RAND_156 = {1{`RANDOM}};
  phv_data_156 = _RAND_156[7:0];
  _RAND_157 = {1{`RANDOM}};
  phv_data_157 = _RAND_157[7:0];
  _RAND_158 = {1{`RANDOM}};
  phv_data_158 = _RAND_158[7:0];
  _RAND_159 = {1{`RANDOM}};
  phv_data_159 = _RAND_159[7:0];
  _RAND_160 = {1{`RANDOM}};
  phv_header_0 = _RAND_160[15:0];
  _RAND_161 = {1{`RANDOM}};
  phv_header_1 = _RAND_161[15:0];
  _RAND_162 = {1{`RANDOM}};
  phv_header_2 = _RAND_162[15:0];
  _RAND_163 = {1{`RANDOM}};
  phv_header_3 = _RAND_163[15:0];
  _RAND_164 = {1{`RANDOM}};
  phv_header_4 = _RAND_164[15:0];
  _RAND_165 = {1{`RANDOM}};
  phv_header_5 = _RAND_165[15:0];
  _RAND_166 = {1{`RANDOM}};
  phv_header_6 = _RAND_166[15:0];
  _RAND_167 = {1{`RANDOM}};
  phv_header_7 = _RAND_167[15:0];
  _RAND_168 = {1{`RANDOM}};
  phv_header_8 = _RAND_168[15:0];
  _RAND_169 = {1{`RANDOM}};
  phv_header_9 = _RAND_169[15:0];
  _RAND_170 = {1{`RANDOM}};
  phv_header_10 = _RAND_170[15:0];
  _RAND_171 = {1{`RANDOM}};
  phv_header_11 = _RAND_171[15:0];
  _RAND_172 = {1{`RANDOM}};
  phv_header_12 = _RAND_172[15:0];
  _RAND_173 = {1{`RANDOM}};
  phv_header_13 = _RAND_173[15:0];
  _RAND_174 = {1{`RANDOM}};
  phv_header_14 = _RAND_174[15:0];
  _RAND_175 = {1{`RANDOM}};
  phv_header_15 = _RAND_175[15:0];
  _RAND_176 = {1{`RANDOM}};
  phv_parse_current_state = _RAND_176[7:0];
  _RAND_177 = {1{`RANDOM}};
  phv_parse_current_offset = _RAND_177[7:0];
  _RAND_178 = {1{`RANDOM}};
  phv_parse_transition_field = _RAND_178[15:0];
  _RAND_179 = {1{`RANDOM}};
  phv_next_processor_id = _RAND_179[3:0];
  _RAND_180 = {1{`RANDOM}};
  phv_next_config_id = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  phv_is_valid_processor = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  offset_0 = _RAND_182[7:0];
  _RAND_183 = {1{`RANDOM}};
  offset_1 = _RAND_183[7:0];
  _RAND_184 = {1{`RANDOM}};
  offset_2 = _RAND_184[7:0];
  _RAND_185 = {1{`RANDOM}};
  offset_3 = _RAND_185[7:0];
  _RAND_186 = {1{`RANDOM}};
  length_0 = _RAND_186[7:0];
  _RAND_187 = {1{`RANDOM}};
  length_1 = _RAND_187[7:0];
  _RAND_188 = {1{`RANDOM}};
  length_2 = _RAND_188[7:0];
  _RAND_189 = {1{`RANDOM}};
  length_3 = _RAND_189[7:0];
  _RAND_190 = {2{`RANDOM}};
  field_0 = _RAND_190[63:0];
  _RAND_191 = {2{`RANDOM}};
  field_1 = _RAND_191[63:0];
  _RAND_192 = {2{`RANDOM}};
  field_2 = _RAND_192[63:0];
  _RAND_193 = {2{`RANDOM}};
  field_3 = _RAND_193[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
