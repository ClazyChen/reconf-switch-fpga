module MatchGetKeyPISA(
  input          clock,
  input  [7:0]   io_pipe_phv_in_data_0,
  input  [7:0]   io_pipe_phv_in_data_1,
  input  [7:0]   io_pipe_phv_in_data_2,
  input  [7:0]   io_pipe_phv_in_data_3,
  input  [7:0]   io_pipe_phv_in_data_4,
  input  [7:0]   io_pipe_phv_in_data_5,
  input  [7:0]   io_pipe_phv_in_data_6,
  input  [7:0]   io_pipe_phv_in_data_7,
  input  [7:0]   io_pipe_phv_in_data_8,
  input  [7:0]   io_pipe_phv_in_data_9,
  input  [7:0]   io_pipe_phv_in_data_10,
  input  [7:0]   io_pipe_phv_in_data_11,
  input  [7:0]   io_pipe_phv_in_data_12,
  input  [7:0]   io_pipe_phv_in_data_13,
  input  [7:0]   io_pipe_phv_in_data_14,
  input  [7:0]   io_pipe_phv_in_data_15,
  input  [7:0]   io_pipe_phv_in_data_16,
  input  [7:0]   io_pipe_phv_in_data_17,
  input  [7:0]   io_pipe_phv_in_data_18,
  input  [7:0]   io_pipe_phv_in_data_19,
  input  [7:0]   io_pipe_phv_in_data_20,
  input  [7:0]   io_pipe_phv_in_data_21,
  input  [7:0]   io_pipe_phv_in_data_22,
  input  [7:0]   io_pipe_phv_in_data_23,
  input  [7:0]   io_pipe_phv_in_data_24,
  input  [7:0]   io_pipe_phv_in_data_25,
  input  [7:0]   io_pipe_phv_in_data_26,
  input  [7:0]   io_pipe_phv_in_data_27,
  input  [7:0]   io_pipe_phv_in_data_28,
  input  [7:0]   io_pipe_phv_in_data_29,
  input  [7:0]   io_pipe_phv_in_data_30,
  input  [7:0]   io_pipe_phv_in_data_31,
  input  [7:0]   io_pipe_phv_in_data_32,
  input  [7:0]   io_pipe_phv_in_data_33,
  input  [7:0]   io_pipe_phv_in_data_34,
  input  [7:0]   io_pipe_phv_in_data_35,
  input  [7:0]   io_pipe_phv_in_data_36,
  input  [7:0]   io_pipe_phv_in_data_37,
  input  [7:0]   io_pipe_phv_in_data_38,
  input  [7:0]   io_pipe_phv_in_data_39,
  input  [7:0]   io_pipe_phv_in_data_40,
  input  [7:0]   io_pipe_phv_in_data_41,
  input  [7:0]   io_pipe_phv_in_data_42,
  input  [7:0]   io_pipe_phv_in_data_43,
  input  [7:0]   io_pipe_phv_in_data_44,
  input  [7:0]   io_pipe_phv_in_data_45,
  input  [7:0]   io_pipe_phv_in_data_46,
  input  [7:0]   io_pipe_phv_in_data_47,
  input  [7:0]   io_pipe_phv_in_data_48,
  input  [7:0]   io_pipe_phv_in_data_49,
  input  [7:0]   io_pipe_phv_in_data_50,
  input  [7:0]   io_pipe_phv_in_data_51,
  input  [7:0]   io_pipe_phv_in_data_52,
  input  [7:0]   io_pipe_phv_in_data_53,
  input  [7:0]   io_pipe_phv_in_data_54,
  input  [7:0]   io_pipe_phv_in_data_55,
  input  [7:0]   io_pipe_phv_in_data_56,
  input  [7:0]   io_pipe_phv_in_data_57,
  input  [7:0]   io_pipe_phv_in_data_58,
  input  [7:0]   io_pipe_phv_in_data_59,
  input  [7:0]   io_pipe_phv_in_data_60,
  input  [7:0]   io_pipe_phv_in_data_61,
  input  [7:0]   io_pipe_phv_in_data_62,
  input  [7:0]   io_pipe_phv_in_data_63,
  input  [7:0]   io_pipe_phv_in_data_64,
  input  [7:0]   io_pipe_phv_in_data_65,
  input  [7:0]   io_pipe_phv_in_data_66,
  input  [7:0]   io_pipe_phv_in_data_67,
  input  [7:0]   io_pipe_phv_in_data_68,
  input  [7:0]   io_pipe_phv_in_data_69,
  input  [7:0]   io_pipe_phv_in_data_70,
  input  [7:0]   io_pipe_phv_in_data_71,
  input  [7:0]   io_pipe_phv_in_data_72,
  input  [7:0]   io_pipe_phv_in_data_73,
  input  [7:0]   io_pipe_phv_in_data_74,
  input  [7:0]   io_pipe_phv_in_data_75,
  input  [7:0]   io_pipe_phv_in_data_76,
  input  [7:0]   io_pipe_phv_in_data_77,
  input  [7:0]   io_pipe_phv_in_data_78,
  input  [7:0]   io_pipe_phv_in_data_79,
  input  [7:0]   io_pipe_phv_in_data_80,
  input  [7:0]   io_pipe_phv_in_data_81,
  input  [7:0]   io_pipe_phv_in_data_82,
  input  [7:0]   io_pipe_phv_in_data_83,
  input  [7:0]   io_pipe_phv_in_data_84,
  input  [7:0]   io_pipe_phv_in_data_85,
  input  [7:0]   io_pipe_phv_in_data_86,
  input  [7:0]   io_pipe_phv_in_data_87,
  input  [7:0]   io_pipe_phv_in_data_88,
  input  [7:0]   io_pipe_phv_in_data_89,
  input  [7:0]   io_pipe_phv_in_data_90,
  input  [7:0]   io_pipe_phv_in_data_91,
  input  [7:0]   io_pipe_phv_in_data_92,
  input  [7:0]   io_pipe_phv_in_data_93,
  input  [7:0]   io_pipe_phv_in_data_94,
  input  [7:0]   io_pipe_phv_in_data_95,
  input  [7:0]   io_pipe_phv_in_data_96,
  input  [7:0]   io_pipe_phv_in_data_97,
  input  [7:0]   io_pipe_phv_in_data_98,
  input  [7:0]   io_pipe_phv_in_data_99,
  input  [7:0]   io_pipe_phv_in_data_100,
  input  [7:0]   io_pipe_phv_in_data_101,
  input  [7:0]   io_pipe_phv_in_data_102,
  input  [7:0]   io_pipe_phv_in_data_103,
  input  [7:0]   io_pipe_phv_in_data_104,
  input  [7:0]   io_pipe_phv_in_data_105,
  input  [7:0]   io_pipe_phv_in_data_106,
  input  [7:0]   io_pipe_phv_in_data_107,
  input  [7:0]   io_pipe_phv_in_data_108,
  input  [7:0]   io_pipe_phv_in_data_109,
  input  [7:0]   io_pipe_phv_in_data_110,
  input  [7:0]   io_pipe_phv_in_data_111,
  input  [7:0]   io_pipe_phv_in_data_112,
  input  [7:0]   io_pipe_phv_in_data_113,
  input  [7:0]   io_pipe_phv_in_data_114,
  input  [7:0]   io_pipe_phv_in_data_115,
  input  [7:0]   io_pipe_phv_in_data_116,
  input  [7:0]   io_pipe_phv_in_data_117,
  input  [7:0]   io_pipe_phv_in_data_118,
  input  [7:0]   io_pipe_phv_in_data_119,
  input  [7:0]   io_pipe_phv_in_data_120,
  input  [7:0]   io_pipe_phv_in_data_121,
  input  [7:0]   io_pipe_phv_in_data_122,
  input  [7:0]   io_pipe_phv_in_data_123,
  input  [7:0]   io_pipe_phv_in_data_124,
  input  [7:0]   io_pipe_phv_in_data_125,
  input  [7:0]   io_pipe_phv_in_data_126,
  input  [7:0]   io_pipe_phv_in_data_127,
  input  [7:0]   io_pipe_phv_in_data_128,
  input  [7:0]   io_pipe_phv_in_data_129,
  input  [7:0]   io_pipe_phv_in_data_130,
  input  [7:0]   io_pipe_phv_in_data_131,
  input  [7:0]   io_pipe_phv_in_data_132,
  input  [7:0]   io_pipe_phv_in_data_133,
  input  [7:0]   io_pipe_phv_in_data_134,
  input  [7:0]   io_pipe_phv_in_data_135,
  input  [7:0]   io_pipe_phv_in_data_136,
  input  [7:0]   io_pipe_phv_in_data_137,
  input  [7:0]   io_pipe_phv_in_data_138,
  input  [7:0]   io_pipe_phv_in_data_139,
  input  [7:0]   io_pipe_phv_in_data_140,
  input  [7:0]   io_pipe_phv_in_data_141,
  input  [7:0]   io_pipe_phv_in_data_142,
  input  [7:0]   io_pipe_phv_in_data_143,
  input  [7:0]   io_pipe_phv_in_data_144,
  input  [7:0]   io_pipe_phv_in_data_145,
  input  [7:0]   io_pipe_phv_in_data_146,
  input  [7:0]   io_pipe_phv_in_data_147,
  input  [7:0]   io_pipe_phv_in_data_148,
  input  [7:0]   io_pipe_phv_in_data_149,
  input  [7:0]   io_pipe_phv_in_data_150,
  input  [7:0]   io_pipe_phv_in_data_151,
  input  [7:0]   io_pipe_phv_in_data_152,
  input  [7:0]   io_pipe_phv_in_data_153,
  input  [7:0]   io_pipe_phv_in_data_154,
  input  [7:0]   io_pipe_phv_in_data_155,
  input  [7:0]   io_pipe_phv_in_data_156,
  input  [7:0]   io_pipe_phv_in_data_157,
  input  [7:0]   io_pipe_phv_in_data_158,
  input  [7:0]   io_pipe_phv_in_data_159,
  input  [7:0]   io_pipe_phv_in_data_160,
  input  [7:0]   io_pipe_phv_in_data_161,
  input  [7:0]   io_pipe_phv_in_data_162,
  input  [7:0]   io_pipe_phv_in_data_163,
  input  [7:0]   io_pipe_phv_in_data_164,
  input  [7:0]   io_pipe_phv_in_data_165,
  input  [7:0]   io_pipe_phv_in_data_166,
  input  [7:0]   io_pipe_phv_in_data_167,
  input  [7:0]   io_pipe_phv_in_data_168,
  input  [7:0]   io_pipe_phv_in_data_169,
  input  [7:0]   io_pipe_phv_in_data_170,
  input  [7:0]   io_pipe_phv_in_data_171,
  input  [7:0]   io_pipe_phv_in_data_172,
  input  [7:0]   io_pipe_phv_in_data_173,
  input  [7:0]   io_pipe_phv_in_data_174,
  input  [7:0]   io_pipe_phv_in_data_175,
  input  [7:0]   io_pipe_phv_in_data_176,
  input  [7:0]   io_pipe_phv_in_data_177,
  input  [7:0]   io_pipe_phv_in_data_178,
  input  [7:0]   io_pipe_phv_in_data_179,
  input  [7:0]   io_pipe_phv_in_data_180,
  input  [7:0]   io_pipe_phv_in_data_181,
  input  [7:0]   io_pipe_phv_in_data_182,
  input  [7:0]   io_pipe_phv_in_data_183,
  input  [7:0]   io_pipe_phv_in_data_184,
  input  [7:0]   io_pipe_phv_in_data_185,
  input  [7:0]   io_pipe_phv_in_data_186,
  input  [7:0]   io_pipe_phv_in_data_187,
  input  [7:0]   io_pipe_phv_in_data_188,
  input  [7:0]   io_pipe_phv_in_data_189,
  input  [7:0]   io_pipe_phv_in_data_190,
  input  [7:0]   io_pipe_phv_in_data_191,
  input  [7:0]   io_pipe_phv_in_data_192,
  input  [7:0]   io_pipe_phv_in_data_193,
  input  [7:0]   io_pipe_phv_in_data_194,
  input  [7:0]   io_pipe_phv_in_data_195,
  input  [7:0]   io_pipe_phv_in_data_196,
  input  [7:0]   io_pipe_phv_in_data_197,
  input  [7:0]   io_pipe_phv_in_data_198,
  input  [7:0]   io_pipe_phv_in_data_199,
  input  [7:0]   io_pipe_phv_in_data_200,
  input  [7:0]   io_pipe_phv_in_data_201,
  input  [7:0]   io_pipe_phv_in_data_202,
  input  [7:0]   io_pipe_phv_in_data_203,
  input  [7:0]   io_pipe_phv_in_data_204,
  input  [7:0]   io_pipe_phv_in_data_205,
  input  [7:0]   io_pipe_phv_in_data_206,
  input  [7:0]   io_pipe_phv_in_data_207,
  input  [7:0]   io_pipe_phv_in_data_208,
  input  [7:0]   io_pipe_phv_in_data_209,
  input  [7:0]   io_pipe_phv_in_data_210,
  input  [7:0]   io_pipe_phv_in_data_211,
  input  [7:0]   io_pipe_phv_in_data_212,
  input  [7:0]   io_pipe_phv_in_data_213,
  input  [7:0]   io_pipe_phv_in_data_214,
  input  [7:0]   io_pipe_phv_in_data_215,
  input  [7:0]   io_pipe_phv_in_data_216,
  input  [7:0]   io_pipe_phv_in_data_217,
  input  [7:0]   io_pipe_phv_in_data_218,
  input  [7:0]   io_pipe_phv_in_data_219,
  input  [7:0]   io_pipe_phv_in_data_220,
  input  [7:0]   io_pipe_phv_in_data_221,
  input  [7:0]   io_pipe_phv_in_data_222,
  input  [7:0]   io_pipe_phv_in_data_223,
  input  [7:0]   io_pipe_phv_in_data_224,
  input  [7:0]   io_pipe_phv_in_data_225,
  input  [7:0]   io_pipe_phv_in_data_226,
  input  [7:0]   io_pipe_phv_in_data_227,
  input  [7:0]   io_pipe_phv_in_data_228,
  input  [7:0]   io_pipe_phv_in_data_229,
  input  [7:0]   io_pipe_phv_in_data_230,
  input  [7:0]   io_pipe_phv_in_data_231,
  input  [7:0]   io_pipe_phv_in_data_232,
  input  [7:0]   io_pipe_phv_in_data_233,
  input  [7:0]   io_pipe_phv_in_data_234,
  input  [7:0]   io_pipe_phv_in_data_235,
  input  [7:0]   io_pipe_phv_in_data_236,
  input  [7:0]   io_pipe_phv_in_data_237,
  input  [7:0]   io_pipe_phv_in_data_238,
  input  [7:0]   io_pipe_phv_in_data_239,
  input  [7:0]   io_pipe_phv_in_data_240,
  input  [7:0]   io_pipe_phv_in_data_241,
  input  [7:0]   io_pipe_phv_in_data_242,
  input  [7:0]   io_pipe_phv_in_data_243,
  input  [7:0]   io_pipe_phv_in_data_244,
  input  [7:0]   io_pipe_phv_in_data_245,
  input  [7:0]   io_pipe_phv_in_data_246,
  input  [7:0]   io_pipe_phv_in_data_247,
  input  [7:0]   io_pipe_phv_in_data_248,
  input  [7:0]   io_pipe_phv_in_data_249,
  input  [7:0]   io_pipe_phv_in_data_250,
  input  [7:0]   io_pipe_phv_in_data_251,
  input  [7:0]   io_pipe_phv_in_data_252,
  input  [7:0]   io_pipe_phv_in_data_253,
  input  [7:0]   io_pipe_phv_in_data_254,
  input  [7:0]   io_pipe_phv_in_data_255,
  input  [7:0]   io_pipe_phv_in_data_256,
  input  [7:0]   io_pipe_phv_in_data_257,
  input  [7:0]   io_pipe_phv_in_data_258,
  input  [7:0]   io_pipe_phv_in_data_259,
  input  [7:0]   io_pipe_phv_in_data_260,
  input  [7:0]   io_pipe_phv_in_data_261,
  input  [7:0]   io_pipe_phv_in_data_262,
  input  [7:0]   io_pipe_phv_in_data_263,
  input  [7:0]   io_pipe_phv_in_data_264,
  input  [7:0]   io_pipe_phv_in_data_265,
  input  [7:0]   io_pipe_phv_in_data_266,
  input  [7:0]   io_pipe_phv_in_data_267,
  input  [7:0]   io_pipe_phv_in_data_268,
  input  [7:0]   io_pipe_phv_in_data_269,
  input  [7:0]   io_pipe_phv_in_data_270,
  input  [7:0]   io_pipe_phv_in_data_271,
  input  [7:0]   io_pipe_phv_in_data_272,
  input  [7:0]   io_pipe_phv_in_data_273,
  input  [7:0]   io_pipe_phv_in_data_274,
  input  [7:0]   io_pipe_phv_in_data_275,
  input  [7:0]   io_pipe_phv_in_data_276,
  input  [7:0]   io_pipe_phv_in_data_277,
  input  [7:0]   io_pipe_phv_in_data_278,
  input  [7:0]   io_pipe_phv_in_data_279,
  input  [7:0]   io_pipe_phv_in_data_280,
  input  [7:0]   io_pipe_phv_in_data_281,
  input  [7:0]   io_pipe_phv_in_data_282,
  input  [7:0]   io_pipe_phv_in_data_283,
  input  [7:0]   io_pipe_phv_in_data_284,
  input  [7:0]   io_pipe_phv_in_data_285,
  input  [7:0]   io_pipe_phv_in_data_286,
  input  [7:0]   io_pipe_phv_in_data_287,
  input  [7:0]   io_pipe_phv_in_data_288,
  input  [7:0]   io_pipe_phv_in_data_289,
  input  [7:0]   io_pipe_phv_in_data_290,
  input  [7:0]   io_pipe_phv_in_data_291,
  input  [7:0]   io_pipe_phv_in_data_292,
  input  [7:0]   io_pipe_phv_in_data_293,
  input  [7:0]   io_pipe_phv_in_data_294,
  input  [7:0]   io_pipe_phv_in_data_295,
  input  [7:0]   io_pipe_phv_in_data_296,
  input  [7:0]   io_pipe_phv_in_data_297,
  input  [7:0]   io_pipe_phv_in_data_298,
  input  [7:0]   io_pipe_phv_in_data_299,
  input  [7:0]   io_pipe_phv_in_data_300,
  input  [7:0]   io_pipe_phv_in_data_301,
  input  [7:0]   io_pipe_phv_in_data_302,
  input  [7:0]   io_pipe_phv_in_data_303,
  input  [7:0]   io_pipe_phv_in_data_304,
  input  [7:0]   io_pipe_phv_in_data_305,
  input  [7:0]   io_pipe_phv_in_data_306,
  input  [7:0]   io_pipe_phv_in_data_307,
  input  [7:0]   io_pipe_phv_in_data_308,
  input  [7:0]   io_pipe_phv_in_data_309,
  input  [7:0]   io_pipe_phv_in_data_310,
  input  [7:0]   io_pipe_phv_in_data_311,
  input  [7:0]   io_pipe_phv_in_data_312,
  input  [7:0]   io_pipe_phv_in_data_313,
  input  [7:0]   io_pipe_phv_in_data_314,
  input  [7:0]   io_pipe_phv_in_data_315,
  input  [7:0]   io_pipe_phv_in_data_316,
  input  [7:0]   io_pipe_phv_in_data_317,
  input  [7:0]   io_pipe_phv_in_data_318,
  input  [7:0]   io_pipe_phv_in_data_319,
  input  [7:0]   io_pipe_phv_in_data_320,
  input  [7:0]   io_pipe_phv_in_data_321,
  input  [7:0]   io_pipe_phv_in_data_322,
  input  [7:0]   io_pipe_phv_in_data_323,
  input  [7:0]   io_pipe_phv_in_data_324,
  input  [7:0]   io_pipe_phv_in_data_325,
  input  [7:0]   io_pipe_phv_in_data_326,
  input  [7:0]   io_pipe_phv_in_data_327,
  input  [7:0]   io_pipe_phv_in_data_328,
  input  [7:0]   io_pipe_phv_in_data_329,
  input  [7:0]   io_pipe_phv_in_data_330,
  input  [7:0]   io_pipe_phv_in_data_331,
  input  [7:0]   io_pipe_phv_in_data_332,
  input  [7:0]   io_pipe_phv_in_data_333,
  input  [7:0]   io_pipe_phv_in_data_334,
  input  [7:0]   io_pipe_phv_in_data_335,
  input  [7:0]   io_pipe_phv_in_data_336,
  input  [7:0]   io_pipe_phv_in_data_337,
  input  [7:0]   io_pipe_phv_in_data_338,
  input  [7:0]   io_pipe_phv_in_data_339,
  input  [7:0]   io_pipe_phv_in_data_340,
  input  [7:0]   io_pipe_phv_in_data_341,
  input  [7:0]   io_pipe_phv_in_data_342,
  input  [7:0]   io_pipe_phv_in_data_343,
  input  [7:0]   io_pipe_phv_in_data_344,
  input  [7:0]   io_pipe_phv_in_data_345,
  input  [7:0]   io_pipe_phv_in_data_346,
  input  [7:0]   io_pipe_phv_in_data_347,
  input  [7:0]   io_pipe_phv_in_data_348,
  input  [7:0]   io_pipe_phv_in_data_349,
  input  [7:0]   io_pipe_phv_in_data_350,
  input  [7:0]   io_pipe_phv_in_data_351,
  input  [7:0]   io_pipe_phv_in_data_352,
  input  [7:0]   io_pipe_phv_in_data_353,
  input  [7:0]   io_pipe_phv_in_data_354,
  input  [7:0]   io_pipe_phv_in_data_355,
  input  [7:0]   io_pipe_phv_in_data_356,
  input  [7:0]   io_pipe_phv_in_data_357,
  input  [7:0]   io_pipe_phv_in_data_358,
  input  [7:0]   io_pipe_phv_in_data_359,
  input  [7:0]   io_pipe_phv_in_data_360,
  input  [7:0]   io_pipe_phv_in_data_361,
  input  [7:0]   io_pipe_phv_in_data_362,
  input  [7:0]   io_pipe_phv_in_data_363,
  input  [7:0]   io_pipe_phv_in_data_364,
  input  [7:0]   io_pipe_phv_in_data_365,
  input  [7:0]   io_pipe_phv_in_data_366,
  input  [7:0]   io_pipe_phv_in_data_367,
  input  [7:0]   io_pipe_phv_in_data_368,
  input  [7:0]   io_pipe_phv_in_data_369,
  input  [7:0]   io_pipe_phv_in_data_370,
  input  [7:0]   io_pipe_phv_in_data_371,
  input  [7:0]   io_pipe_phv_in_data_372,
  input  [7:0]   io_pipe_phv_in_data_373,
  input  [7:0]   io_pipe_phv_in_data_374,
  input  [7:0]   io_pipe_phv_in_data_375,
  input  [7:0]   io_pipe_phv_in_data_376,
  input  [7:0]   io_pipe_phv_in_data_377,
  input  [7:0]   io_pipe_phv_in_data_378,
  input  [7:0]   io_pipe_phv_in_data_379,
  input  [7:0]   io_pipe_phv_in_data_380,
  input  [7:0]   io_pipe_phv_in_data_381,
  input  [7:0]   io_pipe_phv_in_data_382,
  input  [7:0]   io_pipe_phv_in_data_383,
  input  [7:0]   io_pipe_phv_in_data_384,
  input  [7:0]   io_pipe_phv_in_data_385,
  input  [7:0]   io_pipe_phv_in_data_386,
  input  [7:0]   io_pipe_phv_in_data_387,
  input  [7:0]   io_pipe_phv_in_data_388,
  input  [7:0]   io_pipe_phv_in_data_389,
  input  [7:0]   io_pipe_phv_in_data_390,
  input  [7:0]   io_pipe_phv_in_data_391,
  input  [7:0]   io_pipe_phv_in_data_392,
  input  [7:0]   io_pipe_phv_in_data_393,
  input  [7:0]   io_pipe_phv_in_data_394,
  input  [7:0]   io_pipe_phv_in_data_395,
  input  [7:0]   io_pipe_phv_in_data_396,
  input  [7:0]   io_pipe_phv_in_data_397,
  input  [7:0]   io_pipe_phv_in_data_398,
  input  [7:0]   io_pipe_phv_in_data_399,
  input  [7:0]   io_pipe_phv_in_data_400,
  input  [7:0]   io_pipe_phv_in_data_401,
  input  [7:0]   io_pipe_phv_in_data_402,
  input  [7:0]   io_pipe_phv_in_data_403,
  input  [7:0]   io_pipe_phv_in_data_404,
  input  [7:0]   io_pipe_phv_in_data_405,
  input  [7:0]   io_pipe_phv_in_data_406,
  input  [7:0]   io_pipe_phv_in_data_407,
  input  [7:0]   io_pipe_phv_in_data_408,
  input  [7:0]   io_pipe_phv_in_data_409,
  input  [7:0]   io_pipe_phv_in_data_410,
  input  [7:0]   io_pipe_phv_in_data_411,
  input  [7:0]   io_pipe_phv_in_data_412,
  input  [7:0]   io_pipe_phv_in_data_413,
  input  [7:0]   io_pipe_phv_in_data_414,
  input  [7:0]   io_pipe_phv_in_data_415,
  input  [7:0]   io_pipe_phv_in_data_416,
  input  [7:0]   io_pipe_phv_in_data_417,
  input  [7:0]   io_pipe_phv_in_data_418,
  input  [7:0]   io_pipe_phv_in_data_419,
  input  [7:0]   io_pipe_phv_in_data_420,
  input  [7:0]   io_pipe_phv_in_data_421,
  input  [7:0]   io_pipe_phv_in_data_422,
  input  [7:0]   io_pipe_phv_in_data_423,
  input  [7:0]   io_pipe_phv_in_data_424,
  input  [7:0]   io_pipe_phv_in_data_425,
  input  [7:0]   io_pipe_phv_in_data_426,
  input  [7:0]   io_pipe_phv_in_data_427,
  input  [7:0]   io_pipe_phv_in_data_428,
  input  [7:0]   io_pipe_phv_in_data_429,
  input  [7:0]   io_pipe_phv_in_data_430,
  input  [7:0]   io_pipe_phv_in_data_431,
  input  [7:0]   io_pipe_phv_in_data_432,
  input  [7:0]   io_pipe_phv_in_data_433,
  input  [7:0]   io_pipe_phv_in_data_434,
  input  [7:0]   io_pipe_phv_in_data_435,
  input  [7:0]   io_pipe_phv_in_data_436,
  input  [7:0]   io_pipe_phv_in_data_437,
  input  [7:0]   io_pipe_phv_in_data_438,
  input  [7:0]   io_pipe_phv_in_data_439,
  input  [7:0]   io_pipe_phv_in_data_440,
  input  [7:0]   io_pipe_phv_in_data_441,
  input  [7:0]   io_pipe_phv_in_data_442,
  input  [7:0]   io_pipe_phv_in_data_443,
  input  [7:0]   io_pipe_phv_in_data_444,
  input  [7:0]   io_pipe_phv_in_data_445,
  input  [7:0]   io_pipe_phv_in_data_446,
  input  [7:0]   io_pipe_phv_in_data_447,
  input  [7:0]   io_pipe_phv_in_data_448,
  input  [7:0]   io_pipe_phv_in_data_449,
  input  [7:0]   io_pipe_phv_in_data_450,
  input  [7:0]   io_pipe_phv_in_data_451,
  input  [7:0]   io_pipe_phv_in_data_452,
  input  [7:0]   io_pipe_phv_in_data_453,
  input  [7:0]   io_pipe_phv_in_data_454,
  input  [7:0]   io_pipe_phv_in_data_455,
  input  [7:0]   io_pipe_phv_in_data_456,
  input  [7:0]   io_pipe_phv_in_data_457,
  input  [7:0]   io_pipe_phv_in_data_458,
  input  [7:0]   io_pipe_phv_in_data_459,
  input  [7:0]   io_pipe_phv_in_data_460,
  input  [7:0]   io_pipe_phv_in_data_461,
  input  [7:0]   io_pipe_phv_in_data_462,
  input  [7:0]   io_pipe_phv_in_data_463,
  input  [7:0]   io_pipe_phv_in_data_464,
  input  [7:0]   io_pipe_phv_in_data_465,
  input  [7:0]   io_pipe_phv_in_data_466,
  input  [7:0]   io_pipe_phv_in_data_467,
  input  [7:0]   io_pipe_phv_in_data_468,
  input  [7:0]   io_pipe_phv_in_data_469,
  input  [7:0]   io_pipe_phv_in_data_470,
  input  [7:0]   io_pipe_phv_in_data_471,
  input  [7:0]   io_pipe_phv_in_data_472,
  input  [7:0]   io_pipe_phv_in_data_473,
  input  [7:0]   io_pipe_phv_in_data_474,
  input  [7:0]   io_pipe_phv_in_data_475,
  input  [7:0]   io_pipe_phv_in_data_476,
  input  [7:0]   io_pipe_phv_in_data_477,
  input  [7:0]   io_pipe_phv_in_data_478,
  input  [7:0]   io_pipe_phv_in_data_479,
  input  [7:0]   io_pipe_phv_in_data_480,
  input  [7:0]   io_pipe_phv_in_data_481,
  input  [7:0]   io_pipe_phv_in_data_482,
  input  [7:0]   io_pipe_phv_in_data_483,
  input  [7:0]   io_pipe_phv_in_data_484,
  input  [7:0]   io_pipe_phv_in_data_485,
  input  [7:0]   io_pipe_phv_in_data_486,
  input  [7:0]   io_pipe_phv_in_data_487,
  input  [7:0]   io_pipe_phv_in_data_488,
  input  [7:0]   io_pipe_phv_in_data_489,
  input  [7:0]   io_pipe_phv_in_data_490,
  input  [7:0]   io_pipe_phv_in_data_491,
  input  [7:0]   io_pipe_phv_in_data_492,
  input  [7:0]   io_pipe_phv_in_data_493,
  input  [7:0]   io_pipe_phv_in_data_494,
  input  [7:0]   io_pipe_phv_in_data_495,
  input  [7:0]   io_pipe_phv_in_data_496,
  input  [7:0]   io_pipe_phv_in_data_497,
  input  [7:0]   io_pipe_phv_in_data_498,
  input  [7:0]   io_pipe_phv_in_data_499,
  input  [7:0]   io_pipe_phv_in_data_500,
  input  [7:0]   io_pipe_phv_in_data_501,
  input  [7:0]   io_pipe_phv_in_data_502,
  input  [7:0]   io_pipe_phv_in_data_503,
  input  [7:0]   io_pipe_phv_in_data_504,
  input  [7:0]   io_pipe_phv_in_data_505,
  input  [7:0]   io_pipe_phv_in_data_506,
  input  [7:0]   io_pipe_phv_in_data_507,
  input  [7:0]   io_pipe_phv_in_data_508,
  input  [7:0]   io_pipe_phv_in_data_509,
  input  [7:0]   io_pipe_phv_in_data_510,
  input  [7:0]   io_pipe_phv_in_data_511,
  input  [3:0]   io_pipe_phv_in_next_processor_id,
  input          io_pipe_phv_in_next_config_id,
  input          io_pipe_phv_in_is_valid_processor,
  output [7:0]   io_pipe_phv_out_data_0,
  output [7:0]   io_pipe_phv_out_data_1,
  output [7:0]   io_pipe_phv_out_data_2,
  output [7:0]   io_pipe_phv_out_data_3,
  output [7:0]   io_pipe_phv_out_data_4,
  output [7:0]   io_pipe_phv_out_data_5,
  output [7:0]   io_pipe_phv_out_data_6,
  output [7:0]   io_pipe_phv_out_data_7,
  output [7:0]   io_pipe_phv_out_data_8,
  output [7:0]   io_pipe_phv_out_data_9,
  output [7:0]   io_pipe_phv_out_data_10,
  output [7:0]   io_pipe_phv_out_data_11,
  output [7:0]   io_pipe_phv_out_data_12,
  output [7:0]   io_pipe_phv_out_data_13,
  output [7:0]   io_pipe_phv_out_data_14,
  output [7:0]   io_pipe_phv_out_data_15,
  output [7:0]   io_pipe_phv_out_data_16,
  output [7:0]   io_pipe_phv_out_data_17,
  output [7:0]   io_pipe_phv_out_data_18,
  output [7:0]   io_pipe_phv_out_data_19,
  output [7:0]   io_pipe_phv_out_data_20,
  output [7:0]   io_pipe_phv_out_data_21,
  output [7:0]   io_pipe_phv_out_data_22,
  output [7:0]   io_pipe_phv_out_data_23,
  output [7:0]   io_pipe_phv_out_data_24,
  output [7:0]   io_pipe_phv_out_data_25,
  output [7:0]   io_pipe_phv_out_data_26,
  output [7:0]   io_pipe_phv_out_data_27,
  output [7:0]   io_pipe_phv_out_data_28,
  output [7:0]   io_pipe_phv_out_data_29,
  output [7:0]   io_pipe_phv_out_data_30,
  output [7:0]   io_pipe_phv_out_data_31,
  output [7:0]   io_pipe_phv_out_data_32,
  output [7:0]   io_pipe_phv_out_data_33,
  output [7:0]   io_pipe_phv_out_data_34,
  output [7:0]   io_pipe_phv_out_data_35,
  output [7:0]   io_pipe_phv_out_data_36,
  output [7:0]   io_pipe_phv_out_data_37,
  output [7:0]   io_pipe_phv_out_data_38,
  output [7:0]   io_pipe_phv_out_data_39,
  output [7:0]   io_pipe_phv_out_data_40,
  output [7:0]   io_pipe_phv_out_data_41,
  output [7:0]   io_pipe_phv_out_data_42,
  output [7:0]   io_pipe_phv_out_data_43,
  output [7:0]   io_pipe_phv_out_data_44,
  output [7:0]   io_pipe_phv_out_data_45,
  output [7:0]   io_pipe_phv_out_data_46,
  output [7:0]   io_pipe_phv_out_data_47,
  output [7:0]   io_pipe_phv_out_data_48,
  output [7:0]   io_pipe_phv_out_data_49,
  output [7:0]   io_pipe_phv_out_data_50,
  output [7:0]   io_pipe_phv_out_data_51,
  output [7:0]   io_pipe_phv_out_data_52,
  output [7:0]   io_pipe_phv_out_data_53,
  output [7:0]   io_pipe_phv_out_data_54,
  output [7:0]   io_pipe_phv_out_data_55,
  output [7:0]   io_pipe_phv_out_data_56,
  output [7:0]   io_pipe_phv_out_data_57,
  output [7:0]   io_pipe_phv_out_data_58,
  output [7:0]   io_pipe_phv_out_data_59,
  output [7:0]   io_pipe_phv_out_data_60,
  output [7:0]   io_pipe_phv_out_data_61,
  output [7:0]   io_pipe_phv_out_data_62,
  output [7:0]   io_pipe_phv_out_data_63,
  output [7:0]   io_pipe_phv_out_data_64,
  output [7:0]   io_pipe_phv_out_data_65,
  output [7:0]   io_pipe_phv_out_data_66,
  output [7:0]   io_pipe_phv_out_data_67,
  output [7:0]   io_pipe_phv_out_data_68,
  output [7:0]   io_pipe_phv_out_data_69,
  output [7:0]   io_pipe_phv_out_data_70,
  output [7:0]   io_pipe_phv_out_data_71,
  output [7:0]   io_pipe_phv_out_data_72,
  output [7:0]   io_pipe_phv_out_data_73,
  output [7:0]   io_pipe_phv_out_data_74,
  output [7:0]   io_pipe_phv_out_data_75,
  output [7:0]   io_pipe_phv_out_data_76,
  output [7:0]   io_pipe_phv_out_data_77,
  output [7:0]   io_pipe_phv_out_data_78,
  output [7:0]   io_pipe_phv_out_data_79,
  output [7:0]   io_pipe_phv_out_data_80,
  output [7:0]   io_pipe_phv_out_data_81,
  output [7:0]   io_pipe_phv_out_data_82,
  output [7:0]   io_pipe_phv_out_data_83,
  output [7:0]   io_pipe_phv_out_data_84,
  output [7:0]   io_pipe_phv_out_data_85,
  output [7:0]   io_pipe_phv_out_data_86,
  output [7:0]   io_pipe_phv_out_data_87,
  output [7:0]   io_pipe_phv_out_data_88,
  output [7:0]   io_pipe_phv_out_data_89,
  output [7:0]   io_pipe_phv_out_data_90,
  output [7:0]   io_pipe_phv_out_data_91,
  output [7:0]   io_pipe_phv_out_data_92,
  output [7:0]   io_pipe_phv_out_data_93,
  output [7:0]   io_pipe_phv_out_data_94,
  output [7:0]   io_pipe_phv_out_data_95,
  output [7:0]   io_pipe_phv_out_data_96,
  output [7:0]   io_pipe_phv_out_data_97,
  output [7:0]   io_pipe_phv_out_data_98,
  output [7:0]   io_pipe_phv_out_data_99,
  output [7:0]   io_pipe_phv_out_data_100,
  output [7:0]   io_pipe_phv_out_data_101,
  output [7:0]   io_pipe_phv_out_data_102,
  output [7:0]   io_pipe_phv_out_data_103,
  output [7:0]   io_pipe_phv_out_data_104,
  output [7:0]   io_pipe_phv_out_data_105,
  output [7:0]   io_pipe_phv_out_data_106,
  output [7:0]   io_pipe_phv_out_data_107,
  output [7:0]   io_pipe_phv_out_data_108,
  output [7:0]   io_pipe_phv_out_data_109,
  output [7:0]   io_pipe_phv_out_data_110,
  output [7:0]   io_pipe_phv_out_data_111,
  output [7:0]   io_pipe_phv_out_data_112,
  output [7:0]   io_pipe_phv_out_data_113,
  output [7:0]   io_pipe_phv_out_data_114,
  output [7:0]   io_pipe_phv_out_data_115,
  output [7:0]   io_pipe_phv_out_data_116,
  output [7:0]   io_pipe_phv_out_data_117,
  output [7:0]   io_pipe_phv_out_data_118,
  output [7:0]   io_pipe_phv_out_data_119,
  output [7:0]   io_pipe_phv_out_data_120,
  output [7:0]   io_pipe_phv_out_data_121,
  output [7:0]   io_pipe_phv_out_data_122,
  output [7:0]   io_pipe_phv_out_data_123,
  output [7:0]   io_pipe_phv_out_data_124,
  output [7:0]   io_pipe_phv_out_data_125,
  output [7:0]   io_pipe_phv_out_data_126,
  output [7:0]   io_pipe_phv_out_data_127,
  output [7:0]   io_pipe_phv_out_data_128,
  output [7:0]   io_pipe_phv_out_data_129,
  output [7:0]   io_pipe_phv_out_data_130,
  output [7:0]   io_pipe_phv_out_data_131,
  output [7:0]   io_pipe_phv_out_data_132,
  output [7:0]   io_pipe_phv_out_data_133,
  output [7:0]   io_pipe_phv_out_data_134,
  output [7:0]   io_pipe_phv_out_data_135,
  output [7:0]   io_pipe_phv_out_data_136,
  output [7:0]   io_pipe_phv_out_data_137,
  output [7:0]   io_pipe_phv_out_data_138,
  output [7:0]   io_pipe_phv_out_data_139,
  output [7:0]   io_pipe_phv_out_data_140,
  output [7:0]   io_pipe_phv_out_data_141,
  output [7:0]   io_pipe_phv_out_data_142,
  output [7:0]   io_pipe_phv_out_data_143,
  output [7:0]   io_pipe_phv_out_data_144,
  output [7:0]   io_pipe_phv_out_data_145,
  output [7:0]   io_pipe_phv_out_data_146,
  output [7:0]   io_pipe_phv_out_data_147,
  output [7:0]   io_pipe_phv_out_data_148,
  output [7:0]   io_pipe_phv_out_data_149,
  output [7:0]   io_pipe_phv_out_data_150,
  output [7:0]   io_pipe_phv_out_data_151,
  output [7:0]   io_pipe_phv_out_data_152,
  output [7:0]   io_pipe_phv_out_data_153,
  output [7:0]   io_pipe_phv_out_data_154,
  output [7:0]   io_pipe_phv_out_data_155,
  output [7:0]   io_pipe_phv_out_data_156,
  output [7:0]   io_pipe_phv_out_data_157,
  output [7:0]   io_pipe_phv_out_data_158,
  output [7:0]   io_pipe_phv_out_data_159,
  output [7:0]   io_pipe_phv_out_data_160,
  output [7:0]   io_pipe_phv_out_data_161,
  output [7:0]   io_pipe_phv_out_data_162,
  output [7:0]   io_pipe_phv_out_data_163,
  output [7:0]   io_pipe_phv_out_data_164,
  output [7:0]   io_pipe_phv_out_data_165,
  output [7:0]   io_pipe_phv_out_data_166,
  output [7:0]   io_pipe_phv_out_data_167,
  output [7:0]   io_pipe_phv_out_data_168,
  output [7:0]   io_pipe_phv_out_data_169,
  output [7:0]   io_pipe_phv_out_data_170,
  output [7:0]   io_pipe_phv_out_data_171,
  output [7:0]   io_pipe_phv_out_data_172,
  output [7:0]   io_pipe_phv_out_data_173,
  output [7:0]   io_pipe_phv_out_data_174,
  output [7:0]   io_pipe_phv_out_data_175,
  output [7:0]   io_pipe_phv_out_data_176,
  output [7:0]   io_pipe_phv_out_data_177,
  output [7:0]   io_pipe_phv_out_data_178,
  output [7:0]   io_pipe_phv_out_data_179,
  output [7:0]   io_pipe_phv_out_data_180,
  output [7:0]   io_pipe_phv_out_data_181,
  output [7:0]   io_pipe_phv_out_data_182,
  output [7:0]   io_pipe_phv_out_data_183,
  output [7:0]   io_pipe_phv_out_data_184,
  output [7:0]   io_pipe_phv_out_data_185,
  output [7:0]   io_pipe_phv_out_data_186,
  output [7:0]   io_pipe_phv_out_data_187,
  output [7:0]   io_pipe_phv_out_data_188,
  output [7:0]   io_pipe_phv_out_data_189,
  output [7:0]   io_pipe_phv_out_data_190,
  output [7:0]   io_pipe_phv_out_data_191,
  output [7:0]   io_pipe_phv_out_data_192,
  output [7:0]   io_pipe_phv_out_data_193,
  output [7:0]   io_pipe_phv_out_data_194,
  output [7:0]   io_pipe_phv_out_data_195,
  output [7:0]   io_pipe_phv_out_data_196,
  output [7:0]   io_pipe_phv_out_data_197,
  output [7:0]   io_pipe_phv_out_data_198,
  output [7:0]   io_pipe_phv_out_data_199,
  output [7:0]   io_pipe_phv_out_data_200,
  output [7:0]   io_pipe_phv_out_data_201,
  output [7:0]   io_pipe_phv_out_data_202,
  output [7:0]   io_pipe_phv_out_data_203,
  output [7:0]   io_pipe_phv_out_data_204,
  output [7:0]   io_pipe_phv_out_data_205,
  output [7:0]   io_pipe_phv_out_data_206,
  output [7:0]   io_pipe_phv_out_data_207,
  output [7:0]   io_pipe_phv_out_data_208,
  output [7:0]   io_pipe_phv_out_data_209,
  output [7:0]   io_pipe_phv_out_data_210,
  output [7:0]   io_pipe_phv_out_data_211,
  output [7:0]   io_pipe_phv_out_data_212,
  output [7:0]   io_pipe_phv_out_data_213,
  output [7:0]   io_pipe_phv_out_data_214,
  output [7:0]   io_pipe_phv_out_data_215,
  output [7:0]   io_pipe_phv_out_data_216,
  output [7:0]   io_pipe_phv_out_data_217,
  output [7:0]   io_pipe_phv_out_data_218,
  output [7:0]   io_pipe_phv_out_data_219,
  output [7:0]   io_pipe_phv_out_data_220,
  output [7:0]   io_pipe_phv_out_data_221,
  output [7:0]   io_pipe_phv_out_data_222,
  output [7:0]   io_pipe_phv_out_data_223,
  output [7:0]   io_pipe_phv_out_data_224,
  output [7:0]   io_pipe_phv_out_data_225,
  output [7:0]   io_pipe_phv_out_data_226,
  output [7:0]   io_pipe_phv_out_data_227,
  output [7:0]   io_pipe_phv_out_data_228,
  output [7:0]   io_pipe_phv_out_data_229,
  output [7:0]   io_pipe_phv_out_data_230,
  output [7:0]   io_pipe_phv_out_data_231,
  output [7:0]   io_pipe_phv_out_data_232,
  output [7:0]   io_pipe_phv_out_data_233,
  output [7:0]   io_pipe_phv_out_data_234,
  output [7:0]   io_pipe_phv_out_data_235,
  output [7:0]   io_pipe_phv_out_data_236,
  output [7:0]   io_pipe_phv_out_data_237,
  output [7:0]   io_pipe_phv_out_data_238,
  output [7:0]   io_pipe_phv_out_data_239,
  output [7:0]   io_pipe_phv_out_data_240,
  output [7:0]   io_pipe_phv_out_data_241,
  output [7:0]   io_pipe_phv_out_data_242,
  output [7:0]   io_pipe_phv_out_data_243,
  output [7:0]   io_pipe_phv_out_data_244,
  output [7:0]   io_pipe_phv_out_data_245,
  output [7:0]   io_pipe_phv_out_data_246,
  output [7:0]   io_pipe_phv_out_data_247,
  output [7:0]   io_pipe_phv_out_data_248,
  output [7:0]   io_pipe_phv_out_data_249,
  output [7:0]   io_pipe_phv_out_data_250,
  output [7:0]   io_pipe_phv_out_data_251,
  output [7:0]   io_pipe_phv_out_data_252,
  output [7:0]   io_pipe_phv_out_data_253,
  output [7:0]   io_pipe_phv_out_data_254,
  output [7:0]   io_pipe_phv_out_data_255,
  output [7:0]   io_pipe_phv_out_data_256,
  output [7:0]   io_pipe_phv_out_data_257,
  output [7:0]   io_pipe_phv_out_data_258,
  output [7:0]   io_pipe_phv_out_data_259,
  output [7:0]   io_pipe_phv_out_data_260,
  output [7:0]   io_pipe_phv_out_data_261,
  output [7:0]   io_pipe_phv_out_data_262,
  output [7:0]   io_pipe_phv_out_data_263,
  output [7:0]   io_pipe_phv_out_data_264,
  output [7:0]   io_pipe_phv_out_data_265,
  output [7:0]   io_pipe_phv_out_data_266,
  output [7:0]   io_pipe_phv_out_data_267,
  output [7:0]   io_pipe_phv_out_data_268,
  output [7:0]   io_pipe_phv_out_data_269,
  output [7:0]   io_pipe_phv_out_data_270,
  output [7:0]   io_pipe_phv_out_data_271,
  output [7:0]   io_pipe_phv_out_data_272,
  output [7:0]   io_pipe_phv_out_data_273,
  output [7:0]   io_pipe_phv_out_data_274,
  output [7:0]   io_pipe_phv_out_data_275,
  output [7:0]   io_pipe_phv_out_data_276,
  output [7:0]   io_pipe_phv_out_data_277,
  output [7:0]   io_pipe_phv_out_data_278,
  output [7:0]   io_pipe_phv_out_data_279,
  output [7:0]   io_pipe_phv_out_data_280,
  output [7:0]   io_pipe_phv_out_data_281,
  output [7:0]   io_pipe_phv_out_data_282,
  output [7:0]   io_pipe_phv_out_data_283,
  output [7:0]   io_pipe_phv_out_data_284,
  output [7:0]   io_pipe_phv_out_data_285,
  output [7:0]   io_pipe_phv_out_data_286,
  output [7:0]   io_pipe_phv_out_data_287,
  output [7:0]   io_pipe_phv_out_data_288,
  output [7:0]   io_pipe_phv_out_data_289,
  output [7:0]   io_pipe_phv_out_data_290,
  output [7:0]   io_pipe_phv_out_data_291,
  output [7:0]   io_pipe_phv_out_data_292,
  output [7:0]   io_pipe_phv_out_data_293,
  output [7:0]   io_pipe_phv_out_data_294,
  output [7:0]   io_pipe_phv_out_data_295,
  output [7:0]   io_pipe_phv_out_data_296,
  output [7:0]   io_pipe_phv_out_data_297,
  output [7:0]   io_pipe_phv_out_data_298,
  output [7:0]   io_pipe_phv_out_data_299,
  output [7:0]   io_pipe_phv_out_data_300,
  output [7:0]   io_pipe_phv_out_data_301,
  output [7:0]   io_pipe_phv_out_data_302,
  output [7:0]   io_pipe_phv_out_data_303,
  output [7:0]   io_pipe_phv_out_data_304,
  output [7:0]   io_pipe_phv_out_data_305,
  output [7:0]   io_pipe_phv_out_data_306,
  output [7:0]   io_pipe_phv_out_data_307,
  output [7:0]   io_pipe_phv_out_data_308,
  output [7:0]   io_pipe_phv_out_data_309,
  output [7:0]   io_pipe_phv_out_data_310,
  output [7:0]   io_pipe_phv_out_data_311,
  output [7:0]   io_pipe_phv_out_data_312,
  output [7:0]   io_pipe_phv_out_data_313,
  output [7:0]   io_pipe_phv_out_data_314,
  output [7:0]   io_pipe_phv_out_data_315,
  output [7:0]   io_pipe_phv_out_data_316,
  output [7:0]   io_pipe_phv_out_data_317,
  output [7:0]   io_pipe_phv_out_data_318,
  output [7:0]   io_pipe_phv_out_data_319,
  output [7:0]   io_pipe_phv_out_data_320,
  output [7:0]   io_pipe_phv_out_data_321,
  output [7:0]   io_pipe_phv_out_data_322,
  output [7:0]   io_pipe_phv_out_data_323,
  output [7:0]   io_pipe_phv_out_data_324,
  output [7:0]   io_pipe_phv_out_data_325,
  output [7:0]   io_pipe_phv_out_data_326,
  output [7:0]   io_pipe_phv_out_data_327,
  output [7:0]   io_pipe_phv_out_data_328,
  output [7:0]   io_pipe_phv_out_data_329,
  output [7:0]   io_pipe_phv_out_data_330,
  output [7:0]   io_pipe_phv_out_data_331,
  output [7:0]   io_pipe_phv_out_data_332,
  output [7:0]   io_pipe_phv_out_data_333,
  output [7:0]   io_pipe_phv_out_data_334,
  output [7:0]   io_pipe_phv_out_data_335,
  output [7:0]   io_pipe_phv_out_data_336,
  output [7:0]   io_pipe_phv_out_data_337,
  output [7:0]   io_pipe_phv_out_data_338,
  output [7:0]   io_pipe_phv_out_data_339,
  output [7:0]   io_pipe_phv_out_data_340,
  output [7:0]   io_pipe_phv_out_data_341,
  output [7:0]   io_pipe_phv_out_data_342,
  output [7:0]   io_pipe_phv_out_data_343,
  output [7:0]   io_pipe_phv_out_data_344,
  output [7:0]   io_pipe_phv_out_data_345,
  output [7:0]   io_pipe_phv_out_data_346,
  output [7:0]   io_pipe_phv_out_data_347,
  output [7:0]   io_pipe_phv_out_data_348,
  output [7:0]   io_pipe_phv_out_data_349,
  output [7:0]   io_pipe_phv_out_data_350,
  output [7:0]   io_pipe_phv_out_data_351,
  output [7:0]   io_pipe_phv_out_data_352,
  output [7:0]   io_pipe_phv_out_data_353,
  output [7:0]   io_pipe_phv_out_data_354,
  output [7:0]   io_pipe_phv_out_data_355,
  output [7:0]   io_pipe_phv_out_data_356,
  output [7:0]   io_pipe_phv_out_data_357,
  output [7:0]   io_pipe_phv_out_data_358,
  output [7:0]   io_pipe_phv_out_data_359,
  output [7:0]   io_pipe_phv_out_data_360,
  output [7:0]   io_pipe_phv_out_data_361,
  output [7:0]   io_pipe_phv_out_data_362,
  output [7:0]   io_pipe_phv_out_data_363,
  output [7:0]   io_pipe_phv_out_data_364,
  output [7:0]   io_pipe_phv_out_data_365,
  output [7:0]   io_pipe_phv_out_data_366,
  output [7:0]   io_pipe_phv_out_data_367,
  output [7:0]   io_pipe_phv_out_data_368,
  output [7:0]   io_pipe_phv_out_data_369,
  output [7:0]   io_pipe_phv_out_data_370,
  output [7:0]   io_pipe_phv_out_data_371,
  output [7:0]   io_pipe_phv_out_data_372,
  output [7:0]   io_pipe_phv_out_data_373,
  output [7:0]   io_pipe_phv_out_data_374,
  output [7:0]   io_pipe_phv_out_data_375,
  output [7:0]   io_pipe_phv_out_data_376,
  output [7:0]   io_pipe_phv_out_data_377,
  output [7:0]   io_pipe_phv_out_data_378,
  output [7:0]   io_pipe_phv_out_data_379,
  output [7:0]   io_pipe_phv_out_data_380,
  output [7:0]   io_pipe_phv_out_data_381,
  output [7:0]   io_pipe_phv_out_data_382,
  output [7:0]   io_pipe_phv_out_data_383,
  output [7:0]   io_pipe_phv_out_data_384,
  output [7:0]   io_pipe_phv_out_data_385,
  output [7:0]   io_pipe_phv_out_data_386,
  output [7:0]   io_pipe_phv_out_data_387,
  output [7:0]   io_pipe_phv_out_data_388,
  output [7:0]   io_pipe_phv_out_data_389,
  output [7:0]   io_pipe_phv_out_data_390,
  output [7:0]   io_pipe_phv_out_data_391,
  output [7:0]   io_pipe_phv_out_data_392,
  output [7:0]   io_pipe_phv_out_data_393,
  output [7:0]   io_pipe_phv_out_data_394,
  output [7:0]   io_pipe_phv_out_data_395,
  output [7:0]   io_pipe_phv_out_data_396,
  output [7:0]   io_pipe_phv_out_data_397,
  output [7:0]   io_pipe_phv_out_data_398,
  output [7:0]   io_pipe_phv_out_data_399,
  output [7:0]   io_pipe_phv_out_data_400,
  output [7:0]   io_pipe_phv_out_data_401,
  output [7:0]   io_pipe_phv_out_data_402,
  output [7:0]   io_pipe_phv_out_data_403,
  output [7:0]   io_pipe_phv_out_data_404,
  output [7:0]   io_pipe_phv_out_data_405,
  output [7:0]   io_pipe_phv_out_data_406,
  output [7:0]   io_pipe_phv_out_data_407,
  output [7:0]   io_pipe_phv_out_data_408,
  output [7:0]   io_pipe_phv_out_data_409,
  output [7:0]   io_pipe_phv_out_data_410,
  output [7:0]   io_pipe_phv_out_data_411,
  output [7:0]   io_pipe_phv_out_data_412,
  output [7:0]   io_pipe_phv_out_data_413,
  output [7:0]   io_pipe_phv_out_data_414,
  output [7:0]   io_pipe_phv_out_data_415,
  output [7:0]   io_pipe_phv_out_data_416,
  output [7:0]   io_pipe_phv_out_data_417,
  output [7:0]   io_pipe_phv_out_data_418,
  output [7:0]   io_pipe_phv_out_data_419,
  output [7:0]   io_pipe_phv_out_data_420,
  output [7:0]   io_pipe_phv_out_data_421,
  output [7:0]   io_pipe_phv_out_data_422,
  output [7:0]   io_pipe_phv_out_data_423,
  output [7:0]   io_pipe_phv_out_data_424,
  output [7:0]   io_pipe_phv_out_data_425,
  output [7:0]   io_pipe_phv_out_data_426,
  output [7:0]   io_pipe_phv_out_data_427,
  output [7:0]   io_pipe_phv_out_data_428,
  output [7:0]   io_pipe_phv_out_data_429,
  output [7:0]   io_pipe_phv_out_data_430,
  output [7:0]   io_pipe_phv_out_data_431,
  output [7:0]   io_pipe_phv_out_data_432,
  output [7:0]   io_pipe_phv_out_data_433,
  output [7:0]   io_pipe_phv_out_data_434,
  output [7:0]   io_pipe_phv_out_data_435,
  output [7:0]   io_pipe_phv_out_data_436,
  output [7:0]   io_pipe_phv_out_data_437,
  output [7:0]   io_pipe_phv_out_data_438,
  output [7:0]   io_pipe_phv_out_data_439,
  output [7:0]   io_pipe_phv_out_data_440,
  output [7:0]   io_pipe_phv_out_data_441,
  output [7:0]   io_pipe_phv_out_data_442,
  output [7:0]   io_pipe_phv_out_data_443,
  output [7:0]   io_pipe_phv_out_data_444,
  output [7:0]   io_pipe_phv_out_data_445,
  output [7:0]   io_pipe_phv_out_data_446,
  output [7:0]   io_pipe_phv_out_data_447,
  output [7:0]   io_pipe_phv_out_data_448,
  output [7:0]   io_pipe_phv_out_data_449,
  output [7:0]   io_pipe_phv_out_data_450,
  output [7:0]   io_pipe_phv_out_data_451,
  output [7:0]   io_pipe_phv_out_data_452,
  output [7:0]   io_pipe_phv_out_data_453,
  output [7:0]   io_pipe_phv_out_data_454,
  output [7:0]   io_pipe_phv_out_data_455,
  output [7:0]   io_pipe_phv_out_data_456,
  output [7:0]   io_pipe_phv_out_data_457,
  output [7:0]   io_pipe_phv_out_data_458,
  output [7:0]   io_pipe_phv_out_data_459,
  output [7:0]   io_pipe_phv_out_data_460,
  output [7:0]   io_pipe_phv_out_data_461,
  output [7:0]   io_pipe_phv_out_data_462,
  output [7:0]   io_pipe_phv_out_data_463,
  output [7:0]   io_pipe_phv_out_data_464,
  output [7:0]   io_pipe_phv_out_data_465,
  output [7:0]   io_pipe_phv_out_data_466,
  output [7:0]   io_pipe_phv_out_data_467,
  output [7:0]   io_pipe_phv_out_data_468,
  output [7:0]   io_pipe_phv_out_data_469,
  output [7:0]   io_pipe_phv_out_data_470,
  output [7:0]   io_pipe_phv_out_data_471,
  output [7:0]   io_pipe_phv_out_data_472,
  output [7:0]   io_pipe_phv_out_data_473,
  output [7:0]   io_pipe_phv_out_data_474,
  output [7:0]   io_pipe_phv_out_data_475,
  output [7:0]   io_pipe_phv_out_data_476,
  output [7:0]   io_pipe_phv_out_data_477,
  output [7:0]   io_pipe_phv_out_data_478,
  output [7:0]   io_pipe_phv_out_data_479,
  output [7:0]   io_pipe_phv_out_data_480,
  output [7:0]   io_pipe_phv_out_data_481,
  output [7:0]   io_pipe_phv_out_data_482,
  output [7:0]   io_pipe_phv_out_data_483,
  output [7:0]   io_pipe_phv_out_data_484,
  output [7:0]   io_pipe_phv_out_data_485,
  output [7:0]   io_pipe_phv_out_data_486,
  output [7:0]   io_pipe_phv_out_data_487,
  output [7:0]   io_pipe_phv_out_data_488,
  output [7:0]   io_pipe_phv_out_data_489,
  output [7:0]   io_pipe_phv_out_data_490,
  output [7:0]   io_pipe_phv_out_data_491,
  output [7:0]   io_pipe_phv_out_data_492,
  output [7:0]   io_pipe_phv_out_data_493,
  output [7:0]   io_pipe_phv_out_data_494,
  output [7:0]   io_pipe_phv_out_data_495,
  output [7:0]   io_pipe_phv_out_data_496,
  output [7:0]   io_pipe_phv_out_data_497,
  output [7:0]   io_pipe_phv_out_data_498,
  output [7:0]   io_pipe_phv_out_data_499,
  output [7:0]   io_pipe_phv_out_data_500,
  output [7:0]   io_pipe_phv_out_data_501,
  output [7:0]   io_pipe_phv_out_data_502,
  output [7:0]   io_pipe_phv_out_data_503,
  output [7:0]   io_pipe_phv_out_data_504,
  output [7:0]   io_pipe_phv_out_data_505,
  output [7:0]   io_pipe_phv_out_data_506,
  output [7:0]   io_pipe_phv_out_data_507,
  output [7:0]   io_pipe_phv_out_data_508,
  output [7:0]   io_pipe_phv_out_data_509,
  output [7:0]   io_pipe_phv_out_data_510,
  output [7:0]   io_pipe_phv_out_data_511,
  output [3:0]   io_pipe_phv_out_next_processor_id,
  output         io_pipe_phv_out_next_config_id,
  output         io_pipe_phv_out_is_valid_processor,
  input  [1:0]   io_key_config_0_field_config_0,
  input  [1:0]   io_key_config_0_field_config_1,
  input  [1:0]   io_key_config_0_field_config_2,
  input  [1:0]   io_key_config_0_field_config_3,
  input  [1:0]   io_key_config_0_field_config_4,
  input  [1:0]   io_key_config_0_field_config_5,
  input          io_key_config_0_field_mask_0_0,
  input          io_key_config_0_field_mask_0_1,
  input          io_key_config_0_field_mask_0_2,
  input          io_key_config_0_field_mask_0_3,
  input          io_key_config_0_field_mask_1_0,
  input          io_key_config_0_field_mask_1_1,
  input          io_key_config_0_field_mask_1_2,
  input          io_key_config_0_field_mask_1_3,
  input          io_key_config_0_field_mask_2_0,
  input          io_key_config_0_field_mask_2_1,
  input          io_key_config_0_field_mask_2_2,
  input          io_key_config_0_field_mask_2_3,
  input          io_key_config_0_field_mask_3_0,
  input          io_key_config_0_field_mask_3_1,
  input          io_key_config_0_field_mask_3_2,
  input          io_key_config_0_field_mask_3_3,
  input          io_key_config_0_field_mask_4_0,
  input          io_key_config_0_field_mask_4_1,
  input          io_key_config_0_field_mask_4_2,
  input          io_key_config_0_field_mask_4_3,
  input          io_key_config_0_field_mask_5_0,
  input          io_key_config_0_field_mask_5_1,
  input          io_key_config_0_field_mask_5_2,
  input          io_key_config_0_field_mask_5_3,
  input  [7:0]   io_key_config_0_field_id_0_0,
  input  [7:0]   io_key_config_0_field_id_0_1,
  input  [7:0]   io_key_config_0_field_id_0_2,
  input  [7:0]   io_key_config_0_field_id_0_3,
  input  [7:0]   io_key_config_0_field_id_1_0,
  input  [7:0]   io_key_config_0_field_id_1_1,
  input  [7:0]   io_key_config_0_field_id_1_2,
  input  [7:0]   io_key_config_0_field_id_1_3,
  input  [7:0]   io_key_config_0_field_id_2_0,
  input  [7:0]   io_key_config_0_field_id_2_1,
  input  [7:0]   io_key_config_0_field_id_2_2,
  input  [7:0]   io_key_config_0_field_id_2_3,
  input  [7:0]   io_key_config_0_field_id_3_0,
  input  [7:0]   io_key_config_0_field_id_3_1,
  input  [7:0]   io_key_config_0_field_id_3_2,
  input  [7:0]   io_key_config_0_field_id_3_3,
  input  [7:0]   io_key_config_0_field_id_4_0,
  input  [7:0]   io_key_config_0_field_id_4_1,
  input  [7:0]   io_key_config_0_field_id_4_2,
  input  [7:0]   io_key_config_0_field_id_4_3,
  input  [7:0]   io_key_config_0_field_id_5_0,
  input  [7:0]   io_key_config_0_field_id_5_1,
  input  [7:0]   io_key_config_0_field_id_5_2,
  input  [7:0]   io_key_config_0_field_id_5_3,
  input  [1:0]   io_key_config_1_field_config_0,
  input  [1:0]   io_key_config_1_field_config_1,
  input  [1:0]   io_key_config_1_field_config_2,
  input  [1:0]   io_key_config_1_field_config_3,
  input  [1:0]   io_key_config_1_field_config_4,
  input  [1:0]   io_key_config_1_field_config_5,
  input          io_key_config_1_field_mask_0_0,
  input          io_key_config_1_field_mask_0_1,
  input          io_key_config_1_field_mask_0_2,
  input          io_key_config_1_field_mask_0_3,
  input          io_key_config_1_field_mask_1_0,
  input          io_key_config_1_field_mask_1_1,
  input          io_key_config_1_field_mask_1_2,
  input          io_key_config_1_field_mask_1_3,
  input          io_key_config_1_field_mask_2_0,
  input          io_key_config_1_field_mask_2_1,
  input          io_key_config_1_field_mask_2_2,
  input          io_key_config_1_field_mask_2_3,
  input          io_key_config_1_field_mask_3_0,
  input          io_key_config_1_field_mask_3_1,
  input          io_key_config_1_field_mask_3_2,
  input          io_key_config_1_field_mask_3_3,
  input          io_key_config_1_field_mask_4_0,
  input          io_key_config_1_field_mask_4_1,
  input          io_key_config_1_field_mask_4_2,
  input          io_key_config_1_field_mask_4_3,
  input          io_key_config_1_field_mask_5_0,
  input          io_key_config_1_field_mask_5_1,
  input          io_key_config_1_field_mask_5_2,
  input          io_key_config_1_field_mask_5_3,
  input  [7:0]   io_key_config_1_field_id_0_0,
  input  [7:0]   io_key_config_1_field_id_0_1,
  input  [7:0]   io_key_config_1_field_id_0_2,
  input  [7:0]   io_key_config_1_field_id_0_3,
  input  [7:0]   io_key_config_1_field_id_1_0,
  input  [7:0]   io_key_config_1_field_id_1_1,
  input  [7:0]   io_key_config_1_field_id_1_2,
  input  [7:0]   io_key_config_1_field_id_1_3,
  input  [7:0]   io_key_config_1_field_id_2_0,
  input  [7:0]   io_key_config_1_field_id_2_1,
  input  [7:0]   io_key_config_1_field_id_2_2,
  input  [7:0]   io_key_config_1_field_id_2_3,
  input  [7:0]   io_key_config_1_field_id_3_0,
  input  [7:0]   io_key_config_1_field_id_3_1,
  input  [7:0]   io_key_config_1_field_id_3_2,
  input  [7:0]   io_key_config_1_field_id_3_3,
  input  [7:0]   io_key_config_1_field_id_4_0,
  input  [7:0]   io_key_config_1_field_id_4_1,
  input  [7:0]   io_key_config_1_field_id_4_2,
  input  [7:0]   io_key_config_1_field_id_4_3,
  input  [7:0]   io_key_config_1_field_id_5_0,
  input  [7:0]   io_key_config_1_field_id_5_1,
  input  [7:0]   io_key_config_1_field_id_5_2,
  input  [7:0]   io_key_config_1_field_id_5_3,
  output [191:0] io_match_key
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] phv_data_0; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_1; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_2; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_3; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_4; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_5; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_6; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_7; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_8; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_9; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_10; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_11; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_12; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_13; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_14; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_15; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_16; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_17; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_18; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_19; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_20; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_21; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_22; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_23; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_24; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_25; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_26; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_27; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_28; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_29; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_30; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_31; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_32; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_33; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_34; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_35; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_36; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_37; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_38; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_39; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_40; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_41; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_42; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_43; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_44; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_45; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_46; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_47; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_48; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_49; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_50; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_51; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_52; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_53; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_54; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_55; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_56; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_57; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_58; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_59; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_60; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_61; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_62; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_63; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_64; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_65; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_66; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_67; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_68; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_69; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_70; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_71; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_72; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_73; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_74; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_75; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_76; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_77; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_78; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_79; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_80; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_81; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_82; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_83; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_84; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_85; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_86; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_87; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_88; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_89; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_90; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_91; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_92; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_93; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_94; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_95; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_96; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_97; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_98; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_99; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_100; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_101; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_102; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_103; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_104; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_105; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_106; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_107; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_108; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_109; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_110; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_111; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_112; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_113; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_114; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_115; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_116; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_117; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_118; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_119; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_120; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_121; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_122; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_123; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_124; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_125; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_126; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_127; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_128; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_129; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_130; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_131; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_132; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_133; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_134; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_135; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_136; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_137; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_138; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_139; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_140; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_141; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_142; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_143; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_144; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_145; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_146; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_147; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_148; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_149; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_150; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_151; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_152; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_153; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_154; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_155; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_156; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_157; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_158; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_159; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_160; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_161; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_162; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_163; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_164; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_165; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_166; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_167; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_168; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_169; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_170; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_171; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_172; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_173; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_174; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_175; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_176; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_177; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_178; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_179; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_180; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_181; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_182; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_183; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_184; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_185; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_186; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_187; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_188; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_189; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_190; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_191; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_192; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_193; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_194; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_195; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_196; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_197; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_198; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_199; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_200; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_201; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_202; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_203; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_204; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_205; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_206; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_207; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_208; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_209; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_210; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_211; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_212; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_213; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_214; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_215; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_216; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_217; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_218; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_219; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_220; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_221; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_222; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_223; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_224; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_225; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_226; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_227; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_228; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_229; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_230; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_231; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_232; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_233; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_234; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_235; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_236; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_237; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_238; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_239; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_240; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_241; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_242; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_243; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_244; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_245; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_246; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_247; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_248; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_249; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_250; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_251; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_252; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_253; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_254; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_255; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_256; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_257; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_258; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_259; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_260; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_261; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_262; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_263; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_264; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_265; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_266; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_267; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_268; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_269; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_270; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_271; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_272; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_273; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_274; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_275; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_276; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_277; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_278; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_279; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_280; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_281; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_282; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_283; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_284; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_285; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_286; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_287; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_288; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_289; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_290; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_291; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_292; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_293; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_294; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_295; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_296; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_297; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_298; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_299; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_300; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_301; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_302; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_303; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_304; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_305; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_306; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_307; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_308; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_309; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_310; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_311; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_312; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_313; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_314; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_315; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_316; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_317; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_318; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_319; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_320; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_321; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_322; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_323; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_324; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_325; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_326; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_327; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_328; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_329; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_330; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_331; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_332; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_333; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_334; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_335; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_336; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_337; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_338; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_339; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_340; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_341; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_342; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_343; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_344; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_345; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_346; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_347; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_348; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_349; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_350; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_351; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_352; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_353; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_354; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_355; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_356; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_357; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_358; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_359; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_360; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_361; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_362; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_363; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_364; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_365; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_366; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_367; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_368; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_369; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_370; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_371; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_372; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_373; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_374; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_375; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_376; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_377; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_378; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_379; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_380; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_381; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_382; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_383; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_384; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_385; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_386; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_387; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_388; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_389; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_390; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_391; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_392; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_393; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_394; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_395; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_396; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_397; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_398; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_399; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_400; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_401; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_402; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_403; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_404; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_405; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_406; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_407; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_408; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_409; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_410; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_411; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_412; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_413; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_414; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_415; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_416; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_417; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_418; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_419; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_420; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_421; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_422; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_423; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_424; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_425; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_426; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_427; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_428; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_429; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_430; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_431; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_432; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_433; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_434; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_435; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_436; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_437; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_438; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_439; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_440; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_441; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_442; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_443; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_444; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_445; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_446; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_447; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_448; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_449; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_450; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_451; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_452; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_453; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_454; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_455; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_456; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_457; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_458; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_459; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_460; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_461; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_462; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_463; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_464; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_465; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_466; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_467; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_468; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_469; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_470; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_471; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_472; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_473; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_474; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_475; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_476; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_477; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_478; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_479; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_480; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_481; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_482; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_483; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_484; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_485; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_486; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_487; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_488; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_489; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_490; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_491; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_492; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_493; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_494; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_495; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_496; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_497; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_498; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_499; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_500; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_501; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_502; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_503; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_504; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_505; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_506; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_507; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_508; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_509; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_510; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_511; // @[matcher_pisa.scala 110:22]
  reg [3:0] phv_next_processor_id; // @[matcher_pisa.scala 110:22]
  reg  phv_next_config_id; // @[matcher_pisa.scala 110:22]
  reg  phv_is_valid_processor; // @[matcher_pisa.scala 110:22]
  wire [1:0] _GEN_56 = phv_next_config_id ? io_key_config_1_field_config_0 : io_key_config_0_field_config_0; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire [1:0] _GEN_57 = phv_next_config_id ? io_key_config_1_field_config_1 : io_key_config_0_field_config_1; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire [1:0] _GEN_58 = phv_next_config_id ? io_key_config_1_field_config_2 : io_key_config_0_field_config_2; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire [1:0] _GEN_59 = phv_next_config_id ? io_key_config_1_field_config_3 : io_key_config_0_field_config_3; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire [1:0] _GEN_60 = phv_next_config_id ? io_key_config_1_field_config_4 : io_key_config_0_field_config_4; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire [1:0] _GEN_61 = phv_next_config_id ? io_key_config_1_field_config_5 : io_key_config_0_field_config_5; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire  _GEN_62 = phv_next_config_id ? io_key_config_1_field_mask_0_0 : io_key_config_0_field_mask_0_0; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire  _GEN_63 = phv_next_config_id ? io_key_config_1_field_mask_0_1 : io_key_config_0_field_mask_0_1; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire  _GEN_64 = phv_next_config_id ? io_key_config_1_field_mask_0_2 : io_key_config_0_field_mask_0_2; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire  _GEN_65 = phv_next_config_id ? io_key_config_1_field_mask_0_3 : io_key_config_0_field_mask_0_3; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire  _GEN_66 = phv_next_config_id ? io_key_config_1_field_mask_1_0 : io_key_config_0_field_mask_1_0; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire  _GEN_67 = phv_next_config_id ? io_key_config_1_field_mask_1_1 : io_key_config_0_field_mask_1_1; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire  _GEN_68 = phv_next_config_id ? io_key_config_1_field_mask_1_2 : io_key_config_0_field_mask_1_2; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire  _GEN_69 = phv_next_config_id ? io_key_config_1_field_mask_1_3 : io_key_config_0_field_mask_1_3; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire  _GEN_70 = phv_next_config_id ? io_key_config_1_field_mask_2_0 : io_key_config_0_field_mask_2_0; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire  _GEN_71 = phv_next_config_id ? io_key_config_1_field_mask_2_1 : io_key_config_0_field_mask_2_1; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire  _GEN_72 = phv_next_config_id ? io_key_config_1_field_mask_2_2 : io_key_config_0_field_mask_2_2; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire  _GEN_73 = phv_next_config_id ? io_key_config_1_field_mask_2_3 : io_key_config_0_field_mask_2_3; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire  _GEN_74 = phv_next_config_id ? io_key_config_1_field_mask_3_0 : io_key_config_0_field_mask_3_0; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire  _GEN_75 = phv_next_config_id ? io_key_config_1_field_mask_3_1 : io_key_config_0_field_mask_3_1; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire  _GEN_76 = phv_next_config_id ? io_key_config_1_field_mask_3_2 : io_key_config_0_field_mask_3_2; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire  _GEN_77 = phv_next_config_id ? io_key_config_1_field_mask_3_3 : io_key_config_0_field_mask_3_3; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire  _GEN_78 = phv_next_config_id ? io_key_config_1_field_mask_4_0 : io_key_config_0_field_mask_4_0; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire  _GEN_79 = phv_next_config_id ? io_key_config_1_field_mask_4_1 : io_key_config_0_field_mask_4_1; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire  _GEN_80 = phv_next_config_id ? io_key_config_1_field_mask_4_2 : io_key_config_0_field_mask_4_2; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire  _GEN_81 = phv_next_config_id ? io_key_config_1_field_mask_4_3 : io_key_config_0_field_mask_4_3; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire  _GEN_82 = phv_next_config_id ? io_key_config_1_field_mask_5_0 : io_key_config_0_field_mask_5_0; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire  _GEN_83 = phv_next_config_id ? io_key_config_1_field_mask_5_1 : io_key_config_0_field_mask_5_1; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire  _GEN_84 = phv_next_config_id ? io_key_config_1_field_mask_5_2 : io_key_config_0_field_mask_5_2; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire  _GEN_85 = phv_next_config_id ? io_key_config_1_field_mask_5_3 : io_key_config_0_field_mask_5_3; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire [7:0] _GEN_86 = phv_next_config_id ? io_key_config_1_field_id_0_0 : io_key_config_0_field_id_0_0; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire [7:0] _GEN_87 = phv_next_config_id ? io_key_config_1_field_id_0_1 : io_key_config_0_field_id_0_1; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire [7:0] _GEN_88 = phv_next_config_id ? io_key_config_1_field_id_0_2 : io_key_config_0_field_id_0_2; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire [7:0] _GEN_89 = phv_next_config_id ? io_key_config_1_field_id_0_3 : io_key_config_0_field_id_0_3; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire [7:0] _GEN_90 = phv_next_config_id ? io_key_config_1_field_id_1_0 : io_key_config_0_field_id_1_0; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire [7:0] _GEN_91 = phv_next_config_id ? io_key_config_1_field_id_1_1 : io_key_config_0_field_id_1_1; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire [7:0] _GEN_92 = phv_next_config_id ? io_key_config_1_field_id_1_2 : io_key_config_0_field_id_1_2; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire [7:0] _GEN_93 = phv_next_config_id ? io_key_config_1_field_id_1_3 : io_key_config_0_field_id_1_3; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire [7:0] _GEN_94 = phv_next_config_id ? io_key_config_1_field_id_2_0 : io_key_config_0_field_id_2_0; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire [7:0] _GEN_95 = phv_next_config_id ? io_key_config_1_field_id_2_1 : io_key_config_0_field_id_2_1; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire [7:0] _GEN_96 = phv_next_config_id ? io_key_config_1_field_id_2_2 : io_key_config_0_field_id_2_2; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire [7:0] _GEN_97 = phv_next_config_id ? io_key_config_1_field_id_2_3 : io_key_config_0_field_id_2_3; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire [7:0] _GEN_98 = phv_next_config_id ? io_key_config_1_field_id_3_0 : io_key_config_0_field_id_3_0; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire [7:0] _GEN_99 = phv_next_config_id ? io_key_config_1_field_id_3_1 : io_key_config_0_field_id_3_1; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire [7:0] _GEN_100 = phv_next_config_id ? io_key_config_1_field_id_3_2 : io_key_config_0_field_id_3_2; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire [7:0] _GEN_101 = phv_next_config_id ? io_key_config_1_field_id_3_3 : io_key_config_0_field_id_3_3; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire [7:0] _GEN_102 = phv_next_config_id ? io_key_config_1_field_id_4_0 : io_key_config_0_field_id_4_0; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire [7:0] _GEN_103 = phv_next_config_id ? io_key_config_1_field_id_4_1 : io_key_config_0_field_id_4_1; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire [7:0] _GEN_104 = phv_next_config_id ? io_key_config_1_field_id_4_2 : io_key_config_0_field_id_4_2; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire [7:0] _GEN_105 = phv_next_config_id ? io_key_config_1_field_id_4_3 : io_key_config_0_field_id_4_3; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire [7:0] _GEN_106 = phv_next_config_id ? io_key_config_1_field_id_5_0 : io_key_config_0_field_id_5_0; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire [7:0] _GEN_107 = phv_next_config_id ? io_key_config_1_field_id_5_1 : io_key_config_0_field_id_5_1; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire [7:0] _GEN_108 = phv_next_config_id ? io_key_config_1_field_id_5_2 : io_key_config_0_field_id_5_2; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire [7:0] _GEN_109 = phv_next_config_id ? io_key_config_1_field_id_5_3 : io_key_config_0_field_id_5_3; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire [7:0] _GEN_110 = 8'h0 == _GEN_86 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_111 = 8'h1 == _GEN_86 ? phv_data_1 : _GEN_110; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_112 = 8'h2 == _GEN_86 ? phv_data_2 : _GEN_111; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_113 = 8'h3 == _GEN_86 ? phv_data_3 : _GEN_112; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_114 = 8'h4 == _GEN_86 ? phv_data_4 : _GEN_113; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_115 = 8'h5 == _GEN_86 ? phv_data_5 : _GEN_114; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_116 = 8'h6 == _GEN_86 ? phv_data_6 : _GEN_115; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_117 = 8'h7 == _GEN_86 ? phv_data_7 : _GEN_116; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_118 = 8'h8 == _GEN_86 ? phv_data_8 : _GEN_117; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_119 = 8'h9 == _GEN_86 ? phv_data_9 : _GEN_118; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_120 = 8'ha == _GEN_86 ? phv_data_10 : _GEN_119; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_121 = 8'hb == _GEN_86 ? phv_data_11 : _GEN_120; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_122 = 8'hc == _GEN_86 ? phv_data_12 : _GEN_121; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_123 = 8'hd == _GEN_86 ? phv_data_13 : _GEN_122; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_124 = 8'he == _GEN_86 ? phv_data_14 : _GEN_123; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_125 = 8'hf == _GEN_86 ? phv_data_15 : _GEN_124; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_126 = 8'h10 == _GEN_86 ? phv_data_16 : _GEN_125; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_127 = 8'h11 == _GEN_86 ? phv_data_17 : _GEN_126; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_128 = 8'h12 == _GEN_86 ? phv_data_18 : _GEN_127; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_129 = 8'h13 == _GEN_86 ? phv_data_19 : _GEN_128; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_130 = 8'h14 == _GEN_86 ? phv_data_20 : _GEN_129; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_131 = 8'h15 == _GEN_86 ? phv_data_21 : _GEN_130; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_132 = 8'h16 == _GEN_86 ? phv_data_22 : _GEN_131; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_133 = 8'h17 == _GEN_86 ? phv_data_23 : _GEN_132; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_134 = 8'h18 == _GEN_86 ? phv_data_24 : _GEN_133; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_135 = 8'h19 == _GEN_86 ? phv_data_25 : _GEN_134; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_136 = 8'h1a == _GEN_86 ? phv_data_26 : _GEN_135; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_137 = 8'h1b == _GEN_86 ? phv_data_27 : _GEN_136; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_138 = 8'h1c == _GEN_86 ? phv_data_28 : _GEN_137; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_139 = 8'h1d == _GEN_86 ? phv_data_29 : _GEN_138; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_140 = 8'h1e == _GEN_86 ? phv_data_30 : _GEN_139; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_141 = 8'h1f == _GEN_86 ? phv_data_31 : _GEN_140; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_142 = 8'h20 == _GEN_86 ? phv_data_32 : _GEN_141; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_143 = 8'h21 == _GEN_86 ? phv_data_33 : _GEN_142; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_144 = 8'h22 == _GEN_86 ? phv_data_34 : _GEN_143; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_145 = 8'h23 == _GEN_86 ? phv_data_35 : _GEN_144; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_146 = 8'h24 == _GEN_86 ? phv_data_36 : _GEN_145; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_147 = 8'h25 == _GEN_86 ? phv_data_37 : _GEN_146; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_148 = 8'h26 == _GEN_86 ? phv_data_38 : _GEN_147; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_149 = 8'h27 == _GEN_86 ? phv_data_39 : _GEN_148; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_150 = 8'h28 == _GEN_86 ? phv_data_40 : _GEN_149; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_151 = 8'h29 == _GEN_86 ? phv_data_41 : _GEN_150; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_152 = 8'h2a == _GEN_86 ? phv_data_42 : _GEN_151; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_153 = 8'h2b == _GEN_86 ? phv_data_43 : _GEN_152; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_154 = 8'h2c == _GEN_86 ? phv_data_44 : _GEN_153; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_155 = 8'h2d == _GEN_86 ? phv_data_45 : _GEN_154; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_156 = 8'h2e == _GEN_86 ? phv_data_46 : _GEN_155; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_157 = 8'h2f == _GEN_86 ? phv_data_47 : _GEN_156; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_158 = 8'h30 == _GEN_86 ? phv_data_48 : _GEN_157; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_159 = 8'h31 == _GEN_86 ? phv_data_49 : _GEN_158; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_160 = 8'h32 == _GEN_86 ? phv_data_50 : _GEN_159; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_161 = 8'h33 == _GEN_86 ? phv_data_51 : _GEN_160; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_162 = 8'h34 == _GEN_86 ? phv_data_52 : _GEN_161; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_163 = 8'h35 == _GEN_86 ? phv_data_53 : _GEN_162; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_164 = 8'h36 == _GEN_86 ? phv_data_54 : _GEN_163; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_165 = 8'h37 == _GEN_86 ? phv_data_55 : _GEN_164; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_166 = 8'h38 == _GEN_86 ? phv_data_56 : _GEN_165; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_167 = 8'h39 == _GEN_86 ? phv_data_57 : _GEN_166; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_168 = 8'h3a == _GEN_86 ? phv_data_58 : _GEN_167; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_169 = 8'h3b == _GEN_86 ? phv_data_59 : _GEN_168; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_170 = 8'h3c == _GEN_86 ? phv_data_60 : _GEN_169; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_171 = 8'h3d == _GEN_86 ? phv_data_61 : _GEN_170; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_172 = 8'h3e == _GEN_86 ? phv_data_62 : _GEN_171; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_173 = 8'h3f == _GEN_86 ? phv_data_63 : _GEN_172; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] bytes__0 = _GEN_62 ? _GEN_173 : 8'h0; // @[matcher_pisa.scala 129:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_175 = 8'h0 == _GEN_87 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_176 = 8'h1 == _GEN_87 ? phv_data_1 : _GEN_175; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_177 = 8'h2 == _GEN_87 ? phv_data_2 : _GEN_176; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_178 = 8'h3 == _GEN_87 ? phv_data_3 : _GEN_177; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_179 = 8'h4 == _GEN_87 ? phv_data_4 : _GEN_178; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_180 = 8'h5 == _GEN_87 ? phv_data_5 : _GEN_179; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_181 = 8'h6 == _GEN_87 ? phv_data_6 : _GEN_180; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_182 = 8'h7 == _GEN_87 ? phv_data_7 : _GEN_181; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_183 = 8'h8 == _GEN_87 ? phv_data_8 : _GEN_182; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_184 = 8'h9 == _GEN_87 ? phv_data_9 : _GEN_183; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_185 = 8'ha == _GEN_87 ? phv_data_10 : _GEN_184; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_186 = 8'hb == _GEN_87 ? phv_data_11 : _GEN_185; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_187 = 8'hc == _GEN_87 ? phv_data_12 : _GEN_186; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_188 = 8'hd == _GEN_87 ? phv_data_13 : _GEN_187; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_189 = 8'he == _GEN_87 ? phv_data_14 : _GEN_188; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_190 = 8'hf == _GEN_87 ? phv_data_15 : _GEN_189; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_191 = 8'h10 == _GEN_87 ? phv_data_16 : _GEN_190; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_192 = 8'h11 == _GEN_87 ? phv_data_17 : _GEN_191; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_193 = 8'h12 == _GEN_87 ? phv_data_18 : _GEN_192; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_194 = 8'h13 == _GEN_87 ? phv_data_19 : _GEN_193; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_195 = 8'h14 == _GEN_87 ? phv_data_20 : _GEN_194; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_196 = 8'h15 == _GEN_87 ? phv_data_21 : _GEN_195; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_197 = 8'h16 == _GEN_87 ? phv_data_22 : _GEN_196; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_198 = 8'h17 == _GEN_87 ? phv_data_23 : _GEN_197; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_199 = 8'h18 == _GEN_87 ? phv_data_24 : _GEN_198; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_200 = 8'h19 == _GEN_87 ? phv_data_25 : _GEN_199; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_201 = 8'h1a == _GEN_87 ? phv_data_26 : _GEN_200; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_202 = 8'h1b == _GEN_87 ? phv_data_27 : _GEN_201; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_203 = 8'h1c == _GEN_87 ? phv_data_28 : _GEN_202; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_204 = 8'h1d == _GEN_87 ? phv_data_29 : _GEN_203; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_205 = 8'h1e == _GEN_87 ? phv_data_30 : _GEN_204; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_206 = 8'h1f == _GEN_87 ? phv_data_31 : _GEN_205; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_207 = 8'h20 == _GEN_87 ? phv_data_32 : _GEN_206; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_208 = 8'h21 == _GEN_87 ? phv_data_33 : _GEN_207; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_209 = 8'h22 == _GEN_87 ? phv_data_34 : _GEN_208; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_210 = 8'h23 == _GEN_87 ? phv_data_35 : _GEN_209; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_211 = 8'h24 == _GEN_87 ? phv_data_36 : _GEN_210; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_212 = 8'h25 == _GEN_87 ? phv_data_37 : _GEN_211; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_213 = 8'h26 == _GEN_87 ? phv_data_38 : _GEN_212; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_214 = 8'h27 == _GEN_87 ? phv_data_39 : _GEN_213; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_215 = 8'h28 == _GEN_87 ? phv_data_40 : _GEN_214; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_216 = 8'h29 == _GEN_87 ? phv_data_41 : _GEN_215; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_217 = 8'h2a == _GEN_87 ? phv_data_42 : _GEN_216; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_218 = 8'h2b == _GEN_87 ? phv_data_43 : _GEN_217; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_219 = 8'h2c == _GEN_87 ? phv_data_44 : _GEN_218; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_220 = 8'h2d == _GEN_87 ? phv_data_45 : _GEN_219; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_221 = 8'h2e == _GEN_87 ? phv_data_46 : _GEN_220; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_222 = 8'h2f == _GEN_87 ? phv_data_47 : _GEN_221; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_223 = 8'h30 == _GEN_87 ? phv_data_48 : _GEN_222; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_224 = 8'h31 == _GEN_87 ? phv_data_49 : _GEN_223; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_225 = 8'h32 == _GEN_87 ? phv_data_50 : _GEN_224; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_226 = 8'h33 == _GEN_87 ? phv_data_51 : _GEN_225; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_227 = 8'h34 == _GEN_87 ? phv_data_52 : _GEN_226; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_228 = 8'h35 == _GEN_87 ? phv_data_53 : _GEN_227; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_229 = 8'h36 == _GEN_87 ? phv_data_54 : _GEN_228; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_230 = 8'h37 == _GEN_87 ? phv_data_55 : _GEN_229; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_231 = 8'h38 == _GEN_87 ? phv_data_56 : _GEN_230; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_232 = 8'h39 == _GEN_87 ? phv_data_57 : _GEN_231; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_233 = 8'h3a == _GEN_87 ? phv_data_58 : _GEN_232; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_234 = 8'h3b == _GEN_87 ? phv_data_59 : _GEN_233; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_235 = 8'h3c == _GEN_87 ? phv_data_60 : _GEN_234; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_236 = 8'h3d == _GEN_87 ? phv_data_61 : _GEN_235; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_237 = 8'h3e == _GEN_87 ? phv_data_62 : _GEN_236; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_238 = 8'h3f == _GEN_87 ? phv_data_63 : _GEN_237; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] bytes__1 = _GEN_63 ? _GEN_238 : 8'h0; // @[matcher_pisa.scala 129:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_240 = 8'h0 == _GEN_88 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_241 = 8'h1 == _GEN_88 ? phv_data_1 : _GEN_240; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_242 = 8'h2 == _GEN_88 ? phv_data_2 : _GEN_241; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_243 = 8'h3 == _GEN_88 ? phv_data_3 : _GEN_242; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_244 = 8'h4 == _GEN_88 ? phv_data_4 : _GEN_243; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_245 = 8'h5 == _GEN_88 ? phv_data_5 : _GEN_244; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_246 = 8'h6 == _GEN_88 ? phv_data_6 : _GEN_245; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_247 = 8'h7 == _GEN_88 ? phv_data_7 : _GEN_246; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_248 = 8'h8 == _GEN_88 ? phv_data_8 : _GEN_247; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_249 = 8'h9 == _GEN_88 ? phv_data_9 : _GEN_248; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_250 = 8'ha == _GEN_88 ? phv_data_10 : _GEN_249; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_251 = 8'hb == _GEN_88 ? phv_data_11 : _GEN_250; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_252 = 8'hc == _GEN_88 ? phv_data_12 : _GEN_251; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_253 = 8'hd == _GEN_88 ? phv_data_13 : _GEN_252; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_254 = 8'he == _GEN_88 ? phv_data_14 : _GEN_253; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_255 = 8'hf == _GEN_88 ? phv_data_15 : _GEN_254; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_256 = 8'h10 == _GEN_88 ? phv_data_16 : _GEN_255; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_257 = 8'h11 == _GEN_88 ? phv_data_17 : _GEN_256; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_258 = 8'h12 == _GEN_88 ? phv_data_18 : _GEN_257; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_259 = 8'h13 == _GEN_88 ? phv_data_19 : _GEN_258; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_260 = 8'h14 == _GEN_88 ? phv_data_20 : _GEN_259; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_261 = 8'h15 == _GEN_88 ? phv_data_21 : _GEN_260; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_262 = 8'h16 == _GEN_88 ? phv_data_22 : _GEN_261; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_263 = 8'h17 == _GEN_88 ? phv_data_23 : _GEN_262; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_264 = 8'h18 == _GEN_88 ? phv_data_24 : _GEN_263; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_265 = 8'h19 == _GEN_88 ? phv_data_25 : _GEN_264; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_266 = 8'h1a == _GEN_88 ? phv_data_26 : _GEN_265; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_267 = 8'h1b == _GEN_88 ? phv_data_27 : _GEN_266; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_268 = 8'h1c == _GEN_88 ? phv_data_28 : _GEN_267; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_269 = 8'h1d == _GEN_88 ? phv_data_29 : _GEN_268; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_270 = 8'h1e == _GEN_88 ? phv_data_30 : _GEN_269; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_271 = 8'h1f == _GEN_88 ? phv_data_31 : _GEN_270; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_272 = 8'h20 == _GEN_88 ? phv_data_32 : _GEN_271; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_273 = 8'h21 == _GEN_88 ? phv_data_33 : _GEN_272; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_274 = 8'h22 == _GEN_88 ? phv_data_34 : _GEN_273; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_275 = 8'h23 == _GEN_88 ? phv_data_35 : _GEN_274; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_276 = 8'h24 == _GEN_88 ? phv_data_36 : _GEN_275; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_277 = 8'h25 == _GEN_88 ? phv_data_37 : _GEN_276; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_278 = 8'h26 == _GEN_88 ? phv_data_38 : _GEN_277; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_279 = 8'h27 == _GEN_88 ? phv_data_39 : _GEN_278; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_280 = 8'h28 == _GEN_88 ? phv_data_40 : _GEN_279; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_281 = 8'h29 == _GEN_88 ? phv_data_41 : _GEN_280; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_282 = 8'h2a == _GEN_88 ? phv_data_42 : _GEN_281; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_283 = 8'h2b == _GEN_88 ? phv_data_43 : _GEN_282; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_284 = 8'h2c == _GEN_88 ? phv_data_44 : _GEN_283; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_285 = 8'h2d == _GEN_88 ? phv_data_45 : _GEN_284; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_286 = 8'h2e == _GEN_88 ? phv_data_46 : _GEN_285; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_287 = 8'h2f == _GEN_88 ? phv_data_47 : _GEN_286; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_288 = 8'h30 == _GEN_88 ? phv_data_48 : _GEN_287; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_289 = 8'h31 == _GEN_88 ? phv_data_49 : _GEN_288; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_290 = 8'h32 == _GEN_88 ? phv_data_50 : _GEN_289; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_291 = 8'h33 == _GEN_88 ? phv_data_51 : _GEN_290; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_292 = 8'h34 == _GEN_88 ? phv_data_52 : _GEN_291; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_293 = 8'h35 == _GEN_88 ? phv_data_53 : _GEN_292; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_294 = 8'h36 == _GEN_88 ? phv_data_54 : _GEN_293; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_295 = 8'h37 == _GEN_88 ? phv_data_55 : _GEN_294; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_296 = 8'h38 == _GEN_88 ? phv_data_56 : _GEN_295; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_297 = 8'h39 == _GEN_88 ? phv_data_57 : _GEN_296; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_298 = 8'h3a == _GEN_88 ? phv_data_58 : _GEN_297; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_299 = 8'h3b == _GEN_88 ? phv_data_59 : _GEN_298; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_300 = 8'h3c == _GEN_88 ? phv_data_60 : _GEN_299; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_301 = 8'h3d == _GEN_88 ? phv_data_61 : _GEN_300; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_302 = 8'h3e == _GEN_88 ? phv_data_62 : _GEN_301; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_303 = 8'h3f == _GEN_88 ? phv_data_63 : _GEN_302; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] bytes__2 = _GEN_64 ? _GEN_303 : 8'h0; // @[matcher_pisa.scala 129:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_305 = 8'h0 == _GEN_89 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_306 = 8'h1 == _GEN_89 ? phv_data_1 : _GEN_305; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_307 = 8'h2 == _GEN_89 ? phv_data_2 : _GEN_306; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_308 = 8'h3 == _GEN_89 ? phv_data_3 : _GEN_307; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_309 = 8'h4 == _GEN_89 ? phv_data_4 : _GEN_308; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_310 = 8'h5 == _GEN_89 ? phv_data_5 : _GEN_309; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_311 = 8'h6 == _GEN_89 ? phv_data_6 : _GEN_310; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_312 = 8'h7 == _GEN_89 ? phv_data_7 : _GEN_311; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_313 = 8'h8 == _GEN_89 ? phv_data_8 : _GEN_312; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_314 = 8'h9 == _GEN_89 ? phv_data_9 : _GEN_313; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_315 = 8'ha == _GEN_89 ? phv_data_10 : _GEN_314; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_316 = 8'hb == _GEN_89 ? phv_data_11 : _GEN_315; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_317 = 8'hc == _GEN_89 ? phv_data_12 : _GEN_316; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_318 = 8'hd == _GEN_89 ? phv_data_13 : _GEN_317; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_319 = 8'he == _GEN_89 ? phv_data_14 : _GEN_318; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_320 = 8'hf == _GEN_89 ? phv_data_15 : _GEN_319; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_321 = 8'h10 == _GEN_89 ? phv_data_16 : _GEN_320; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_322 = 8'h11 == _GEN_89 ? phv_data_17 : _GEN_321; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_323 = 8'h12 == _GEN_89 ? phv_data_18 : _GEN_322; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_324 = 8'h13 == _GEN_89 ? phv_data_19 : _GEN_323; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_325 = 8'h14 == _GEN_89 ? phv_data_20 : _GEN_324; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_326 = 8'h15 == _GEN_89 ? phv_data_21 : _GEN_325; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_327 = 8'h16 == _GEN_89 ? phv_data_22 : _GEN_326; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_328 = 8'h17 == _GEN_89 ? phv_data_23 : _GEN_327; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_329 = 8'h18 == _GEN_89 ? phv_data_24 : _GEN_328; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_330 = 8'h19 == _GEN_89 ? phv_data_25 : _GEN_329; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_331 = 8'h1a == _GEN_89 ? phv_data_26 : _GEN_330; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_332 = 8'h1b == _GEN_89 ? phv_data_27 : _GEN_331; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_333 = 8'h1c == _GEN_89 ? phv_data_28 : _GEN_332; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_334 = 8'h1d == _GEN_89 ? phv_data_29 : _GEN_333; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_335 = 8'h1e == _GEN_89 ? phv_data_30 : _GEN_334; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_336 = 8'h1f == _GEN_89 ? phv_data_31 : _GEN_335; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_337 = 8'h20 == _GEN_89 ? phv_data_32 : _GEN_336; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_338 = 8'h21 == _GEN_89 ? phv_data_33 : _GEN_337; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_339 = 8'h22 == _GEN_89 ? phv_data_34 : _GEN_338; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_340 = 8'h23 == _GEN_89 ? phv_data_35 : _GEN_339; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_341 = 8'h24 == _GEN_89 ? phv_data_36 : _GEN_340; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_342 = 8'h25 == _GEN_89 ? phv_data_37 : _GEN_341; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_343 = 8'h26 == _GEN_89 ? phv_data_38 : _GEN_342; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_344 = 8'h27 == _GEN_89 ? phv_data_39 : _GEN_343; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_345 = 8'h28 == _GEN_89 ? phv_data_40 : _GEN_344; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_346 = 8'h29 == _GEN_89 ? phv_data_41 : _GEN_345; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_347 = 8'h2a == _GEN_89 ? phv_data_42 : _GEN_346; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_348 = 8'h2b == _GEN_89 ? phv_data_43 : _GEN_347; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_349 = 8'h2c == _GEN_89 ? phv_data_44 : _GEN_348; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_350 = 8'h2d == _GEN_89 ? phv_data_45 : _GEN_349; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_351 = 8'h2e == _GEN_89 ? phv_data_46 : _GEN_350; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_352 = 8'h2f == _GEN_89 ? phv_data_47 : _GEN_351; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_353 = 8'h30 == _GEN_89 ? phv_data_48 : _GEN_352; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_354 = 8'h31 == _GEN_89 ? phv_data_49 : _GEN_353; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_355 = 8'h32 == _GEN_89 ? phv_data_50 : _GEN_354; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_356 = 8'h33 == _GEN_89 ? phv_data_51 : _GEN_355; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_357 = 8'h34 == _GEN_89 ? phv_data_52 : _GEN_356; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_358 = 8'h35 == _GEN_89 ? phv_data_53 : _GEN_357; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_359 = 8'h36 == _GEN_89 ? phv_data_54 : _GEN_358; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_360 = 8'h37 == _GEN_89 ? phv_data_55 : _GEN_359; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_361 = 8'h38 == _GEN_89 ? phv_data_56 : _GEN_360; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_362 = 8'h39 == _GEN_89 ? phv_data_57 : _GEN_361; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_363 = 8'h3a == _GEN_89 ? phv_data_58 : _GEN_362; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_364 = 8'h3b == _GEN_89 ? phv_data_59 : _GEN_363; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_365 = 8'h3c == _GEN_89 ? phv_data_60 : _GEN_364; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_366 = 8'h3d == _GEN_89 ? phv_data_61 : _GEN_365; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_367 = 8'h3e == _GEN_89 ? phv_data_62 : _GEN_366; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_368 = 8'h3f == _GEN_89 ? phv_data_63 : _GEN_367; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] bytes__3 = _GEN_65 ? _GEN_368 : 8'h0; // @[matcher_pisa.scala 129:46 matcher_pisa.scala 128:34]
  wire [31:0] _groups_0_T = {bytes__0,bytes__1,bytes__2,bytes__3}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_370 = _GEN_56 == 2'h1 ? _groups_0_T : 32'h0; // @[matcher_pisa.scala 123:50 matcher_pisa.scala 137:31 matcher_pisa.scala 122:27]
  wire [15:0] _double_bytes_0_T = {phv_data_64,phv_data_65}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_371 = 8'h40 == _GEN_86 ? _double_bytes_0_T : 16'h0; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53 matcher_pisa.scala 144:41]
  wire [15:0] _double_bytes_0_T_1 = {phv_data_66,phv_data_67}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_372 = 8'h41 == _GEN_86 ? _double_bytes_0_T_1 : _GEN_371; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_2 = {phv_data_68,phv_data_69}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_373 = 8'h42 == _GEN_86 ? _double_bytes_0_T_2 : _GEN_372; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_3 = {phv_data_70,phv_data_71}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_374 = 8'h43 == _GEN_86 ? _double_bytes_0_T_3 : _GEN_373; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_4 = {phv_data_72,phv_data_73}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_375 = 8'h44 == _GEN_86 ? _double_bytes_0_T_4 : _GEN_374; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_5 = {phv_data_74,phv_data_75}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_376 = 8'h45 == _GEN_86 ? _double_bytes_0_T_5 : _GEN_375; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_6 = {phv_data_76,phv_data_77}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_377 = 8'h46 == _GEN_86 ? _double_bytes_0_T_6 : _GEN_376; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_7 = {phv_data_78,phv_data_79}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_378 = 8'h47 == _GEN_86 ? _double_bytes_0_T_7 : _GEN_377; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_8 = {phv_data_80,phv_data_81}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_379 = 8'h48 == _GEN_86 ? _double_bytes_0_T_8 : _GEN_378; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_9 = {phv_data_82,phv_data_83}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_380 = 8'h49 == _GEN_86 ? _double_bytes_0_T_9 : _GEN_379; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_10 = {phv_data_84,phv_data_85}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_381 = 8'h4a == _GEN_86 ? _double_bytes_0_T_10 : _GEN_380; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_11 = {phv_data_86,phv_data_87}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_382 = 8'h4b == _GEN_86 ? _double_bytes_0_T_11 : _GEN_381; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_12 = {phv_data_88,phv_data_89}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_383 = 8'h4c == _GEN_86 ? _double_bytes_0_T_12 : _GEN_382; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_13 = {phv_data_90,phv_data_91}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_384 = 8'h4d == _GEN_86 ? _double_bytes_0_T_13 : _GEN_383; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_14 = {phv_data_92,phv_data_93}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_385 = 8'h4e == _GEN_86 ? _double_bytes_0_T_14 : _GEN_384; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_15 = {phv_data_94,phv_data_95}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_386 = 8'h4f == _GEN_86 ? _double_bytes_0_T_15 : _GEN_385; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_16 = {phv_data_96,phv_data_97}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_387 = 8'h50 == _GEN_86 ? _double_bytes_0_T_16 : _GEN_386; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_17 = {phv_data_98,phv_data_99}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_388 = 8'h51 == _GEN_86 ? _double_bytes_0_T_17 : _GEN_387; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_18 = {phv_data_100,phv_data_101}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_389 = 8'h52 == _GEN_86 ? _double_bytes_0_T_18 : _GEN_388; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_19 = {phv_data_102,phv_data_103}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_390 = 8'h53 == _GEN_86 ? _double_bytes_0_T_19 : _GEN_389; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_20 = {phv_data_104,phv_data_105}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_391 = 8'h54 == _GEN_86 ? _double_bytes_0_T_20 : _GEN_390; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_21 = {phv_data_106,phv_data_107}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_392 = 8'h55 == _GEN_86 ? _double_bytes_0_T_21 : _GEN_391; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_22 = {phv_data_108,phv_data_109}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_393 = 8'h56 == _GEN_86 ? _double_bytes_0_T_22 : _GEN_392; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_23 = {phv_data_110,phv_data_111}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_394 = 8'h57 == _GEN_86 ? _double_bytes_0_T_23 : _GEN_393; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_24 = {phv_data_112,phv_data_113}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_395 = 8'h58 == _GEN_86 ? _double_bytes_0_T_24 : _GEN_394; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_25 = {phv_data_114,phv_data_115}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_396 = 8'h59 == _GEN_86 ? _double_bytes_0_T_25 : _GEN_395; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_26 = {phv_data_116,phv_data_117}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_397 = 8'h5a == _GEN_86 ? _double_bytes_0_T_26 : _GEN_396; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_27 = {phv_data_118,phv_data_119}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_398 = 8'h5b == _GEN_86 ? _double_bytes_0_T_27 : _GEN_397; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_28 = {phv_data_120,phv_data_121}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_399 = 8'h5c == _GEN_86 ? _double_bytes_0_T_28 : _GEN_398; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_29 = {phv_data_122,phv_data_123}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_400 = 8'h5d == _GEN_86 ? _double_bytes_0_T_29 : _GEN_399; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_30 = {phv_data_124,phv_data_125}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_401 = 8'h5e == _GEN_86 ? _double_bytes_0_T_30 : _GEN_400; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_31 = {phv_data_126,phv_data_127}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_402 = 8'h5f == _GEN_86 ? _double_bytes_0_T_31 : _GEN_401; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_32 = {phv_data_128,phv_data_129}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_403 = 8'h60 == _GEN_86 ? _double_bytes_0_T_32 : _GEN_402; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_33 = {phv_data_130,phv_data_131}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_404 = 8'h61 == _GEN_86 ? _double_bytes_0_T_33 : _GEN_403; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_34 = {phv_data_132,phv_data_133}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_405 = 8'h62 == _GEN_86 ? _double_bytes_0_T_34 : _GEN_404; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_35 = {phv_data_134,phv_data_135}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_406 = 8'h63 == _GEN_86 ? _double_bytes_0_T_35 : _GEN_405; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_36 = {phv_data_136,phv_data_137}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_407 = 8'h64 == _GEN_86 ? _double_bytes_0_T_36 : _GEN_406; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_37 = {phv_data_138,phv_data_139}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_408 = 8'h65 == _GEN_86 ? _double_bytes_0_T_37 : _GEN_407; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_38 = {phv_data_140,phv_data_141}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_409 = 8'h66 == _GEN_86 ? _double_bytes_0_T_38 : _GEN_408; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_39 = {phv_data_142,phv_data_143}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_410 = 8'h67 == _GEN_86 ? _double_bytes_0_T_39 : _GEN_409; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_40 = {phv_data_144,phv_data_145}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_411 = 8'h68 == _GEN_86 ? _double_bytes_0_T_40 : _GEN_410; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_41 = {phv_data_146,phv_data_147}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_412 = 8'h69 == _GEN_86 ? _double_bytes_0_T_41 : _GEN_411; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_42 = {phv_data_148,phv_data_149}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_413 = 8'h6a == _GEN_86 ? _double_bytes_0_T_42 : _GEN_412; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_43 = {phv_data_150,phv_data_151}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_414 = 8'h6b == _GEN_86 ? _double_bytes_0_T_43 : _GEN_413; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_44 = {phv_data_152,phv_data_153}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_415 = 8'h6c == _GEN_86 ? _double_bytes_0_T_44 : _GEN_414; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_45 = {phv_data_154,phv_data_155}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_416 = 8'h6d == _GEN_86 ? _double_bytes_0_T_45 : _GEN_415; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_46 = {phv_data_156,phv_data_157}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_417 = 8'h6e == _GEN_86 ? _double_bytes_0_T_46 : _GEN_416; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_47 = {phv_data_158,phv_data_159}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_418 = 8'h6f == _GEN_86 ? _double_bytes_0_T_47 : _GEN_417; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_48 = {phv_data_160,phv_data_161}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_419 = 8'h70 == _GEN_86 ? _double_bytes_0_T_48 : _GEN_418; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_49 = {phv_data_162,phv_data_163}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_420 = 8'h71 == _GEN_86 ? _double_bytes_0_T_49 : _GEN_419; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_50 = {phv_data_164,phv_data_165}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_421 = 8'h72 == _GEN_86 ? _double_bytes_0_T_50 : _GEN_420; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_51 = {phv_data_166,phv_data_167}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_422 = 8'h73 == _GEN_86 ? _double_bytes_0_T_51 : _GEN_421; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_52 = {phv_data_168,phv_data_169}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_423 = 8'h74 == _GEN_86 ? _double_bytes_0_T_52 : _GEN_422; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_53 = {phv_data_170,phv_data_171}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_424 = 8'h75 == _GEN_86 ? _double_bytes_0_T_53 : _GEN_423; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_54 = {phv_data_172,phv_data_173}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_425 = 8'h76 == _GEN_86 ? _double_bytes_0_T_54 : _GEN_424; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_55 = {phv_data_174,phv_data_175}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_426 = 8'h77 == _GEN_86 ? _double_bytes_0_T_55 : _GEN_425; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_56 = {phv_data_176,phv_data_177}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_427 = 8'h78 == _GEN_86 ? _double_bytes_0_T_56 : _GEN_426; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_57 = {phv_data_178,phv_data_179}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_428 = 8'h79 == _GEN_86 ? _double_bytes_0_T_57 : _GEN_427; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_58 = {phv_data_180,phv_data_181}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_429 = 8'h7a == _GEN_86 ? _double_bytes_0_T_58 : _GEN_428; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_59 = {phv_data_182,phv_data_183}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_430 = 8'h7b == _GEN_86 ? _double_bytes_0_T_59 : _GEN_429; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_60 = {phv_data_184,phv_data_185}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_431 = 8'h7c == _GEN_86 ? _double_bytes_0_T_60 : _GEN_430; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_61 = {phv_data_186,phv_data_187}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_432 = 8'h7d == _GEN_86 ? _double_bytes_0_T_61 : _GEN_431; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_62 = {phv_data_188,phv_data_189}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_433 = 8'h7e == _GEN_86 ? _double_bytes_0_T_62 : _GEN_432; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_63 = {phv_data_190,phv_data_191}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_434 = 8'h7f == _GEN_86 ? _double_bytes_0_T_63 : _GEN_433; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_64 = {phv_data_192,phv_data_193}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_435 = 8'h80 == _GEN_86 ? _double_bytes_0_T_64 : _GEN_434; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_65 = {phv_data_194,phv_data_195}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_436 = 8'h81 == _GEN_86 ? _double_bytes_0_T_65 : _GEN_435; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_66 = {phv_data_196,phv_data_197}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_437 = 8'h82 == _GEN_86 ? _double_bytes_0_T_66 : _GEN_436; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_67 = {phv_data_198,phv_data_199}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_438 = 8'h83 == _GEN_86 ? _double_bytes_0_T_67 : _GEN_437; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_68 = {phv_data_200,phv_data_201}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_439 = 8'h84 == _GEN_86 ? _double_bytes_0_T_68 : _GEN_438; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_69 = {phv_data_202,phv_data_203}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_440 = 8'h85 == _GEN_86 ? _double_bytes_0_T_69 : _GEN_439; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_70 = {phv_data_204,phv_data_205}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_441 = 8'h86 == _GEN_86 ? _double_bytes_0_T_70 : _GEN_440; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_71 = {phv_data_206,phv_data_207}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_442 = 8'h87 == _GEN_86 ? _double_bytes_0_T_71 : _GEN_441; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_72 = {phv_data_208,phv_data_209}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_443 = 8'h88 == _GEN_86 ? _double_bytes_0_T_72 : _GEN_442; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_73 = {phv_data_210,phv_data_211}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_444 = 8'h89 == _GEN_86 ? _double_bytes_0_T_73 : _GEN_443; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_74 = {phv_data_212,phv_data_213}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_445 = 8'h8a == _GEN_86 ? _double_bytes_0_T_74 : _GEN_444; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_75 = {phv_data_214,phv_data_215}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_446 = 8'h8b == _GEN_86 ? _double_bytes_0_T_75 : _GEN_445; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_76 = {phv_data_216,phv_data_217}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_447 = 8'h8c == _GEN_86 ? _double_bytes_0_T_76 : _GEN_446; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_77 = {phv_data_218,phv_data_219}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_448 = 8'h8d == _GEN_86 ? _double_bytes_0_T_77 : _GEN_447; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_78 = {phv_data_220,phv_data_221}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_449 = 8'h8e == _GEN_86 ? _double_bytes_0_T_78 : _GEN_448; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_79 = {phv_data_222,phv_data_223}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_450 = 8'h8f == _GEN_86 ? _double_bytes_0_T_79 : _GEN_449; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_80 = {phv_data_224,phv_data_225}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_451 = 8'h90 == _GEN_86 ? _double_bytes_0_T_80 : _GEN_450; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_81 = {phv_data_226,phv_data_227}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_452 = 8'h91 == _GEN_86 ? _double_bytes_0_T_81 : _GEN_451; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_82 = {phv_data_228,phv_data_229}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_453 = 8'h92 == _GEN_86 ? _double_bytes_0_T_82 : _GEN_452; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_83 = {phv_data_230,phv_data_231}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_454 = 8'h93 == _GEN_86 ? _double_bytes_0_T_83 : _GEN_453; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_84 = {phv_data_232,phv_data_233}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_455 = 8'h94 == _GEN_86 ? _double_bytes_0_T_84 : _GEN_454; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_85 = {phv_data_234,phv_data_235}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_456 = 8'h95 == _GEN_86 ? _double_bytes_0_T_85 : _GEN_455; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_86 = {phv_data_236,phv_data_237}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_457 = 8'h96 == _GEN_86 ? _double_bytes_0_T_86 : _GEN_456; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_87 = {phv_data_238,phv_data_239}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_458 = 8'h97 == _GEN_86 ? _double_bytes_0_T_87 : _GEN_457; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_88 = {phv_data_240,phv_data_241}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_459 = 8'h98 == _GEN_86 ? _double_bytes_0_T_88 : _GEN_458; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_89 = {phv_data_242,phv_data_243}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_460 = 8'h99 == _GEN_86 ? _double_bytes_0_T_89 : _GEN_459; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_90 = {phv_data_244,phv_data_245}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_461 = 8'h9a == _GEN_86 ? _double_bytes_0_T_90 : _GEN_460; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_91 = {phv_data_246,phv_data_247}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_462 = 8'h9b == _GEN_86 ? _double_bytes_0_T_91 : _GEN_461; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_92 = {phv_data_248,phv_data_249}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_463 = 8'h9c == _GEN_86 ? _double_bytes_0_T_92 : _GEN_462; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_93 = {phv_data_250,phv_data_251}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_464 = 8'h9d == _GEN_86 ? _double_bytes_0_T_93 : _GEN_463; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_94 = {phv_data_252,phv_data_253}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_465 = 8'h9e == _GEN_86 ? _double_bytes_0_T_94 : _GEN_464; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_95 = {phv_data_254,phv_data_255}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_466 = 8'h9f == _GEN_86 ? _double_bytes_0_T_95 : _GEN_465; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] double_bytes__0 = _GEN_62 ? _GEN_466 : 16'h0; // @[matcher_pisa.scala 145:46 matcher_pisa.scala 144:41]
  wire [15:0] _GEN_468 = 8'h40 == _GEN_87 ? _double_bytes_0_T : 16'h0; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53 matcher_pisa.scala 144:41]
  wire [15:0] _GEN_469 = 8'h41 == _GEN_87 ? _double_bytes_0_T_1 : _GEN_468; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_470 = 8'h42 == _GEN_87 ? _double_bytes_0_T_2 : _GEN_469; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_471 = 8'h43 == _GEN_87 ? _double_bytes_0_T_3 : _GEN_470; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_472 = 8'h44 == _GEN_87 ? _double_bytes_0_T_4 : _GEN_471; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_473 = 8'h45 == _GEN_87 ? _double_bytes_0_T_5 : _GEN_472; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_474 = 8'h46 == _GEN_87 ? _double_bytes_0_T_6 : _GEN_473; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_475 = 8'h47 == _GEN_87 ? _double_bytes_0_T_7 : _GEN_474; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_476 = 8'h48 == _GEN_87 ? _double_bytes_0_T_8 : _GEN_475; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_477 = 8'h49 == _GEN_87 ? _double_bytes_0_T_9 : _GEN_476; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_478 = 8'h4a == _GEN_87 ? _double_bytes_0_T_10 : _GEN_477; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_479 = 8'h4b == _GEN_87 ? _double_bytes_0_T_11 : _GEN_478; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_480 = 8'h4c == _GEN_87 ? _double_bytes_0_T_12 : _GEN_479; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_481 = 8'h4d == _GEN_87 ? _double_bytes_0_T_13 : _GEN_480; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_482 = 8'h4e == _GEN_87 ? _double_bytes_0_T_14 : _GEN_481; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_483 = 8'h4f == _GEN_87 ? _double_bytes_0_T_15 : _GEN_482; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_484 = 8'h50 == _GEN_87 ? _double_bytes_0_T_16 : _GEN_483; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_485 = 8'h51 == _GEN_87 ? _double_bytes_0_T_17 : _GEN_484; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_486 = 8'h52 == _GEN_87 ? _double_bytes_0_T_18 : _GEN_485; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_487 = 8'h53 == _GEN_87 ? _double_bytes_0_T_19 : _GEN_486; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_488 = 8'h54 == _GEN_87 ? _double_bytes_0_T_20 : _GEN_487; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_489 = 8'h55 == _GEN_87 ? _double_bytes_0_T_21 : _GEN_488; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_490 = 8'h56 == _GEN_87 ? _double_bytes_0_T_22 : _GEN_489; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_491 = 8'h57 == _GEN_87 ? _double_bytes_0_T_23 : _GEN_490; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_492 = 8'h58 == _GEN_87 ? _double_bytes_0_T_24 : _GEN_491; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_493 = 8'h59 == _GEN_87 ? _double_bytes_0_T_25 : _GEN_492; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_494 = 8'h5a == _GEN_87 ? _double_bytes_0_T_26 : _GEN_493; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_495 = 8'h5b == _GEN_87 ? _double_bytes_0_T_27 : _GEN_494; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_496 = 8'h5c == _GEN_87 ? _double_bytes_0_T_28 : _GEN_495; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_497 = 8'h5d == _GEN_87 ? _double_bytes_0_T_29 : _GEN_496; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_498 = 8'h5e == _GEN_87 ? _double_bytes_0_T_30 : _GEN_497; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_499 = 8'h5f == _GEN_87 ? _double_bytes_0_T_31 : _GEN_498; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_500 = 8'h60 == _GEN_87 ? _double_bytes_0_T_32 : _GEN_499; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_501 = 8'h61 == _GEN_87 ? _double_bytes_0_T_33 : _GEN_500; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_502 = 8'h62 == _GEN_87 ? _double_bytes_0_T_34 : _GEN_501; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_503 = 8'h63 == _GEN_87 ? _double_bytes_0_T_35 : _GEN_502; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_504 = 8'h64 == _GEN_87 ? _double_bytes_0_T_36 : _GEN_503; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_505 = 8'h65 == _GEN_87 ? _double_bytes_0_T_37 : _GEN_504; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_506 = 8'h66 == _GEN_87 ? _double_bytes_0_T_38 : _GEN_505; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_507 = 8'h67 == _GEN_87 ? _double_bytes_0_T_39 : _GEN_506; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_508 = 8'h68 == _GEN_87 ? _double_bytes_0_T_40 : _GEN_507; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_509 = 8'h69 == _GEN_87 ? _double_bytes_0_T_41 : _GEN_508; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_510 = 8'h6a == _GEN_87 ? _double_bytes_0_T_42 : _GEN_509; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_511 = 8'h6b == _GEN_87 ? _double_bytes_0_T_43 : _GEN_510; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_512 = 8'h6c == _GEN_87 ? _double_bytes_0_T_44 : _GEN_511; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_513 = 8'h6d == _GEN_87 ? _double_bytes_0_T_45 : _GEN_512; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_514 = 8'h6e == _GEN_87 ? _double_bytes_0_T_46 : _GEN_513; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_515 = 8'h6f == _GEN_87 ? _double_bytes_0_T_47 : _GEN_514; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_516 = 8'h70 == _GEN_87 ? _double_bytes_0_T_48 : _GEN_515; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_517 = 8'h71 == _GEN_87 ? _double_bytes_0_T_49 : _GEN_516; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_518 = 8'h72 == _GEN_87 ? _double_bytes_0_T_50 : _GEN_517; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_519 = 8'h73 == _GEN_87 ? _double_bytes_0_T_51 : _GEN_518; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_520 = 8'h74 == _GEN_87 ? _double_bytes_0_T_52 : _GEN_519; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_521 = 8'h75 == _GEN_87 ? _double_bytes_0_T_53 : _GEN_520; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_522 = 8'h76 == _GEN_87 ? _double_bytes_0_T_54 : _GEN_521; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_523 = 8'h77 == _GEN_87 ? _double_bytes_0_T_55 : _GEN_522; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_524 = 8'h78 == _GEN_87 ? _double_bytes_0_T_56 : _GEN_523; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_525 = 8'h79 == _GEN_87 ? _double_bytes_0_T_57 : _GEN_524; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_526 = 8'h7a == _GEN_87 ? _double_bytes_0_T_58 : _GEN_525; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_527 = 8'h7b == _GEN_87 ? _double_bytes_0_T_59 : _GEN_526; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_528 = 8'h7c == _GEN_87 ? _double_bytes_0_T_60 : _GEN_527; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_529 = 8'h7d == _GEN_87 ? _double_bytes_0_T_61 : _GEN_528; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_530 = 8'h7e == _GEN_87 ? _double_bytes_0_T_62 : _GEN_529; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_531 = 8'h7f == _GEN_87 ? _double_bytes_0_T_63 : _GEN_530; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_532 = 8'h80 == _GEN_87 ? _double_bytes_0_T_64 : _GEN_531; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_533 = 8'h81 == _GEN_87 ? _double_bytes_0_T_65 : _GEN_532; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_534 = 8'h82 == _GEN_87 ? _double_bytes_0_T_66 : _GEN_533; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_535 = 8'h83 == _GEN_87 ? _double_bytes_0_T_67 : _GEN_534; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_536 = 8'h84 == _GEN_87 ? _double_bytes_0_T_68 : _GEN_535; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_537 = 8'h85 == _GEN_87 ? _double_bytes_0_T_69 : _GEN_536; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_538 = 8'h86 == _GEN_87 ? _double_bytes_0_T_70 : _GEN_537; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_539 = 8'h87 == _GEN_87 ? _double_bytes_0_T_71 : _GEN_538; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_540 = 8'h88 == _GEN_87 ? _double_bytes_0_T_72 : _GEN_539; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_541 = 8'h89 == _GEN_87 ? _double_bytes_0_T_73 : _GEN_540; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_542 = 8'h8a == _GEN_87 ? _double_bytes_0_T_74 : _GEN_541; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_543 = 8'h8b == _GEN_87 ? _double_bytes_0_T_75 : _GEN_542; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_544 = 8'h8c == _GEN_87 ? _double_bytes_0_T_76 : _GEN_543; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_545 = 8'h8d == _GEN_87 ? _double_bytes_0_T_77 : _GEN_544; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_546 = 8'h8e == _GEN_87 ? _double_bytes_0_T_78 : _GEN_545; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_547 = 8'h8f == _GEN_87 ? _double_bytes_0_T_79 : _GEN_546; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_548 = 8'h90 == _GEN_87 ? _double_bytes_0_T_80 : _GEN_547; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_549 = 8'h91 == _GEN_87 ? _double_bytes_0_T_81 : _GEN_548; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_550 = 8'h92 == _GEN_87 ? _double_bytes_0_T_82 : _GEN_549; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_551 = 8'h93 == _GEN_87 ? _double_bytes_0_T_83 : _GEN_550; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_552 = 8'h94 == _GEN_87 ? _double_bytes_0_T_84 : _GEN_551; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_553 = 8'h95 == _GEN_87 ? _double_bytes_0_T_85 : _GEN_552; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_554 = 8'h96 == _GEN_87 ? _double_bytes_0_T_86 : _GEN_553; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_555 = 8'h97 == _GEN_87 ? _double_bytes_0_T_87 : _GEN_554; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_556 = 8'h98 == _GEN_87 ? _double_bytes_0_T_88 : _GEN_555; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_557 = 8'h99 == _GEN_87 ? _double_bytes_0_T_89 : _GEN_556; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_558 = 8'h9a == _GEN_87 ? _double_bytes_0_T_90 : _GEN_557; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_559 = 8'h9b == _GEN_87 ? _double_bytes_0_T_91 : _GEN_558; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_560 = 8'h9c == _GEN_87 ? _double_bytes_0_T_92 : _GEN_559; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_561 = 8'h9d == _GEN_87 ? _double_bytes_0_T_93 : _GEN_560; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_562 = 8'h9e == _GEN_87 ? _double_bytes_0_T_94 : _GEN_561; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_563 = 8'h9f == _GEN_87 ? _double_bytes_0_T_95 : _GEN_562; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] double_bytes__1 = _GEN_63 ? _GEN_563 : 16'h0; // @[matcher_pisa.scala 145:46 matcher_pisa.scala 144:41]
  wire [31:0] _groups_0_T_1 = {double_bytes__0,double_bytes__1}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_565 = _GEN_56 == 2'h2 ? _groups_0_T_1 : _GEN_370; // @[matcher_pisa.scala 139:50 matcher_pisa.scala 153:31]
  wire [31:0] _groups_0_T_2 = {phv_data_256,phv_data_257,phv_data_258,phv_data_259}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_566 = 8'ha0 == _GEN_86 ? _groups_0_T_2 : 32'h0; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39 matcher_pisa.scala 158:31]
  wire [31:0] _groups_0_T_3 = {phv_data_260,phv_data_261,phv_data_262,phv_data_263}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_567 = 8'ha1 == _GEN_86 ? _groups_0_T_3 : _GEN_566; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_4 = {phv_data_264,phv_data_265,phv_data_266,phv_data_267}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_568 = 8'ha2 == _GEN_86 ? _groups_0_T_4 : _GEN_567; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_5 = {phv_data_268,phv_data_269,phv_data_270,phv_data_271}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_569 = 8'ha3 == _GEN_86 ? _groups_0_T_5 : _GEN_568; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_6 = {phv_data_272,phv_data_273,phv_data_274,phv_data_275}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_570 = 8'ha4 == _GEN_86 ? _groups_0_T_6 : _GEN_569; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_7 = {phv_data_276,phv_data_277,phv_data_278,phv_data_279}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_571 = 8'ha5 == _GEN_86 ? _groups_0_T_7 : _GEN_570; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_8 = {phv_data_280,phv_data_281,phv_data_282,phv_data_283}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_572 = 8'ha6 == _GEN_86 ? _groups_0_T_8 : _GEN_571; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_9 = {phv_data_284,phv_data_285,phv_data_286,phv_data_287}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_573 = 8'ha7 == _GEN_86 ? _groups_0_T_9 : _GEN_572; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_10 = {phv_data_288,phv_data_289,phv_data_290,phv_data_291}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_574 = 8'ha8 == _GEN_86 ? _groups_0_T_10 : _GEN_573; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_11 = {phv_data_292,phv_data_293,phv_data_294,phv_data_295}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_575 = 8'ha9 == _GEN_86 ? _groups_0_T_11 : _GEN_574; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_12 = {phv_data_296,phv_data_297,phv_data_298,phv_data_299}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_576 = 8'haa == _GEN_86 ? _groups_0_T_12 : _GEN_575; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_13 = {phv_data_300,phv_data_301,phv_data_302,phv_data_303}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_577 = 8'hab == _GEN_86 ? _groups_0_T_13 : _GEN_576; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_14 = {phv_data_304,phv_data_305,phv_data_306,phv_data_307}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_578 = 8'hac == _GEN_86 ? _groups_0_T_14 : _GEN_577; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_15 = {phv_data_308,phv_data_309,phv_data_310,phv_data_311}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_579 = 8'had == _GEN_86 ? _groups_0_T_15 : _GEN_578; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_16 = {phv_data_312,phv_data_313,phv_data_314,phv_data_315}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_580 = 8'hae == _GEN_86 ? _groups_0_T_16 : _GEN_579; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_17 = {phv_data_316,phv_data_317,phv_data_318,phv_data_319}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_581 = 8'haf == _GEN_86 ? _groups_0_T_17 : _GEN_580; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_18 = {phv_data_320,phv_data_321,phv_data_322,phv_data_323}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_582 = 8'hb0 == _GEN_86 ? _groups_0_T_18 : _GEN_581; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_19 = {phv_data_324,phv_data_325,phv_data_326,phv_data_327}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_583 = 8'hb1 == _GEN_86 ? _groups_0_T_19 : _GEN_582; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_20 = {phv_data_328,phv_data_329,phv_data_330,phv_data_331}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_584 = 8'hb2 == _GEN_86 ? _groups_0_T_20 : _GEN_583; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_21 = {phv_data_332,phv_data_333,phv_data_334,phv_data_335}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_585 = 8'hb3 == _GEN_86 ? _groups_0_T_21 : _GEN_584; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_22 = {phv_data_336,phv_data_337,phv_data_338,phv_data_339}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_586 = 8'hb4 == _GEN_86 ? _groups_0_T_22 : _GEN_585; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_23 = {phv_data_340,phv_data_341,phv_data_342,phv_data_343}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_587 = 8'hb5 == _GEN_86 ? _groups_0_T_23 : _GEN_586; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_24 = {phv_data_344,phv_data_345,phv_data_346,phv_data_347}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_588 = 8'hb6 == _GEN_86 ? _groups_0_T_24 : _GEN_587; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_25 = {phv_data_348,phv_data_349,phv_data_350,phv_data_351}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_589 = 8'hb7 == _GEN_86 ? _groups_0_T_25 : _GEN_588; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_26 = {phv_data_352,phv_data_353,phv_data_354,phv_data_355}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_590 = 8'hb8 == _GEN_86 ? _groups_0_T_26 : _GEN_589; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_27 = {phv_data_356,phv_data_357,phv_data_358,phv_data_359}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_591 = 8'hb9 == _GEN_86 ? _groups_0_T_27 : _GEN_590; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_28 = {phv_data_360,phv_data_361,phv_data_362,phv_data_363}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_592 = 8'hba == _GEN_86 ? _groups_0_T_28 : _GEN_591; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_29 = {phv_data_364,phv_data_365,phv_data_366,phv_data_367}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_593 = 8'hbb == _GEN_86 ? _groups_0_T_29 : _GEN_592; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_30 = {phv_data_368,phv_data_369,phv_data_370,phv_data_371}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_594 = 8'hbc == _GEN_86 ? _groups_0_T_30 : _GEN_593; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_31 = {phv_data_372,phv_data_373,phv_data_374,phv_data_375}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_595 = 8'hbd == _GEN_86 ? _groups_0_T_31 : _GEN_594; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_32 = {phv_data_376,phv_data_377,phv_data_378,phv_data_379}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_596 = 8'hbe == _GEN_86 ? _groups_0_T_32 : _GEN_595; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_33 = {phv_data_380,phv_data_381,phv_data_382,phv_data_383}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_597 = 8'hbf == _GEN_86 ? _groups_0_T_33 : _GEN_596; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_34 = {phv_data_384,phv_data_385,phv_data_386,phv_data_387}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_598 = 8'hc0 == _GEN_86 ? _groups_0_T_34 : _GEN_597; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_35 = {phv_data_388,phv_data_389,phv_data_390,phv_data_391}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_599 = 8'hc1 == _GEN_86 ? _groups_0_T_35 : _GEN_598; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_36 = {phv_data_392,phv_data_393,phv_data_394,phv_data_395}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_600 = 8'hc2 == _GEN_86 ? _groups_0_T_36 : _GEN_599; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_37 = {phv_data_396,phv_data_397,phv_data_398,phv_data_399}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_601 = 8'hc3 == _GEN_86 ? _groups_0_T_37 : _GEN_600; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_38 = {phv_data_400,phv_data_401,phv_data_402,phv_data_403}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_602 = 8'hc4 == _GEN_86 ? _groups_0_T_38 : _GEN_601; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_39 = {phv_data_404,phv_data_405,phv_data_406,phv_data_407}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_603 = 8'hc5 == _GEN_86 ? _groups_0_T_39 : _GEN_602; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_40 = {phv_data_408,phv_data_409,phv_data_410,phv_data_411}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_604 = 8'hc6 == _GEN_86 ? _groups_0_T_40 : _GEN_603; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_41 = {phv_data_412,phv_data_413,phv_data_414,phv_data_415}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_605 = 8'hc7 == _GEN_86 ? _groups_0_T_41 : _GEN_604; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_42 = {phv_data_416,phv_data_417,phv_data_418,phv_data_419}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_606 = 8'hc8 == _GEN_86 ? _groups_0_T_42 : _GEN_605; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_43 = {phv_data_420,phv_data_421,phv_data_422,phv_data_423}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_607 = 8'hc9 == _GEN_86 ? _groups_0_T_43 : _GEN_606; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_44 = {phv_data_424,phv_data_425,phv_data_426,phv_data_427}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_608 = 8'hca == _GEN_86 ? _groups_0_T_44 : _GEN_607; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_45 = {phv_data_428,phv_data_429,phv_data_430,phv_data_431}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_609 = 8'hcb == _GEN_86 ? _groups_0_T_45 : _GEN_608; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_46 = {phv_data_432,phv_data_433,phv_data_434,phv_data_435}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_610 = 8'hcc == _GEN_86 ? _groups_0_T_46 : _GEN_609; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_47 = {phv_data_436,phv_data_437,phv_data_438,phv_data_439}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_611 = 8'hcd == _GEN_86 ? _groups_0_T_47 : _GEN_610; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_48 = {phv_data_440,phv_data_441,phv_data_442,phv_data_443}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_612 = 8'hce == _GEN_86 ? _groups_0_T_48 : _GEN_611; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_49 = {phv_data_444,phv_data_445,phv_data_446,phv_data_447}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_613 = 8'hcf == _GEN_86 ? _groups_0_T_49 : _GEN_612; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_50 = {phv_data_448,phv_data_449,phv_data_450,phv_data_451}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_614 = 8'hd0 == _GEN_86 ? _groups_0_T_50 : _GEN_613; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_51 = {phv_data_452,phv_data_453,phv_data_454,phv_data_455}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_615 = 8'hd1 == _GEN_86 ? _groups_0_T_51 : _GEN_614; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_52 = {phv_data_456,phv_data_457,phv_data_458,phv_data_459}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_616 = 8'hd2 == _GEN_86 ? _groups_0_T_52 : _GEN_615; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_53 = {phv_data_460,phv_data_461,phv_data_462,phv_data_463}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_617 = 8'hd3 == _GEN_86 ? _groups_0_T_53 : _GEN_616; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_54 = {phv_data_464,phv_data_465,phv_data_466,phv_data_467}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_618 = 8'hd4 == _GEN_86 ? _groups_0_T_54 : _GEN_617; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_55 = {phv_data_468,phv_data_469,phv_data_470,phv_data_471}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_619 = 8'hd5 == _GEN_86 ? _groups_0_T_55 : _GEN_618; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_56 = {phv_data_472,phv_data_473,phv_data_474,phv_data_475}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_620 = 8'hd6 == _GEN_86 ? _groups_0_T_56 : _GEN_619; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_57 = {phv_data_476,phv_data_477,phv_data_478,phv_data_479}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_621 = 8'hd7 == _GEN_86 ? _groups_0_T_57 : _GEN_620; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_58 = {phv_data_480,phv_data_481,phv_data_482,phv_data_483}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_622 = 8'hd8 == _GEN_86 ? _groups_0_T_58 : _GEN_621; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_59 = {phv_data_484,phv_data_485,phv_data_486,phv_data_487}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_623 = 8'hd9 == _GEN_86 ? _groups_0_T_59 : _GEN_622; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_60 = {phv_data_488,phv_data_489,phv_data_490,phv_data_491}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_624 = 8'hda == _GEN_86 ? _groups_0_T_60 : _GEN_623; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_61 = {phv_data_492,phv_data_493,phv_data_494,phv_data_495}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_625 = 8'hdb == _GEN_86 ? _groups_0_T_61 : _GEN_624; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_62 = {phv_data_496,phv_data_497,phv_data_498,phv_data_499}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_626 = 8'hdc == _GEN_86 ? _groups_0_T_62 : _GEN_625; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_63 = {phv_data_500,phv_data_501,phv_data_502,phv_data_503}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_627 = 8'hdd == _GEN_86 ? _groups_0_T_63 : _GEN_626; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_64 = {phv_data_504,phv_data_505,phv_data_506,phv_data_507}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_628 = 8'hde == _GEN_86 ? _groups_0_T_64 : _GEN_627; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_65 = {phv_data_508,phv_data_509,phv_data_510,phv_data_511}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_629 = 8'hdf == _GEN_86 ? _groups_0_T_65 : _GEN_628; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] groups_0 = _GEN_56 == 2'h3 ? _GEN_629 : _GEN_565; // @[matcher_pisa.scala 155:50]
  wire [7:0] _GEN_631 = 8'h0 == _GEN_90 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_632 = 8'h1 == _GEN_90 ? phv_data_1 : _GEN_631; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_633 = 8'h2 == _GEN_90 ? phv_data_2 : _GEN_632; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_634 = 8'h3 == _GEN_90 ? phv_data_3 : _GEN_633; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_635 = 8'h4 == _GEN_90 ? phv_data_4 : _GEN_634; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_636 = 8'h5 == _GEN_90 ? phv_data_5 : _GEN_635; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_637 = 8'h6 == _GEN_90 ? phv_data_6 : _GEN_636; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_638 = 8'h7 == _GEN_90 ? phv_data_7 : _GEN_637; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_639 = 8'h8 == _GEN_90 ? phv_data_8 : _GEN_638; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_640 = 8'h9 == _GEN_90 ? phv_data_9 : _GEN_639; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_641 = 8'ha == _GEN_90 ? phv_data_10 : _GEN_640; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_642 = 8'hb == _GEN_90 ? phv_data_11 : _GEN_641; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_643 = 8'hc == _GEN_90 ? phv_data_12 : _GEN_642; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_644 = 8'hd == _GEN_90 ? phv_data_13 : _GEN_643; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_645 = 8'he == _GEN_90 ? phv_data_14 : _GEN_644; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_646 = 8'hf == _GEN_90 ? phv_data_15 : _GEN_645; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_647 = 8'h10 == _GEN_90 ? phv_data_16 : _GEN_646; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_648 = 8'h11 == _GEN_90 ? phv_data_17 : _GEN_647; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_649 = 8'h12 == _GEN_90 ? phv_data_18 : _GEN_648; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_650 = 8'h13 == _GEN_90 ? phv_data_19 : _GEN_649; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_651 = 8'h14 == _GEN_90 ? phv_data_20 : _GEN_650; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_652 = 8'h15 == _GEN_90 ? phv_data_21 : _GEN_651; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_653 = 8'h16 == _GEN_90 ? phv_data_22 : _GEN_652; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_654 = 8'h17 == _GEN_90 ? phv_data_23 : _GEN_653; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_655 = 8'h18 == _GEN_90 ? phv_data_24 : _GEN_654; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_656 = 8'h19 == _GEN_90 ? phv_data_25 : _GEN_655; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_657 = 8'h1a == _GEN_90 ? phv_data_26 : _GEN_656; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_658 = 8'h1b == _GEN_90 ? phv_data_27 : _GEN_657; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_659 = 8'h1c == _GEN_90 ? phv_data_28 : _GEN_658; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_660 = 8'h1d == _GEN_90 ? phv_data_29 : _GEN_659; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_661 = 8'h1e == _GEN_90 ? phv_data_30 : _GEN_660; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_662 = 8'h1f == _GEN_90 ? phv_data_31 : _GEN_661; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_663 = 8'h20 == _GEN_90 ? phv_data_32 : _GEN_662; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_664 = 8'h21 == _GEN_90 ? phv_data_33 : _GEN_663; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_665 = 8'h22 == _GEN_90 ? phv_data_34 : _GEN_664; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_666 = 8'h23 == _GEN_90 ? phv_data_35 : _GEN_665; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_667 = 8'h24 == _GEN_90 ? phv_data_36 : _GEN_666; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_668 = 8'h25 == _GEN_90 ? phv_data_37 : _GEN_667; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_669 = 8'h26 == _GEN_90 ? phv_data_38 : _GEN_668; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_670 = 8'h27 == _GEN_90 ? phv_data_39 : _GEN_669; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_671 = 8'h28 == _GEN_90 ? phv_data_40 : _GEN_670; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_672 = 8'h29 == _GEN_90 ? phv_data_41 : _GEN_671; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_673 = 8'h2a == _GEN_90 ? phv_data_42 : _GEN_672; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_674 = 8'h2b == _GEN_90 ? phv_data_43 : _GEN_673; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_675 = 8'h2c == _GEN_90 ? phv_data_44 : _GEN_674; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_676 = 8'h2d == _GEN_90 ? phv_data_45 : _GEN_675; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_677 = 8'h2e == _GEN_90 ? phv_data_46 : _GEN_676; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_678 = 8'h2f == _GEN_90 ? phv_data_47 : _GEN_677; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_679 = 8'h30 == _GEN_90 ? phv_data_48 : _GEN_678; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_680 = 8'h31 == _GEN_90 ? phv_data_49 : _GEN_679; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_681 = 8'h32 == _GEN_90 ? phv_data_50 : _GEN_680; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_682 = 8'h33 == _GEN_90 ? phv_data_51 : _GEN_681; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_683 = 8'h34 == _GEN_90 ? phv_data_52 : _GEN_682; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_684 = 8'h35 == _GEN_90 ? phv_data_53 : _GEN_683; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_685 = 8'h36 == _GEN_90 ? phv_data_54 : _GEN_684; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_686 = 8'h37 == _GEN_90 ? phv_data_55 : _GEN_685; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_687 = 8'h38 == _GEN_90 ? phv_data_56 : _GEN_686; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_688 = 8'h39 == _GEN_90 ? phv_data_57 : _GEN_687; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_689 = 8'h3a == _GEN_90 ? phv_data_58 : _GEN_688; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_690 = 8'h3b == _GEN_90 ? phv_data_59 : _GEN_689; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_691 = 8'h3c == _GEN_90 ? phv_data_60 : _GEN_690; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_692 = 8'h3d == _GEN_90 ? phv_data_61 : _GEN_691; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_693 = 8'h3e == _GEN_90 ? phv_data_62 : _GEN_692; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_694 = 8'h3f == _GEN_90 ? phv_data_63 : _GEN_693; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] bytes_1_0 = _GEN_66 ? _GEN_694 : 8'h0; // @[matcher_pisa.scala 129:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_696 = 8'h0 == _GEN_91 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_697 = 8'h1 == _GEN_91 ? phv_data_1 : _GEN_696; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_698 = 8'h2 == _GEN_91 ? phv_data_2 : _GEN_697; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_699 = 8'h3 == _GEN_91 ? phv_data_3 : _GEN_698; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_700 = 8'h4 == _GEN_91 ? phv_data_4 : _GEN_699; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_701 = 8'h5 == _GEN_91 ? phv_data_5 : _GEN_700; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_702 = 8'h6 == _GEN_91 ? phv_data_6 : _GEN_701; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_703 = 8'h7 == _GEN_91 ? phv_data_7 : _GEN_702; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_704 = 8'h8 == _GEN_91 ? phv_data_8 : _GEN_703; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_705 = 8'h9 == _GEN_91 ? phv_data_9 : _GEN_704; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_706 = 8'ha == _GEN_91 ? phv_data_10 : _GEN_705; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_707 = 8'hb == _GEN_91 ? phv_data_11 : _GEN_706; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_708 = 8'hc == _GEN_91 ? phv_data_12 : _GEN_707; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_709 = 8'hd == _GEN_91 ? phv_data_13 : _GEN_708; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_710 = 8'he == _GEN_91 ? phv_data_14 : _GEN_709; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_711 = 8'hf == _GEN_91 ? phv_data_15 : _GEN_710; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_712 = 8'h10 == _GEN_91 ? phv_data_16 : _GEN_711; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_713 = 8'h11 == _GEN_91 ? phv_data_17 : _GEN_712; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_714 = 8'h12 == _GEN_91 ? phv_data_18 : _GEN_713; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_715 = 8'h13 == _GEN_91 ? phv_data_19 : _GEN_714; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_716 = 8'h14 == _GEN_91 ? phv_data_20 : _GEN_715; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_717 = 8'h15 == _GEN_91 ? phv_data_21 : _GEN_716; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_718 = 8'h16 == _GEN_91 ? phv_data_22 : _GEN_717; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_719 = 8'h17 == _GEN_91 ? phv_data_23 : _GEN_718; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_720 = 8'h18 == _GEN_91 ? phv_data_24 : _GEN_719; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_721 = 8'h19 == _GEN_91 ? phv_data_25 : _GEN_720; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_722 = 8'h1a == _GEN_91 ? phv_data_26 : _GEN_721; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_723 = 8'h1b == _GEN_91 ? phv_data_27 : _GEN_722; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_724 = 8'h1c == _GEN_91 ? phv_data_28 : _GEN_723; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_725 = 8'h1d == _GEN_91 ? phv_data_29 : _GEN_724; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_726 = 8'h1e == _GEN_91 ? phv_data_30 : _GEN_725; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_727 = 8'h1f == _GEN_91 ? phv_data_31 : _GEN_726; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_728 = 8'h20 == _GEN_91 ? phv_data_32 : _GEN_727; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_729 = 8'h21 == _GEN_91 ? phv_data_33 : _GEN_728; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_730 = 8'h22 == _GEN_91 ? phv_data_34 : _GEN_729; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_731 = 8'h23 == _GEN_91 ? phv_data_35 : _GEN_730; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_732 = 8'h24 == _GEN_91 ? phv_data_36 : _GEN_731; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_733 = 8'h25 == _GEN_91 ? phv_data_37 : _GEN_732; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_734 = 8'h26 == _GEN_91 ? phv_data_38 : _GEN_733; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_735 = 8'h27 == _GEN_91 ? phv_data_39 : _GEN_734; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_736 = 8'h28 == _GEN_91 ? phv_data_40 : _GEN_735; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_737 = 8'h29 == _GEN_91 ? phv_data_41 : _GEN_736; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_738 = 8'h2a == _GEN_91 ? phv_data_42 : _GEN_737; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_739 = 8'h2b == _GEN_91 ? phv_data_43 : _GEN_738; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_740 = 8'h2c == _GEN_91 ? phv_data_44 : _GEN_739; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_741 = 8'h2d == _GEN_91 ? phv_data_45 : _GEN_740; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_742 = 8'h2e == _GEN_91 ? phv_data_46 : _GEN_741; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_743 = 8'h2f == _GEN_91 ? phv_data_47 : _GEN_742; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_744 = 8'h30 == _GEN_91 ? phv_data_48 : _GEN_743; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_745 = 8'h31 == _GEN_91 ? phv_data_49 : _GEN_744; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_746 = 8'h32 == _GEN_91 ? phv_data_50 : _GEN_745; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_747 = 8'h33 == _GEN_91 ? phv_data_51 : _GEN_746; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_748 = 8'h34 == _GEN_91 ? phv_data_52 : _GEN_747; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_749 = 8'h35 == _GEN_91 ? phv_data_53 : _GEN_748; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_750 = 8'h36 == _GEN_91 ? phv_data_54 : _GEN_749; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_751 = 8'h37 == _GEN_91 ? phv_data_55 : _GEN_750; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_752 = 8'h38 == _GEN_91 ? phv_data_56 : _GEN_751; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_753 = 8'h39 == _GEN_91 ? phv_data_57 : _GEN_752; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_754 = 8'h3a == _GEN_91 ? phv_data_58 : _GEN_753; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_755 = 8'h3b == _GEN_91 ? phv_data_59 : _GEN_754; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_756 = 8'h3c == _GEN_91 ? phv_data_60 : _GEN_755; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_757 = 8'h3d == _GEN_91 ? phv_data_61 : _GEN_756; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_758 = 8'h3e == _GEN_91 ? phv_data_62 : _GEN_757; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_759 = 8'h3f == _GEN_91 ? phv_data_63 : _GEN_758; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] bytes_1_1 = _GEN_67 ? _GEN_759 : 8'h0; // @[matcher_pisa.scala 129:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_761 = 8'h0 == _GEN_92 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_762 = 8'h1 == _GEN_92 ? phv_data_1 : _GEN_761; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_763 = 8'h2 == _GEN_92 ? phv_data_2 : _GEN_762; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_764 = 8'h3 == _GEN_92 ? phv_data_3 : _GEN_763; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_765 = 8'h4 == _GEN_92 ? phv_data_4 : _GEN_764; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_766 = 8'h5 == _GEN_92 ? phv_data_5 : _GEN_765; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_767 = 8'h6 == _GEN_92 ? phv_data_6 : _GEN_766; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_768 = 8'h7 == _GEN_92 ? phv_data_7 : _GEN_767; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_769 = 8'h8 == _GEN_92 ? phv_data_8 : _GEN_768; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_770 = 8'h9 == _GEN_92 ? phv_data_9 : _GEN_769; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_771 = 8'ha == _GEN_92 ? phv_data_10 : _GEN_770; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_772 = 8'hb == _GEN_92 ? phv_data_11 : _GEN_771; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_773 = 8'hc == _GEN_92 ? phv_data_12 : _GEN_772; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_774 = 8'hd == _GEN_92 ? phv_data_13 : _GEN_773; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_775 = 8'he == _GEN_92 ? phv_data_14 : _GEN_774; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_776 = 8'hf == _GEN_92 ? phv_data_15 : _GEN_775; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_777 = 8'h10 == _GEN_92 ? phv_data_16 : _GEN_776; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_778 = 8'h11 == _GEN_92 ? phv_data_17 : _GEN_777; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_779 = 8'h12 == _GEN_92 ? phv_data_18 : _GEN_778; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_780 = 8'h13 == _GEN_92 ? phv_data_19 : _GEN_779; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_781 = 8'h14 == _GEN_92 ? phv_data_20 : _GEN_780; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_782 = 8'h15 == _GEN_92 ? phv_data_21 : _GEN_781; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_783 = 8'h16 == _GEN_92 ? phv_data_22 : _GEN_782; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_784 = 8'h17 == _GEN_92 ? phv_data_23 : _GEN_783; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_785 = 8'h18 == _GEN_92 ? phv_data_24 : _GEN_784; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_786 = 8'h19 == _GEN_92 ? phv_data_25 : _GEN_785; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_787 = 8'h1a == _GEN_92 ? phv_data_26 : _GEN_786; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_788 = 8'h1b == _GEN_92 ? phv_data_27 : _GEN_787; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_789 = 8'h1c == _GEN_92 ? phv_data_28 : _GEN_788; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_790 = 8'h1d == _GEN_92 ? phv_data_29 : _GEN_789; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_791 = 8'h1e == _GEN_92 ? phv_data_30 : _GEN_790; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_792 = 8'h1f == _GEN_92 ? phv_data_31 : _GEN_791; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_793 = 8'h20 == _GEN_92 ? phv_data_32 : _GEN_792; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_794 = 8'h21 == _GEN_92 ? phv_data_33 : _GEN_793; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_795 = 8'h22 == _GEN_92 ? phv_data_34 : _GEN_794; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_796 = 8'h23 == _GEN_92 ? phv_data_35 : _GEN_795; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_797 = 8'h24 == _GEN_92 ? phv_data_36 : _GEN_796; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_798 = 8'h25 == _GEN_92 ? phv_data_37 : _GEN_797; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_799 = 8'h26 == _GEN_92 ? phv_data_38 : _GEN_798; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_800 = 8'h27 == _GEN_92 ? phv_data_39 : _GEN_799; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_801 = 8'h28 == _GEN_92 ? phv_data_40 : _GEN_800; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_802 = 8'h29 == _GEN_92 ? phv_data_41 : _GEN_801; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_803 = 8'h2a == _GEN_92 ? phv_data_42 : _GEN_802; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_804 = 8'h2b == _GEN_92 ? phv_data_43 : _GEN_803; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_805 = 8'h2c == _GEN_92 ? phv_data_44 : _GEN_804; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_806 = 8'h2d == _GEN_92 ? phv_data_45 : _GEN_805; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_807 = 8'h2e == _GEN_92 ? phv_data_46 : _GEN_806; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_808 = 8'h2f == _GEN_92 ? phv_data_47 : _GEN_807; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_809 = 8'h30 == _GEN_92 ? phv_data_48 : _GEN_808; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_810 = 8'h31 == _GEN_92 ? phv_data_49 : _GEN_809; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_811 = 8'h32 == _GEN_92 ? phv_data_50 : _GEN_810; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_812 = 8'h33 == _GEN_92 ? phv_data_51 : _GEN_811; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_813 = 8'h34 == _GEN_92 ? phv_data_52 : _GEN_812; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_814 = 8'h35 == _GEN_92 ? phv_data_53 : _GEN_813; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_815 = 8'h36 == _GEN_92 ? phv_data_54 : _GEN_814; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_816 = 8'h37 == _GEN_92 ? phv_data_55 : _GEN_815; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_817 = 8'h38 == _GEN_92 ? phv_data_56 : _GEN_816; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_818 = 8'h39 == _GEN_92 ? phv_data_57 : _GEN_817; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_819 = 8'h3a == _GEN_92 ? phv_data_58 : _GEN_818; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_820 = 8'h3b == _GEN_92 ? phv_data_59 : _GEN_819; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_821 = 8'h3c == _GEN_92 ? phv_data_60 : _GEN_820; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_822 = 8'h3d == _GEN_92 ? phv_data_61 : _GEN_821; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_823 = 8'h3e == _GEN_92 ? phv_data_62 : _GEN_822; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_824 = 8'h3f == _GEN_92 ? phv_data_63 : _GEN_823; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] bytes_1_2 = _GEN_68 ? _GEN_824 : 8'h0; // @[matcher_pisa.scala 129:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_826 = 8'h0 == _GEN_93 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_827 = 8'h1 == _GEN_93 ? phv_data_1 : _GEN_826; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_828 = 8'h2 == _GEN_93 ? phv_data_2 : _GEN_827; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_829 = 8'h3 == _GEN_93 ? phv_data_3 : _GEN_828; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_830 = 8'h4 == _GEN_93 ? phv_data_4 : _GEN_829; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_831 = 8'h5 == _GEN_93 ? phv_data_5 : _GEN_830; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_832 = 8'h6 == _GEN_93 ? phv_data_6 : _GEN_831; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_833 = 8'h7 == _GEN_93 ? phv_data_7 : _GEN_832; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_834 = 8'h8 == _GEN_93 ? phv_data_8 : _GEN_833; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_835 = 8'h9 == _GEN_93 ? phv_data_9 : _GEN_834; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_836 = 8'ha == _GEN_93 ? phv_data_10 : _GEN_835; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_837 = 8'hb == _GEN_93 ? phv_data_11 : _GEN_836; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_838 = 8'hc == _GEN_93 ? phv_data_12 : _GEN_837; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_839 = 8'hd == _GEN_93 ? phv_data_13 : _GEN_838; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_840 = 8'he == _GEN_93 ? phv_data_14 : _GEN_839; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_841 = 8'hf == _GEN_93 ? phv_data_15 : _GEN_840; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_842 = 8'h10 == _GEN_93 ? phv_data_16 : _GEN_841; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_843 = 8'h11 == _GEN_93 ? phv_data_17 : _GEN_842; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_844 = 8'h12 == _GEN_93 ? phv_data_18 : _GEN_843; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_845 = 8'h13 == _GEN_93 ? phv_data_19 : _GEN_844; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_846 = 8'h14 == _GEN_93 ? phv_data_20 : _GEN_845; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_847 = 8'h15 == _GEN_93 ? phv_data_21 : _GEN_846; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_848 = 8'h16 == _GEN_93 ? phv_data_22 : _GEN_847; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_849 = 8'h17 == _GEN_93 ? phv_data_23 : _GEN_848; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_850 = 8'h18 == _GEN_93 ? phv_data_24 : _GEN_849; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_851 = 8'h19 == _GEN_93 ? phv_data_25 : _GEN_850; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_852 = 8'h1a == _GEN_93 ? phv_data_26 : _GEN_851; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_853 = 8'h1b == _GEN_93 ? phv_data_27 : _GEN_852; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_854 = 8'h1c == _GEN_93 ? phv_data_28 : _GEN_853; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_855 = 8'h1d == _GEN_93 ? phv_data_29 : _GEN_854; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_856 = 8'h1e == _GEN_93 ? phv_data_30 : _GEN_855; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_857 = 8'h1f == _GEN_93 ? phv_data_31 : _GEN_856; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_858 = 8'h20 == _GEN_93 ? phv_data_32 : _GEN_857; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_859 = 8'h21 == _GEN_93 ? phv_data_33 : _GEN_858; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_860 = 8'h22 == _GEN_93 ? phv_data_34 : _GEN_859; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_861 = 8'h23 == _GEN_93 ? phv_data_35 : _GEN_860; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_862 = 8'h24 == _GEN_93 ? phv_data_36 : _GEN_861; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_863 = 8'h25 == _GEN_93 ? phv_data_37 : _GEN_862; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_864 = 8'h26 == _GEN_93 ? phv_data_38 : _GEN_863; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_865 = 8'h27 == _GEN_93 ? phv_data_39 : _GEN_864; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_866 = 8'h28 == _GEN_93 ? phv_data_40 : _GEN_865; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_867 = 8'h29 == _GEN_93 ? phv_data_41 : _GEN_866; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_868 = 8'h2a == _GEN_93 ? phv_data_42 : _GEN_867; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_869 = 8'h2b == _GEN_93 ? phv_data_43 : _GEN_868; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_870 = 8'h2c == _GEN_93 ? phv_data_44 : _GEN_869; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_871 = 8'h2d == _GEN_93 ? phv_data_45 : _GEN_870; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_872 = 8'h2e == _GEN_93 ? phv_data_46 : _GEN_871; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_873 = 8'h2f == _GEN_93 ? phv_data_47 : _GEN_872; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_874 = 8'h30 == _GEN_93 ? phv_data_48 : _GEN_873; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_875 = 8'h31 == _GEN_93 ? phv_data_49 : _GEN_874; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_876 = 8'h32 == _GEN_93 ? phv_data_50 : _GEN_875; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_877 = 8'h33 == _GEN_93 ? phv_data_51 : _GEN_876; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_878 = 8'h34 == _GEN_93 ? phv_data_52 : _GEN_877; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_879 = 8'h35 == _GEN_93 ? phv_data_53 : _GEN_878; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_880 = 8'h36 == _GEN_93 ? phv_data_54 : _GEN_879; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_881 = 8'h37 == _GEN_93 ? phv_data_55 : _GEN_880; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_882 = 8'h38 == _GEN_93 ? phv_data_56 : _GEN_881; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_883 = 8'h39 == _GEN_93 ? phv_data_57 : _GEN_882; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_884 = 8'h3a == _GEN_93 ? phv_data_58 : _GEN_883; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_885 = 8'h3b == _GEN_93 ? phv_data_59 : _GEN_884; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_886 = 8'h3c == _GEN_93 ? phv_data_60 : _GEN_885; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_887 = 8'h3d == _GEN_93 ? phv_data_61 : _GEN_886; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_888 = 8'h3e == _GEN_93 ? phv_data_62 : _GEN_887; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_889 = 8'h3f == _GEN_93 ? phv_data_63 : _GEN_888; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] bytes_1_3 = _GEN_69 ? _GEN_889 : 8'h0; // @[matcher_pisa.scala 129:46 matcher_pisa.scala 128:34]
  wire [31:0] _groups_1_T = {bytes_1_0,bytes_1_1,bytes_1_2,bytes_1_3}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_891 = _GEN_57 == 2'h1 ? _groups_1_T : 32'h0; // @[matcher_pisa.scala 123:50 matcher_pisa.scala 137:31 matcher_pisa.scala 122:27]
  wire [15:0] _GEN_892 = 8'h40 == _GEN_90 ? _double_bytes_0_T : 16'h0; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53 matcher_pisa.scala 144:41]
  wire [15:0] _GEN_893 = 8'h41 == _GEN_90 ? _double_bytes_0_T_1 : _GEN_892; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_894 = 8'h42 == _GEN_90 ? _double_bytes_0_T_2 : _GEN_893; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_895 = 8'h43 == _GEN_90 ? _double_bytes_0_T_3 : _GEN_894; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_896 = 8'h44 == _GEN_90 ? _double_bytes_0_T_4 : _GEN_895; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_897 = 8'h45 == _GEN_90 ? _double_bytes_0_T_5 : _GEN_896; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_898 = 8'h46 == _GEN_90 ? _double_bytes_0_T_6 : _GEN_897; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_899 = 8'h47 == _GEN_90 ? _double_bytes_0_T_7 : _GEN_898; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_900 = 8'h48 == _GEN_90 ? _double_bytes_0_T_8 : _GEN_899; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_901 = 8'h49 == _GEN_90 ? _double_bytes_0_T_9 : _GEN_900; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_902 = 8'h4a == _GEN_90 ? _double_bytes_0_T_10 : _GEN_901; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_903 = 8'h4b == _GEN_90 ? _double_bytes_0_T_11 : _GEN_902; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_904 = 8'h4c == _GEN_90 ? _double_bytes_0_T_12 : _GEN_903; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_905 = 8'h4d == _GEN_90 ? _double_bytes_0_T_13 : _GEN_904; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_906 = 8'h4e == _GEN_90 ? _double_bytes_0_T_14 : _GEN_905; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_907 = 8'h4f == _GEN_90 ? _double_bytes_0_T_15 : _GEN_906; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_908 = 8'h50 == _GEN_90 ? _double_bytes_0_T_16 : _GEN_907; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_909 = 8'h51 == _GEN_90 ? _double_bytes_0_T_17 : _GEN_908; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_910 = 8'h52 == _GEN_90 ? _double_bytes_0_T_18 : _GEN_909; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_911 = 8'h53 == _GEN_90 ? _double_bytes_0_T_19 : _GEN_910; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_912 = 8'h54 == _GEN_90 ? _double_bytes_0_T_20 : _GEN_911; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_913 = 8'h55 == _GEN_90 ? _double_bytes_0_T_21 : _GEN_912; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_914 = 8'h56 == _GEN_90 ? _double_bytes_0_T_22 : _GEN_913; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_915 = 8'h57 == _GEN_90 ? _double_bytes_0_T_23 : _GEN_914; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_916 = 8'h58 == _GEN_90 ? _double_bytes_0_T_24 : _GEN_915; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_917 = 8'h59 == _GEN_90 ? _double_bytes_0_T_25 : _GEN_916; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_918 = 8'h5a == _GEN_90 ? _double_bytes_0_T_26 : _GEN_917; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_919 = 8'h5b == _GEN_90 ? _double_bytes_0_T_27 : _GEN_918; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_920 = 8'h5c == _GEN_90 ? _double_bytes_0_T_28 : _GEN_919; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_921 = 8'h5d == _GEN_90 ? _double_bytes_0_T_29 : _GEN_920; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_922 = 8'h5e == _GEN_90 ? _double_bytes_0_T_30 : _GEN_921; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_923 = 8'h5f == _GEN_90 ? _double_bytes_0_T_31 : _GEN_922; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_924 = 8'h60 == _GEN_90 ? _double_bytes_0_T_32 : _GEN_923; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_925 = 8'h61 == _GEN_90 ? _double_bytes_0_T_33 : _GEN_924; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_926 = 8'h62 == _GEN_90 ? _double_bytes_0_T_34 : _GEN_925; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_927 = 8'h63 == _GEN_90 ? _double_bytes_0_T_35 : _GEN_926; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_928 = 8'h64 == _GEN_90 ? _double_bytes_0_T_36 : _GEN_927; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_929 = 8'h65 == _GEN_90 ? _double_bytes_0_T_37 : _GEN_928; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_930 = 8'h66 == _GEN_90 ? _double_bytes_0_T_38 : _GEN_929; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_931 = 8'h67 == _GEN_90 ? _double_bytes_0_T_39 : _GEN_930; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_932 = 8'h68 == _GEN_90 ? _double_bytes_0_T_40 : _GEN_931; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_933 = 8'h69 == _GEN_90 ? _double_bytes_0_T_41 : _GEN_932; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_934 = 8'h6a == _GEN_90 ? _double_bytes_0_T_42 : _GEN_933; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_935 = 8'h6b == _GEN_90 ? _double_bytes_0_T_43 : _GEN_934; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_936 = 8'h6c == _GEN_90 ? _double_bytes_0_T_44 : _GEN_935; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_937 = 8'h6d == _GEN_90 ? _double_bytes_0_T_45 : _GEN_936; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_938 = 8'h6e == _GEN_90 ? _double_bytes_0_T_46 : _GEN_937; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_939 = 8'h6f == _GEN_90 ? _double_bytes_0_T_47 : _GEN_938; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_940 = 8'h70 == _GEN_90 ? _double_bytes_0_T_48 : _GEN_939; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_941 = 8'h71 == _GEN_90 ? _double_bytes_0_T_49 : _GEN_940; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_942 = 8'h72 == _GEN_90 ? _double_bytes_0_T_50 : _GEN_941; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_943 = 8'h73 == _GEN_90 ? _double_bytes_0_T_51 : _GEN_942; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_944 = 8'h74 == _GEN_90 ? _double_bytes_0_T_52 : _GEN_943; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_945 = 8'h75 == _GEN_90 ? _double_bytes_0_T_53 : _GEN_944; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_946 = 8'h76 == _GEN_90 ? _double_bytes_0_T_54 : _GEN_945; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_947 = 8'h77 == _GEN_90 ? _double_bytes_0_T_55 : _GEN_946; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_948 = 8'h78 == _GEN_90 ? _double_bytes_0_T_56 : _GEN_947; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_949 = 8'h79 == _GEN_90 ? _double_bytes_0_T_57 : _GEN_948; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_950 = 8'h7a == _GEN_90 ? _double_bytes_0_T_58 : _GEN_949; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_951 = 8'h7b == _GEN_90 ? _double_bytes_0_T_59 : _GEN_950; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_952 = 8'h7c == _GEN_90 ? _double_bytes_0_T_60 : _GEN_951; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_953 = 8'h7d == _GEN_90 ? _double_bytes_0_T_61 : _GEN_952; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_954 = 8'h7e == _GEN_90 ? _double_bytes_0_T_62 : _GEN_953; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_955 = 8'h7f == _GEN_90 ? _double_bytes_0_T_63 : _GEN_954; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_956 = 8'h80 == _GEN_90 ? _double_bytes_0_T_64 : _GEN_955; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_957 = 8'h81 == _GEN_90 ? _double_bytes_0_T_65 : _GEN_956; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_958 = 8'h82 == _GEN_90 ? _double_bytes_0_T_66 : _GEN_957; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_959 = 8'h83 == _GEN_90 ? _double_bytes_0_T_67 : _GEN_958; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_960 = 8'h84 == _GEN_90 ? _double_bytes_0_T_68 : _GEN_959; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_961 = 8'h85 == _GEN_90 ? _double_bytes_0_T_69 : _GEN_960; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_962 = 8'h86 == _GEN_90 ? _double_bytes_0_T_70 : _GEN_961; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_963 = 8'h87 == _GEN_90 ? _double_bytes_0_T_71 : _GEN_962; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_964 = 8'h88 == _GEN_90 ? _double_bytes_0_T_72 : _GEN_963; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_965 = 8'h89 == _GEN_90 ? _double_bytes_0_T_73 : _GEN_964; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_966 = 8'h8a == _GEN_90 ? _double_bytes_0_T_74 : _GEN_965; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_967 = 8'h8b == _GEN_90 ? _double_bytes_0_T_75 : _GEN_966; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_968 = 8'h8c == _GEN_90 ? _double_bytes_0_T_76 : _GEN_967; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_969 = 8'h8d == _GEN_90 ? _double_bytes_0_T_77 : _GEN_968; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_970 = 8'h8e == _GEN_90 ? _double_bytes_0_T_78 : _GEN_969; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_971 = 8'h8f == _GEN_90 ? _double_bytes_0_T_79 : _GEN_970; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_972 = 8'h90 == _GEN_90 ? _double_bytes_0_T_80 : _GEN_971; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_973 = 8'h91 == _GEN_90 ? _double_bytes_0_T_81 : _GEN_972; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_974 = 8'h92 == _GEN_90 ? _double_bytes_0_T_82 : _GEN_973; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_975 = 8'h93 == _GEN_90 ? _double_bytes_0_T_83 : _GEN_974; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_976 = 8'h94 == _GEN_90 ? _double_bytes_0_T_84 : _GEN_975; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_977 = 8'h95 == _GEN_90 ? _double_bytes_0_T_85 : _GEN_976; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_978 = 8'h96 == _GEN_90 ? _double_bytes_0_T_86 : _GEN_977; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_979 = 8'h97 == _GEN_90 ? _double_bytes_0_T_87 : _GEN_978; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_980 = 8'h98 == _GEN_90 ? _double_bytes_0_T_88 : _GEN_979; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_981 = 8'h99 == _GEN_90 ? _double_bytes_0_T_89 : _GEN_980; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_982 = 8'h9a == _GEN_90 ? _double_bytes_0_T_90 : _GEN_981; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_983 = 8'h9b == _GEN_90 ? _double_bytes_0_T_91 : _GEN_982; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_984 = 8'h9c == _GEN_90 ? _double_bytes_0_T_92 : _GEN_983; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_985 = 8'h9d == _GEN_90 ? _double_bytes_0_T_93 : _GEN_984; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_986 = 8'h9e == _GEN_90 ? _double_bytes_0_T_94 : _GEN_985; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_987 = 8'h9f == _GEN_90 ? _double_bytes_0_T_95 : _GEN_986; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] double_bytes_1_0 = _GEN_66 ? _GEN_987 : 16'h0; // @[matcher_pisa.scala 145:46 matcher_pisa.scala 144:41]
  wire [15:0] _GEN_989 = 8'h40 == _GEN_91 ? _double_bytes_0_T : 16'h0; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53 matcher_pisa.scala 144:41]
  wire [15:0] _GEN_990 = 8'h41 == _GEN_91 ? _double_bytes_0_T_1 : _GEN_989; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_991 = 8'h42 == _GEN_91 ? _double_bytes_0_T_2 : _GEN_990; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_992 = 8'h43 == _GEN_91 ? _double_bytes_0_T_3 : _GEN_991; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_993 = 8'h44 == _GEN_91 ? _double_bytes_0_T_4 : _GEN_992; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_994 = 8'h45 == _GEN_91 ? _double_bytes_0_T_5 : _GEN_993; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_995 = 8'h46 == _GEN_91 ? _double_bytes_0_T_6 : _GEN_994; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_996 = 8'h47 == _GEN_91 ? _double_bytes_0_T_7 : _GEN_995; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_997 = 8'h48 == _GEN_91 ? _double_bytes_0_T_8 : _GEN_996; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_998 = 8'h49 == _GEN_91 ? _double_bytes_0_T_9 : _GEN_997; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_999 = 8'h4a == _GEN_91 ? _double_bytes_0_T_10 : _GEN_998; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1000 = 8'h4b == _GEN_91 ? _double_bytes_0_T_11 : _GEN_999; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1001 = 8'h4c == _GEN_91 ? _double_bytes_0_T_12 : _GEN_1000; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1002 = 8'h4d == _GEN_91 ? _double_bytes_0_T_13 : _GEN_1001; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1003 = 8'h4e == _GEN_91 ? _double_bytes_0_T_14 : _GEN_1002; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1004 = 8'h4f == _GEN_91 ? _double_bytes_0_T_15 : _GEN_1003; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1005 = 8'h50 == _GEN_91 ? _double_bytes_0_T_16 : _GEN_1004; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1006 = 8'h51 == _GEN_91 ? _double_bytes_0_T_17 : _GEN_1005; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1007 = 8'h52 == _GEN_91 ? _double_bytes_0_T_18 : _GEN_1006; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1008 = 8'h53 == _GEN_91 ? _double_bytes_0_T_19 : _GEN_1007; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1009 = 8'h54 == _GEN_91 ? _double_bytes_0_T_20 : _GEN_1008; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1010 = 8'h55 == _GEN_91 ? _double_bytes_0_T_21 : _GEN_1009; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1011 = 8'h56 == _GEN_91 ? _double_bytes_0_T_22 : _GEN_1010; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1012 = 8'h57 == _GEN_91 ? _double_bytes_0_T_23 : _GEN_1011; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1013 = 8'h58 == _GEN_91 ? _double_bytes_0_T_24 : _GEN_1012; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1014 = 8'h59 == _GEN_91 ? _double_bytes_0_T_25 : _GEN_1013; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1015 = 8'h5a == _GEN_91 ? _double_bytes_0_T_26 : _GEN_1014; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1016 = 8'h5b == _GEN_91 ? _double_bytes_0_T_27 : _GEN_1015; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1017 = 8'h5c == _GEN_91 ? _double_bytes_0_T_28 : _GEN_1016; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1018 = 8'h5d == _GEN_91 ? _double_bytes_0_T_29 : _GEN_1017; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1019 = 8'h5e == _GEN_91 ? _double_bytes_0_T_30 : _GEN_1018; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1020 = 8'h5f == _GEN_91 ? _double_bytes_0_T_31 : _GEN_1019; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1021 = 8'h60 == _GEN_91 ? _double_bytes_0_T_32 : _GEN_1020; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1022 = 8'h61 == _GEN_91 ? _double_bytes_0_T_33 : _GEN_1021; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1023 = 8'h62 == _GEN_91 ? _double_bytes_0_T_34 : _GEN_1022; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1024 = 8'h63 == _GEN_91 ? _double_bytes_0_T_35 : _GEN_1023; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1025 = 8'h64 == _GEN_91 ? _double_bytes_0_T_36 : _GEN_1024; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1026 = 8'h65 == _GEN_91 ? _double_bytes_0_T_37 : _GEN_1025; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1027 = 8'h66 == _GEN_91 ? _double_bytes_0_T_38 : _GEN_1026; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1028 = 8'h67 == _GEN_91 ? _double_bytes_0_T_39 : _GEN_1027; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1029 = 8'h68 == _GEN_91 ? _double_bytes_0_T_40 : _GEN_1028; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1030 = 8'h69 == _GEN_91 ? _double_bytes_0_T_41 : _GEN_1029; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1031 = 8'h6a == _GEN_91 ? _double_bytes_0_T_42 : _GEN_1030; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1032 = 8'h6b == _GEN_91 ? _double_bytes_0_T_43 : _GEN_1031; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1033 = 8'h6c == _GEN_91 ? _double_bytes_0_T_44 : _GEN_1032; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1034 = 8'h6d == _GEN_91 ? _double_bytes_0_T_45 : _GEN_1033; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1035 = 8'h6e == _GEN_91 ? _double_bytes_0_T_46 : _GEN_1034; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1036 = 8'h6f == _GEN_91 ? _double_bytes_0_T_47 : _GEN_1035; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1037 = 8'h70 == _GEN_91 ? _double_bytes_0_T_48 : _GEN_1036; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1038 = 8'h71 == _GEN_91 ? _double_bytes_0_T_49 : _GEN_1037; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1039 = 8'h72 == _GEN_91 ? _double_bytes_0_T_50 : _GEN_1038; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1040 = 8'h73 == _GEN_91 ? _double_bytes_0_T_51 : _GEN_1039; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1041 = 8'h74 == _GEN_91 ? _double_bytes_0_T_52 : _GEN_1040; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1042 = 8'h75 == _GEN_91 ? _double_bytes_0_T_53 : _GEN_1041; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1043 = 8'h76 == _GEN_91 ? _double_bytes_0_T_54 : _GEN_1042; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1044 = 8'h77 == _GEN_91 ? _double_bytes_0_T_55 : _GEN_1043; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1045 = 8'h78 == _GEN_91 ? _double_bytes_0_T_56 : _GEN_1044; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1046 = 8'h79 == _GEN_91 ? _double_bytes_0_T_57 : _GEN_1045; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1047 = 8'h7a == _GEN_91 ? _double_bytes_0_T_58 : _GEN_1046; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1048 = 8'h7b == _GEN_91 ? _double_bytes_0_T_59 : _GEN_1047; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1049 = 8'h7c == _GEN_91 ? _double_bytes_0_T_60 : _GEN_1048; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1050 = 8'h7d == _GEN_91 ? _double_bytes_0_T_61 : _GEN_1049; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1051 = 8'h7e == _GEN_91 ? _double_bytes_0_T_62 : _GEN_1050; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1052 = 8'h7f == _GEN_91 ? _double_bytes_0_T_63 : _GEN_1051; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1053 = 8'h80 == _GEN_91 ? _double_bytes_0_T_64 : _GEN_1052; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1054 = 8'h81 == _GEN_91 ? _double_bytes_0_T_65 : _GEN_1053; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1055 = 8'h82 == _GEN_91 ? _double_bytes_0_T_66 : _GEN_1054; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1056 = 8'h83 == _GEN_91 ? _double_bytes_0_T_67 : _GEN_1055; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1057 = 8'h84 == _GEN_91 ? _double_bytes_0_T_68 : _GEN_1056; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1058 = 8'h85 == _GEN_91 ? _double_bytes_0_T_69 : _GEN_1057; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1059 = 8'h86 == _GEN_91 ? _double_bytes_0_T_70 : _GEN_1058; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1060 = 8'h87 == _GEN_91 ? _double_bytes_0_T_71 : _GEN_1059; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1061 = 8'h88 == _GEN_91 ? _double_bytes_0_T_72 : _GEN_1060; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1062 = 8'h89 == _GEN_91 ? _double_bytes_0_T_73 : _GEN_1061; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1063 = 8'h8a == _GEN_91 ? _double_bytes_0_T_74 : _GEN_1062; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1064 = 8'h8b == _GEN_91 ? _double_bytes_0_T_75 : _GEN_1063; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1065 = 8'h8c == _GEN_91 ? _double_bytes_0_T_76 : _GEN_1064; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1066 = 8'h8d == _GEN_91 ? _double_bytes_0_T_77 : _GEN_1065; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1067 = 8'h8e == _GEN_91 ? _double_bytes_0_T_78 : _GEN_1066; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1068 = 8'h8f == _GEN_91 ? _double_bytes_0_T_79 : _GEN_1067; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1069 = 8'h90 == _GEN_91 ? _double_bytes_0_T_80 : _GEN_1068; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1070 = 8'h91 == _GEN_91 ? _double_bytes_0_T_81 : _GEN_1069; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1071 = 8'h92 == _GEN_91 ? _double_bytes_0_T_82 : _GEN_1070; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1072 = 8'h93 == _GEN_91 ? _double_bytes_0_T_83 : _GEN_1071; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1073 = 8'h94 == _GEN_91 ? _double_bytes_0_T_84 : _GEN_1072; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1074 = 8'h95 == _GEN_91 ? _double_bytes_0_T_85 : _GEN_1073; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1075 = 8'h96 == _GEN_91 ? _double_bytes_0_T_86 : _GEN_1074; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1076 = 8'h97 == _GEN_91 ? _double_bytes_0_T_87 : _GEN_1075; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1077 = 8'h98 == _GEN_91 ? _double_bytes_0_T_88 : _GEN_1076; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1078 = 8'h99 == _GEN_91 ? _double_bytes_0_T_89 : _GEN_1077; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1079 = 8'h9a == _GEN_91 ? _double_bytes_0_T_90 : _GEN_1078; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1080 = 8'h9b == _GEN_91 ? _double_bytes_0_T_91 : _GEN_1079; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1081 = 8'h9c == _GEN_91 ? _double_bytes_0_T_92 : _GEN_1080; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1082 = 8'h9d == _GEN_91 ? _double_bytes_0_T_93 : _GEN_1081; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1083 = 8'h9e == _GEN_91 ? _double_bytes_0_T_94 : _GEN_1082; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1084 = 8'h9f == _GEN_91 ? _double_bytes_0_T_95 : _GEN_1083; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] double_bytes_1_1 = _GEN_67 ? _GEN_1084 : 16'h0; // @[matcher_pisa.scala 145:46 matcher_pisa.scala 144:41]
  wire [31:0] _groups_1_T_1 = {double_bytes_1_0,double_bytes_1_1}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_1086 = _GEN_57 == 2'h2 ? _groups_1_T_1 : _GEN_891; // @[matcher_pisa.scala 139:50 matcher_pisa.scala 153:31]
  wire [31:0] _GEN_1087 = 8'ha0 == _GEN_90 ? _groups_0_T_2 : 32'h0; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39 matcher_pisa.scala 158:31]
  wire [31:0] _GEN_1088 = 8'ha1 == _GEN_90 ? _groups_0_T_3 : _GEN_1087; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1089 = 8'ha2 == _GEN_90 ? _groups_0_T_4 : _GEN_1088; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1090 = 8'ha3 == _GEN_90 ? _groups_0_T_5 : _GEN_1089; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1091 = 8'ha4 == _GEN_90 ? _groups_0_T_6 : _GEN_1090; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1092 = 8'ha5 == _GEN_90 ? _groups_0_T_7 : _GEN_1091; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1093 = 8'ha6 == _GEN_90 ? _groups_0_T_8 : _GEN_1092; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1094 = 8'ha7 == _GEN_90 ? _groups_0_T_9 : _GEN_1093; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1095 = 8'ha8 == _GEN_90 ? _groups_0_T_10 : _GEN_1094; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1096 = 8'ha9 == _GEN_90 ? _groups_0_T_11 : _GEN_1095; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1097 = 8'haa == _GEN_90 ? _groups_0_T_12 : _GEN_1096; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1098 = 8'hab == _GEN_90 ? _groups_0_T_13 : _GEN_1097; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1099 = 8'hac == _GEN_90 ? _groups_0_T_14 : _GEN_1098; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1100 = 8'had == _GEN_90 ? _groups_0_T_15 : _GEN_1099; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1101 = 8'hae == _GEN_90 ? _groups_0_T_16 : _GEN_1100; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1102 = 8'haf == _GEN_90 ? _groups_0_T_17 : _GEN_1101; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1103 = 8'hb0 == _GEN_90 ? _groups_0_T_18 : _GEN_1102; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1104 = 8'hb1 == _GEN_90 ? _groups_0_T_19 : _GEN_1103; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1105 = 8'hb2 == _GEN_90 ? _groups_0_T_20 : _GEN_1104; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1106 = 8'hb3 == _GEN_90 ? _groups_0_T_21 : _GEN_1105; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1107 = 8'hb4 == _GEN_90 ? _groups_0_T_22 : _GEN_1106; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1108 = 8'hb5 == _GEN_90 ? _groups_0_T_23 : _GEN_1107; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1109 = 8'hb6 == _GEN_90 ? _groups_0_T_24 : _GEN_1108; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1110 = 8'hb7 == _GEN_90 ? _groups_0_T_25 : _GEN_1109; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1111 = 8'hb8 == _GEN_90 ? _groups_0_T_26 : _GEN_1110; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1112 = 8'hb9 == _GEN_90 ? _groups_0_T_27 : _GEN_1111; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1113 = 8'hba == _GEN_90 ? _groups_0_T_28 : _GEN_1112; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1114 = 8'hbb == _GEN_90 ? _groups_0_T_29 : _GEN_1113; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1115 = 8'hbc == _GEN_90 ? _groups_0_T_30 : _GEN_1114; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1116 = 8'hbd == _GEN_90 ? _groups_0_T_31 : _GEN_1115; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1117 = 8'hbe == _GEN_90 ? _groups_0_T_32 : _GEN_1116; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1118 = 8'hbf == _GEN_90 ? _groups_0_T_33 : _GEN_1117; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1119 = 8'hc0 == _GEN_90 ? _groups_0_T_34 : _GEN_1118; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1120 = 8'hc1 == _GEN_90 ? _groups_0_T_35 : _GEN_1119; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1121 = 8'hc2 == _GEN_90 ? _groups_0_T_36 : _GEN_1120; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1122 = 8'hc3 == _GEN_90 ? _groups_0_T_37 : _GEN_1121; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1123 = 8'hc4 == _GEN_90 ? _groups_0_T_38 : _GEN_1122; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1124 = 8'hc5 == _GEN_90 ? _groups_0_T_39 : _GEN_1123; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1125 = 8'hc6 == _GEN_90 ? _groups_0_T_40 : _GEN_1124; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1126 = 8'hc7 == _GEN_90 ? _groups_0_T_41 : _GEN_1125; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1127 = 8'hc8 == _GEN_90 ? _groups_0_T_42 : _GEN_1126; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1128 = 8'hc9 == _GEN_90 ? _groups_0_T_43 : _GEN_1127; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1129 = 8'hca == _GEN_90 ? _groups_0_T_44 : _GEN_1128; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1130 = 8'hcb == _GEN_90 ? _groups_0_T_45 : _GEN_1129; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1131 = 8'hcc == _GEN_90 ? _groups_0_T_46 : _GEN_1130; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1132 = 8'hcd == _GEN_90 ? _groups_0_T_47 : _GEN_1131; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1133 = 8'hce == _GEN_90 ? _groups_0_T_48 : _GEN_1132; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1134 = 8'hcf == _GEN_90 ? _groups_0_T_49 : _GEN_1133; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1135 = 8'hd0 == _GEN_90 ? _groups_0_T_50 : _GEN_1134; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1136 = 8'hd1 == _GEN_90 ? _groups_0_T_51 : _GEN_1135; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1137 = 8'hd2 == _GEN_90 ? _groups_0_T_52 : _GEN_1136; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1138 = 8'hd3 == _GEN_90 ? _groups_0_T_53 : _GEN_1137; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1139 = 8'hd4 == _GEN_90 ? _groups_0_T_54 : _GEN_1138; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1140 = 8'hd5 == _GEN_90 ? _groups_0_T_55 : _GEN_1139; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1141 = 8'hd6 == _GEN_90 ? _groups_0_T_56 : _GEN_1140; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1142 = 8'hd7 == _GEN_90 ? _groups_0_T_57 : _GEN_1141; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1143 = 8'hd8 == _GEN_90 ? _groups_0_T_58 : _GEN_1142; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1144 = 8'hd9 == _GEN_90 ? _groups_0_T_59 : _GEN_1143; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1145 = 8'hda == _GEN_90 ? _groups_0_T_60 : _GEN_1144; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1146 = 8'hdb == _GEN_90 ? _groups_0_T_61 : _GEN_1145; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1147 = 8'hdc == _GEN_90 ? _groups_0_T_62 : _GEN_1146; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1148 = 8'hdd == _GEN_90 ? _groups_0_T_63 : _GEN_1147; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1149 = 8'hde == _GEN_90 ? _groups_0_T_64 : _GEN_1148; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1150 = 8'hdf == _GEN_90 ? _groups_0_T_65 : _GEN_1149; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] groups_1 = _GEN_57 == 2'h3 ? _GEN_1150 : _GEN_1086; // @[matcher_pisa.scala 155:50]
  wire [7:0] _GEN_1152 = 8'h0 == _GEN_94 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_1153 = 8'h1 == _GEN_94 ? phv_data_1 : _GEN_1152; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1154 = 8'h2 == _GEN_94 ? phv_data_2 : _GEN_1153; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1155 = 8'h3 == _GEN_94 ? phv_data_3 : _GEN_1154; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1156 = 8'h4 == _GEN_94 ? phv_data_4 : _GEN_1155; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1157 = 8'h5 == _GEN_94 ? phv_data_5 : _GEN_1156; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1158 = 8'h6 == _GEN_94 ? phv_data_6 : _GEN_1157; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1159 = 8'h7 == _GEN_94 ? phv_data_7 : _GEN_1158; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1160 = 8'h8 == _GEN_94 ? phv_data_8 : _GEN_1159; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1161 = 8'h9 == _GEN_94 ? phv_data_9 : _GEN_1160; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1162 = 8'ha == _GEN_94 ? phv_data_10 : _GEN_1161; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1163 = 8'hb == _GEN_94 ? phv_data_11 : _GEN_1162; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1164 = 8'hc == _GEN_94 ? phv_data_12 : _GEN_1163; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1165 = 8'hd == _GEN_94 ? phv_data_13 : _GEN_1164; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1166 = 8'he == _GEN_94 ? phv_data_14 : _GEN_1165; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1167 = 8'hf == _GEN_94 ? phv_data_15 : _GEN_1166; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1168 = 8'h10 == _GEN_94 ? phv_data_16 : _GEN_1167; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1169 = 8'h11 == _GEN_94 ? phv_data_17 : _GEN_1168; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1170 = 8'h12 == _GEN_94 ? phv_data_18 : _GEN_1169; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1171 = 8'h13 == _GEN_94 ? phv_data_19 : _GEN_1170; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1172 = 8'h14 == _GEN_94 ? phv_data_20 : _GEN_1171; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1173 = 8'h15 == _GEN_94 ? phv_data_21 : _GEN_1172; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1174 = 8'h16 == _GEN_94 ? phv_data_22 : _GEN_1173; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1175 = 8'h17 == _GEN_94 ? phv_data_23 : _GEN_1174; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1176 = 8'h18 == _GEN_94 ? phv_data_24 : _GEN_1175; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1177 = 8'h19 == _GEN_94 ? phv_data_25 : _GEN_1176; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1178 = 8'h1a == _GEN_94 ? phv_data_26 : _GEN_1177; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1179 = 8'h1b == _GEN_94 ? phv_data_27 : _GEN_1178; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1180 = 8'h1c == _GEN_94 ? phv_data_28 : _GEN_1179; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1181 = 8'h1d == _GEN_94 ? phv_data_29 : _GEN_1180; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1182 = 8'h1e == _GEN_94 ? phv_data_30 : _GEN_1181; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1183 = 8'h1f == _GEN_94 ? phv_data_31 : _GEN_1182; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1184 = 8'h20 == _GEN_94 ? phv_data_32 : _GEN_1183; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1185 = 8'h21 == _GEN_94 ? phv_data_33 : _GEN_1184; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1186 = 8'h22 == _GEN_94 ? phv_data_34 : _GEN_1185; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1187 = 8'h23 == _GEN_94 ? phv_data_35 : _GEN_1186; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1188 = 8'h24 == _GEN_94 ? phv_data_36 : _GEN_1187; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1189 = 8'h25 == _GEN_94 ? phv_data_37 : _GEN_1188; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1190 = 8'h26 == _GEN_94 ? phv_data_38 : _GEN_1189; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1191 = 8'h27 == _GEN_94 ? phv_data_39 : _GEN_1190; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1192 = 8'h28 == _GEN_94 ? phv_data_40 : _GEN_1191; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1193 = 8'h29 == _GEN_94 ? phv_data_41 : _GEN_1192; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1194 = 8'h2a == _GEN_94 ? phv_data_42 : _GEN_1193; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1195 = 8'h2b == _GEN_94 ? phv_data_43 : _GEN_1194; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1196 = 8'h2c == _GEN_94 ? phv_data_44 : _GEN_1195; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1197 = 8'h2d == _GEN_94 ? phv_data_45 : _GEN_1196; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1198 = 8'h2e == _GEN_94 ? phv_data_46 : _GEN_1197; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1199 = 8'h2f == _GEN_94 ? phv_data_47 : _GEN_1198; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1200 = 8'h30 == _GEN_94 ? phv_data_48 : _GEN_1199; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1201 = 8'h31 == _GEN_94 ? phv_data_49 : _GEN_1200; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1202 = 8'h32 == _GEN_94 ? phv_data_50 : _GEN_1201; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1203 = 8'h33 == _GEN_94 ? phv_data_51 : _GEN_1202; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1204 = 8'h34 == _GEN_94 ? phv_data_52 : _GEN_1203; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1205 = 8'h35 == _GEN_94 ? phv_data_53 : _GEN_1204; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1206 = 8'h36 == _GEN_94 ? phv_data_54 : _GEN_1205; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1207 = 8'h37 == _GEN_94 ? phv_data_55 : _GEN_1206; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1208 = 8'h38 == _GEN_94 ? phv_data_56 : _GEN_1207; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1209 = 8'h39 == _GEN_94 ? phv_data_57 : _GEN_1208; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1210 = 8'h3a == _GEN_94 ? phv_data_58 : _GEN_1209; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1211 = 8'h3b == _GEN_94 ? phv_data_59 : _GEN_1210; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1212 = 8'h3c == _GEN_94 ? phv_data_60 : _GEN_1211; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1213 = 8'h3d == _GEN_94 ? phv_data_61 : _GEN_1212; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1214 = 8'h3e == _GEN_94 ? phv_data_62 : _GEN_1213; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1215 = 8'h3f == _GEN_94 ? phv_data_63 : _GEN_1214; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] bytes_2_0 = _GEN_70 ? _GEN_1215 : 8'h0; // @[matcher_pisa.scala 129:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_1217 = 8'h0 == _GEN_95 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_1218 = 8'h1 == _GEN_95 ? phv_data_1 : _GEN_1217; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1219 = 8'h2 == _GEN_95 ? phv_data_2 : _GEN_1218; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1220 = 8'h3 == _GEN_95 ? phv_data_3 : _GEN_1219; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1221 = 8'h4 == _GEN_95 ? phv_data_4 : _GEN_1220; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1222 = 8'h5 == _GEN_95 ? phv_data_5 : _GEN_1221; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1223 = 8'h6 == _GEN_95 ? phv_data_6 : _GEN_1222; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1224 = 8'h7 == _GEN_95 ? phv_data_7 : _GEN_1223; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1225 = 8'h8 == _GEN_95 ? phv_data_8 : _GEN_1224; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1226 = 8'h9 == _GEN_95 ? phv_data_9 : _GEN_1225; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1227 = 8'ha == _GEN_95 ? phv_data_10 : _GEN_1226; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1228 = 8'hb == _GEN_95 ? phv_data_11 : _GEN_1227; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1229 = 8'hc == _GEN_95 ? phv_data_12 : _GEN_1228; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1230 = 8'hd == _GEN_95 ? phv_data_13 : _GEN_1229; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1231 = 8'he == _GEN_95 ? phv_data_14 : _GEN_1230; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1232 = 8'hf == _GEN_95 ? phv_data_15 : _GEN_1231; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1233 = 8'h10 == _GEN_95 ? phv_data_16 : _GEN_1232; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1234 = 8'h11 == _GEN_95 ? phv_data_17 : _GEN_1233; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1235 = 8'h12 == _GEN_95 ? phv_data_18 : _GEN_1234; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1236 = 8'h13 == _GEN_95 ? phv_data_19 : _GEN_1235; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1237 = 8'h14 == _GEN_95 ? phv_data_20 : _GEN_1236; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1238 = 8'h15 == _GEN_95 ? phv_data_21 : _GEN_1237; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1239 = 8'h16 == _GEN_95 ? phv_data_22 : _GEN_1238; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1240 = 8'h17 == _GEN_95 ? phv_data_23 : _GEN_1239; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1241 = 8'h18 == _GEN_95 ? phv_data_24 : _GEN_1240; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1242 = 8'h19 == _GEN_95 ? phv_data_25 : _GEN_1241; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1243 = 8'h1a == _GEN_95 ? phv_data_26 : _GEN_1242; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1244 = 8'h1b == _GEN_95 ? phv_data_27 : _GEN_1243; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1245 = 8'h1c == _GEN_95 ? phv_data_28 : _GEN_1244; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1246 = 8'h1d == _GEN_95 ? phv_data_29 : _GEN_1245; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1247 = 8'h1e == _GEN_95 ? phv_data_30 : _GEN_1246; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1248 = 8'h1f == _GEN_95 ? phv_data_31 : _GEN_1247; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1249 = 8'h20 == _GEN_95 ? phv_data_32 : _GEN_1248; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1250 = 8'h21 == _GEN_95 ? phv_data_33 : _GEN_1249; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1251 = 8'h22 == _GEN_95 ? phv_data_34 : _GEN_1250; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1252 = 8'h23 == _GEN_95 ? phv_data_35 : _GEN_1251; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1253 = 8'h24 == _GEN_95 ? phv_data_36 : _GEN_1252; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1254 = 8'h25 == _GEN_95 ? phv_data_37 : _GEN_1253; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1255 = 8'h26 == _GEN_95 ? phv_data_38 : _GEN_1254; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1256 = 8'h27 == _GEN_95 ? phv_data_39 : _GEN_1255; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1257 = 8'h28 == _GEN_95 ? phv_data_40 : _GEN_1256; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1258 = 8'h29 == _GEN_95 ? phv_data_41 : _GEN_1257; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1259 = 8'h2a == _GEN_95 ? phv_data_42 : _GEN_1258; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1260 = 8'h2b == _GEN_95 ? phv_data_43 : _GEN_1259; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1261 = 8'h2c == _GEN_95 ? phv_data_44 : _GEN_1260; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1262 = 8'h2d == _GEN_95 ? phv_data_45 : _GEN_1261; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1263 = 8'h2e == _GEN_95 ? phv_data_46 : _GEN_1262; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1264 = 8'h2f == _GEN_95 ? phv_data_47 : _GEN_1263; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1265 = 8'h30 == _GEN_95 ? phv_data_48 : _GEN_1264; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1266 = 8'h31 == _GEN_95 ? phv_data_49 : _GEN_1265; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1267 = 8'h32 == _GEN_95 ? phv_data_50 : _GEN_1266; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1268 = 8'h33 == _GEN_95 ? phv_data_51 : _GEN_1267; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1269 = 8'h34 == _GEN_95 ? phv_data_52 : _GEN_1268; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1270 = 8'h35 == _GEN_95 ? phv_data_53 : _GEN_1269; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1271 = 8'h36 == _GEN_95 ? phv_data_54 : _GEN_1270; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1272 = 8'h37 == _GEN_95 ? phv_data_55 : _GEN_1271; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1273 = 8'h38 == _GEN_95 ? phv_data_56 : _GEN_1272; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1274 = 8'h39 == _GEN_95 ? phv_data_57 : _GEN_1273; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1275 = 8'h3a == _GEN_95 ? phv_data_58 : _GEN_1274; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1276 = 8'h3b == _GEN_95 ? phv_data_59 : _GEN_1275; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1277 = 8'h3c == _GEN_95 ? phv_data_60 : _GEN_1276; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1278 = 8'h3d == _GEN_95 ? phv_data_61 : _GEN_1277; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1279 = 8'h3e == _GEN_95 ? phv_data_62 : _GEN_1278; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1280 = 8'h3f == _GEN_95 ? phv_data_63 : _GEN_1279; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] bytes_2_1 = _GEN_71 ? _GEN_1280 : 8'h0; // @[matcher_pisa.scala 129:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_1282 = 8'h0 == _GEN_96 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_1283 = 8'h1 == _GEN_96 ? phv_data_1 : _GEN_1282; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1284 = 8'h2 == _GEN_96 ? phv_data_2 : _GEN_1283; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1285 = 8'h3 == _GEN_96 ? phv_data_3 : _GEN_1284; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1286 = 8'h4 == _GEN_96 ? phv_data_4 : _GEN_1285; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1287 = 8'h5 == _GEN_96 ? phv_data_5 : _GEN_1286; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1288 = 8'h6 == _GEN_96 ? phv_data_6 : _GEN_1287; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1289 = 8'h7 == _GEN_96 ? phv_data_7 : _GEN_1288; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1290 = 8'h8 == _GEN_96 ? phv_data_8 : _GEN_1289; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1291 = 8'h9 == _GEN_96 ? phv_data_9 : _GEN_1290; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1292 = 8'ha == _GEN_96 ? phv_data_10 : _GEN_1291; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1293 = 8'hb == _GEN_96 ? phv_data_11 : _GEN_1292; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1294 = 8'hc == _GEN_96 ? phv_data_12 : _GEN_1293; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1295 = 8'hd == _GEN_96 ? phv_data_13 : _GEN_1294; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1296 = 8'he == _GEN_96 ? phv_data_14 : _GEN_1295; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1297 = 8'hf == _GEN_96 ? phv_data_15 : _GEN_1296; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1298 = 8'h10 == _GEN_96 ? phv_data_16 : _GEN_1297; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1299 = 8'h11 == _GEN_96 ? phv_data_17 : _GEN_1298; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1300 = 8'h12 == _GEN_96 ? phv_data_18 : _GEN_1299; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1301 = 8'h13 == _GEN_96 ? phv_data_19 : _GEN_1300; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1302 = 8'h14 == _GEN_96 ? phv_data_20 : _GEN_1301; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1303 = 8'h15 == _GEN_96 ? phv_data_21 : _GEN_1302; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1304 = 8'h16 == _GEN_96 ? phv_data_22 : _GEN_1303; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1305 = 8'h17 == _GEN_96 ? phv_data_23 : _GEN_1304; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1306 = 8'h18 == _GEN_96 ? phv_data_24 : _GEN_1305; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1307 = 8'h19 == _GEN_96 ? phv_data_25 : _GEN_1306; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1308 = 8'h1a == _GEN_96 ? phv_data_26 : _GEN_1307; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1309 = 8'h1b == _GEN_96 ? phv_data_27 : _GEN_1308; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1310 = 8'h1c == _GEN_96 ? phv_data_28 : _GEN_1309; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1311 = 8'h1d == _GEN_96 ? phv_data_29 : _GEN_1310; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1312 = 8'h1e == _GEN_96 ? phv_data_30 : _GEN_1311; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1313 = 8'h1f == _GEN_96 ? phv_data_31 : _GEN_1312; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1314 = 8'h20 == _GEN_96 ? phv_data_32 : _GEN_1313; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1315 = 8'h21 == _GEN_96 ? phv_data_33 : _GEN_1314; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1316 = 8'h22 == _GEN_96 ? phv_data_34 : _GEN_1315; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1317 = 8'h23 == _GEN_96 ? phv_data_35 : _GEN_1316; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1318 = 8'h24 == _GEN_96 ? phv_data_36 : _GEN_1317; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1319 = 8'h25 == _GEN_96 ? phv_data_37 : _GEN_1318; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1320 = 8'h26 == _GEN_96 ? phv_data_38 : _GEN_1319; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1321 = 8'h27 == _GEN_96 ? phv_data_39 : _GEN_1320; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1322 = 8'h28 == _GEN_96 ? phv_data_40 : _GEN_1321; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1323 = 8'h29 == _GEN_96 ? phv_data_41 : _GEN_1322; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1324 = 8'h2a == _GEN_96 ? phv_data_42 : _GEN_1323; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1325 = 8'h2b == _GEN_96 ? phv_data_43 : _GEN_1324; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1326 = 8'h2c == _GEN_96 ? phv_data_44 : _GEN_1325; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1327 = 8'h2d == _GEN_96 ? phv_data_45 : _GEN_1326; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1328 = 8'h2e == _GEN_96 ? phv_data_46 : _GEN_1327; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1329 = 8'h2f == _GEN_96 ? phv_data_47 : _GEN_1328; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1330 = 8'h30 == _GEN_96 ? phv_data_48 : _GEN_1329; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1331 = 8'h31 == _GEN_96 ? phv_data_49 : _GEN_1330; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1332 = 8'h32 == _GEN_96 ? phv_data_50 : _GEN_1331; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1333 = 8'h33 == _GEN_96 ? phv_data_51 : _GEN_1332; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1334 = 8'h34 == _GEN_96 ? phv_data_52 : _GEN_1333; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1335 = 8'h35 == _GEN_96 ? phv_data_53 : _GEN_1334; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1336 = 8'h36 == _GEN_96 ? phv_data_54 : _GEN_1335; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1337 = 8'h37 == _GEN_96 ? phv_data_55 : _GEN_1336; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1338 = 8'h38 == _GEN_96 ? phv_data_56 : _GEN_1337; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1339 = 8'h39 == _GEN_96 ? phv_data_57 : _GEN_1338; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1340 = 8'h3a == _GEN_96 ? phv_data_58 : _GEN_1339; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1341 = 8'h3b == _GEN_96 ? phv_data_59 : _GEN_1340; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1342 = 8'h3c == _GEN_96 ? phv_data_60 : _GEN_1341; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1343 = 8'h3d == _GEN_96 ? phv_data_61 : _GEN_1342; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1344 = 8'h3e == _GEN_96 ? phv_data_62 : _GEN_1343; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1345 = 8'h3f == _GEN_96 ? phv_data_63 : _GEN_1344; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] bytes_2_2 = _GEN_72 ? _GEN_1345 : 8'h0; // @[matcher_pisa.scala 129:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_1347 = 8'h0 == _GEN_97 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_1348 = 8'h1 == _GEN_97 ? phv_data_1 : _GEN_1347; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1349 = 8'h2 == _GEN_97 ? phv_data_2 : _GEN_1348; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1350 = 8'h3 == _GEN_97 ? phv_data_3 : _GEN_1349; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1351 = 8'h4 == _GEN_97 ? phv_data_4 : _GEN_1350; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1352 = 8'h5 == _GEN_97 ? phv_data_5 : _GEN_1351; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1353 = 8'h6 == _GEN_97 ? phv_data_6 : _GEN_1352; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1354 = 8'h7 == _GEN_97 ? phv_data_7 : _GEN_1353; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1355 = 8'h8 == _GEN_97 ? phv_data_8 : _GEN_1354; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1356 = 8'h9 == _GEN_97 ? phv_data_9 : _GEN_1355; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1357 = 8'ha == _GEN_97 ? phv_data_10 : _GEN_1356; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1358 = 8'hb == _GEN_97 ? phv_data_11 : _GEN_1357; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1359 = 8'hc == _GEN_97 ? phv_data_12 : _GEN_1358; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1360 = 8'hd == _GEN_97 ? phv_data_13 : _GEN_1359; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1361 = 8'he == _GEN_97 ? phv_data_14 : _GEN_1360; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1362 = 8'hf == _GEN_97 ? phv_data_15 : _GEN_1361; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1363 = 8'h10 == _GEN_97 ? phv_data_16 : _GEN_1362; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1364 = 8'h11 == _GEN_97 ? phv_data_17 : _GEN_1363; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1365 = 8'h12 == _GEN_97 ? phv_data_18 : _GEN_1364; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1366 = 8'h13 == _GEN_97 ? phv_data_19 : _GEN_1365; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1367 = 8'h14 == _GEN_97 ? phv_data_20 : _GEN_1366; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1368 = 8'h15 == _GEN_97 ? phv_data_21 : _GEN_1367; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1369 = 8'h16 == _GEN_97 ? phv_data_22 : _GEN_1368; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1370 = 8'h17 == _GEN_97 ? phv_data_23 : _GEN_1369; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1371 = 8'h18 == _GEN_97 ? phv_data_24 : _GEN_1370; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1372 = 8'h19 == _GEN_97 ? phv_data_25 : _GEN_1371; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1373 = 8'h1a == _GEN_97 ? phv_data_26 : _GEN_1372; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1374 = 8'h1b == _GEN_97 ? phv_data_27 : _GEN_1373; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1375 = 8'h1c == _GEN_97 ? phv_data_28 : _GEN_1374; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1376 = 8'h1d == _GEN_97 ? phv_data_29 : _GEN_1375; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1377 = 8'h1e == _GEN_97 ? phv_data_30 : _GEN_1376; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1378 = 8'h1f == _GEN_97 ? phv_data_31 : _GEN_1377; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1379 = 8'h20 == _GEN_97 ? phv_data_32 : _GEN_1378; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1380 = 8'h21 == _GEN_97 ? phv_data_33 : _GEN_1379; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1381 = 8'h22 == _GEN_97 ? phv_data_34 : _GEN_1380; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1382 = 8'h23 == _GEN_97 ? phv_data_35 : _GEN_1381; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1383 = 8'h24 == _GEN_97 ? phv_data_36 : _GEN_1382; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1384 = 8'h25 == _GEN_97 ? phv_data_37 : _GEN_1383; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1385 = 8'h26 == _GEN_97 ? phv_data_38 : _GEN_1384; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1386 = 8'h27 == _GEN_97 ? phv_data_39 : _GEN_1385; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1387 = 8'h28 == _GEN_97 ? phv_data_40 : _GEN_1386; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1388 = 8'h29 == _GEN_97 ? phv_data_41 : _GEN_1387; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1389 = 8'h2a == _GEN_97 ? phv_data_42 : _GEN_1388; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1390 = 8'h2b == _GEN_97 ? phv_data_43 : _GEN_1389; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1391 = 8'h2c == _GEN_97 ? phv_data_44 : _GEN_1390; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1392 = 8'h2d == _GEN_97 ? phv_data_45 : _GEN_1391; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1393 = 8'h2e == _GEN_97 ? phv_data_46 : _GEN_1392; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1394 = 8'h2f == _GEN_97 ? phv_data_47 : _GEN_1393; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1395 = 8'h30 == _GEN_97 ? phv_data_48 : _GEN_1394; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1396 = 8'h31 == _GEN_97 ? phv_data_49 : _GEN_1395; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1397 = 8'h32 == _GEN_97 ? phv_data_50 : _GEN_1396; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1398 = 8'h33 == _GEN_97 ? phv_data_51 : _GEN_1397; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1399 = 8'h34 == _GEN_97 ? phv_data_52 : _GEN_1398; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1400 = 8'h35 == _GEN_97 ? phv_data_53 : _GEN_1399; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1401 = 8'h36 == _GEN_97 ? phv_data_54 : _GEN_1400; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1402 = 8'h37 == _GEN_97 ? phv_data_55 : _GEN_1401; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1403 = 8'h38 == _GEN_97 ? phv_data_56 : _GEN_1402; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1404 = 8'h39 == _GEN_97 ? phv_data_57 : _GEN_1403; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1405 = 8'h3a == _GEN_97 ? phv_data_58 : _GEN_1404; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1406 = 8'h3b == _GEN_97 ? phv_data_59 : _GEN_1405; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1407 = 8'h3c == _GEN_97 ? phv_data_60 : _GEN_1406; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1408 = 8'h3d == _GEN_97 ? phv_data_61 : _GEN_1407; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1409 = 8'h3e == _GEN_97 ? phv_data_62 : _GEN_1408; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1410 = 8'h3f == _GEN_97 ? phv_data_63 : _GEN_1409; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] bytes_2_3 = _GEN_73 ? _GEN_1410 : 8'h0; // @[matcher_pisa.scala 129:46 matcher_pisa.scala 128:34]
  wire [31:0] _groups_2_T = {bytes_2_0,bytes_2_1,bytes_2_2,bytes_2_3}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_1412 = _GEN_58 == 2'h1 ? _groups_2_T : 32'h0; // @[matcher_pisa.scala 123:50 matcher_pisa.scala 137:31 matcher_pisa.scala 122:27]
  wire [15:0] _GEN_1413 = 8'h40 == _GEN_94 ? _double_bytes_0_T : 16'h0; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53 matcher_pisa.scala 144:41]
  wire [15:0] _GEN_1414 = 8'h41 == _GEN_94 ? _double_bytes_0_T_1 : _GEN_1413; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1415 = 8'h42 == _GEN_94 ? _double_bytes_0_T_2 : _GEN_1414; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1416 = 8'h43 == _GEN_94 ? _double_bytes_0_T_3 : _GEN_1415; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1417 = 8'h44 == _GEN_94 ? _double_bytes_0_T_4 : _GEN_1416; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1418 = 8'h45 == _GEN_94 ? _double_bytes_0_T_5 : _GEN_1417; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1419 = 8'h46 == _GEN_94 ? _double_bytes_0_T_6 : _GEN_1418; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1420 = 8'h47 == _GEN_94 ? _double_bytes_0_T_7 : _GEN_1419; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1421 = 8'h48 == _GEN_94 ? _double_bytes_0_T_8 : _GEN_1420; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1422 = 8'h49 == _GEN_94 ? _double_bytes_0_T_9 : _GEN_1421; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1423 = 8'h4a == _GEN_94 ? _double_bytes_0_T_10 : _GEN_1422; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1424 = 8'h4b == _GEN_94 ? _double_bytes_0_T_11 : _GEN_1423; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1425 = 8'h4c == _GEN_94 ? _double_bytes_0_T_12 : _GEN_1424; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1426 = 8'h4d == _GEN_94 ? _double_bytes_0_T_13 : _GEN_1425; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1427 = 8'h4e == _GEN_94 ? _double_bytes_0_T_14 : _GEN_1426; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1428 = 8'h4f == _GEN_94 ? _double_bytes_0_T_15 : _GEN_1427; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1429 = 8'h50 == _GEN_94 ? _double_bytes_0_T_16 : _GEN_1428; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1430 = 8'h51 == _GEN_94 ? _double_bytes_0_T_17 : _GEN_1429; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1431 = 8'h52 == _GEN_94 ? _double_bytes_0_T_18 : _GEN_1430; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1432 = 8'h53 == _GEN_94 ? _double_bytes_0_T_19 : _GEN_1431; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1433 = 8'h54 == _GEN_94 ? _double_bytes_0_T_20 : _GEN_1432; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1434 = 8'h55 == _GEN_94 ? _double_bytes_0_T_21 : _GEN_1433; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1435 = 8'h56 == _GEN_94 ? _double_bytes_0_T_22 : _GEN_1434; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1436 = 8'h57 == _GEN_94 ? _double_bytes_0_T_23 : _GEN_1435; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1437 = 8'h58 == _GEN_94 ? _double_bytes_0_T_24 : _GEN_1436; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1438 = 8'h59 == _GEN_94 ? _double_bytes_0_T_25 : _GEN_1437; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1439 = 8'h5a == _GEN_94 ? _double_bytes_0_T_26 : _GEN_1438; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1440 = 8'h5b == _GEN_94 ? _double_bytes_0_T_27 : _GEN_1439; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1441 = 8'h5c == _GEN_94 ? _double_bytes_0_T_28 : _GEN_1440; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1442 = 8'h5d == _GEN_94 ? _double_bytes_0_T_29 : _GEN_1441; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1443 = 8'h5e == _GEN_94 ? _double_bytes_0_T_30 : _GEN_1442; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1444 = 8'h5f == _GEN_94 ? _double_bytes_0_T_31 : _GEN_1443; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1445 = 8'h60 == _GEN_94 ? _double_bytes_0_T_32 : _GEN_1444; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1446 = 8'h61 == _GEN_94 ? _double_bytes_0_T_33 : _GEN_1445; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1447 = 8'h62 == _GEN_94 ? _double_bytes_0_T_34 : _GEN_1446; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1448 = 8'h63 == _GEN_94 ? _double_bytes_0_T_35 : _GEN_1447; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1449 = 8'h64 == _GEN_94 ? _double_bytes_0_T_36 : _GEN_1448; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1450 = 8'h65 == _GEN_94 ? _double_bytes_0_T_37 : _GEN_1449; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1451 = 8'h66 == _GEN_94 ? _double_bytes_0_T_38 : _GEN_1450; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1452 = 8'h67 == _GEN_94 ? _double_bytes_0_T_39 : _GEN_1451; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1453 = 8'h68 == _GEN_94 ? _double_bytes_0_T_40 : _GEN_1452; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1454 = 8'h69 == _GEN_94 ? _double_bytes_0_T_41 : _GEN_1453; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1455 = 8'h6a == _GEN_94 ? _double_bytes_0_T_42 : _GEN_1454; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1456 = 8'h6b == _GEN_94 ? _double_bytes_0_T_43 : _GEN_1455; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1457 = 8'h6c == _GEN_94 ? _double_bytes_0_T_44 : _GEN_1456; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1458 = 8'h6d == _GEN_94 ? _double_bytes_0_T_45 : _GEN_1457; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1459 = 8'h6e == _GEN_94 ? _double_bytes_0_T_46 : _GEN_1458; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1460 = 8'h6f == _GEN_94 ? _double_bytes_0_T_47 : _GEN_1459; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1461 = 8'h70 == _GEN_94 ? _double_bytes_0_T_48 : _GEN_1460; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1462 = 8'h71 == _GEN_94 ? _double_bytes_0_T_49 : _GEN_1461; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1463 = 8'h72 == _GEN_94 ? _double_bytes_0_T_50 : _GEN_1462; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1464 = 8'h73 == _GEN_94 ? _double_bytes_0_T_51 : _GEN_1463; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1465 = 8'h74 == _GEN_94 ? _double_bytes_0_T_52 : _GEN_1464; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1466 = 8'h75 == _GEN_94 ? _double_bytes_0_T_53 : _GEN_1465; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1467 = 8'h76 == _GEN_94 ? _double_bytes_0_T_54 : _GEN_1466; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1468 = 8'h77 == _GEN_94 ? _double_bytes_0_T_55 : _GEN_1467; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1469 = 8'h78 == _GEN_94 ? _double_bytes_0_T_56 : _GEN_1468; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1470 = 8'h79 == _GEN_94 ? _double_bytes_0_T_57 : _GEN_1469; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1471 = 8'h7a == _GEN_94 ? _double_bytes_0_T_58 : _GEN_1470; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1472 = 8'h7b == _GEN_94 ? _double_bytes_0_T_59 : _GEN_1471; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1473 = 8'h7c == _GEN_94 ? _double_bytes_0_T_60 : _GEN_1472; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1474 = 8'h7d == _GEN_94 ? _double_bytes_0_T_61 : _GEN_1473; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1475 = 8'h7e == _GEN_94 ? _double_bytes_0_T_62 : _GEN_1474; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1476 = 8'h7f == _GEN_94 ? _double_bytes_0_T_63 : _GEN_1475; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1477 = 8'h80 == _GEN_94 ? _double_bytes_0_T_64 : _GEN_1476; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1478 = 8'h81 == _GEN_94 ? _double_bytes_0_T_65 : _GEN_1477; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1479 = 8'h82 == _GEN_94 ? _double_bytes_0_T_66 : _GEN_1478; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1480 = 8'h83 == _GEN_94 ? _double_bytes_0_T_67 : _GEN_1479; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1481 = 8'h84 == _GEN_94 ? _double_bytes_0_T_68 : _GEN_1480; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1482 = 8'h85 == _GEN_94 ? _double_bytes_0_T_69 : _GEN_1481; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1483 = 8'h86 == _GEN_94 ? _double_bytes_0_T_70 : _GEN_1482; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1484 = 8'h87 == _GEN_94 ? _double_bytes_0_T_71 : _GEN_1483; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1485 = 8'h88 == _GEN_94 ? _double_bytes_0_T_72 : _GEN_1484; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1486 = 8'h89 == _GEN_94 ? _double_bytes_0_T_73 : _GEN_1485; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1487 = 8'h8a == _GEN_94 ? _double_bytes_0_T_74 : _GEN_1486; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1488 = 8'h8b == _GEN_94 ? _double_bytes_0_T_75 : _GEN_1487; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1489 = 8'h8c == _GEN_94 ? _double_bytes_0_T_76 : _GEN_1488; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1490 = 8'h8d == _GEN_94 ? _double_bytes_0_T_77 : _GEN_1489; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1491 = 8'h8e == _GEN_94 ? _double_bytes_0_T_78 : _GEN_1490; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1492 = 8'h8f == _GEN_94 ? _double_bytes_0_T_79 : _GEN_1491; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1493 = 8'h90 == _GEN_94 ? _double_bytes_0_T_80 : _GEN_1492; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1494 = 8'h91 == _GEN_94 ? _double_bytes_0_T_81 : _GEN_1493; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1495 = 8'h92 == _GEN_94 ? _double_bytes_0_T_82 : _GEN_1494; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1496 = 8'h93 == _GEN_94 ? _double_bytes_0_T_83 : _GEN_1495; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1497 = 8'h94 == _GEN_94 ? _double_bytes_0_T_84 : _GEN_1496; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1498 = 8'h95 == _GEN_94 ? _double_bytes_0_T_85 : _GEN_1497; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1499 = 8'h96 == _GEN_94 ? _double_bytes_0_T_86 : _GEN_1498; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1500 = 8'h97 == _GEN_94 ? _double_bytes_0_T_87 : _GEN_1499; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1501 = 8'h98 == _GEN_94 ? _double_bytes_0_T_88 : _GEN_1500; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1502 = 8'h99 == _GEN_94 ? _double_bytes_0_T_89 : _GEN_1501; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1503 = 8'h9a == _GEN_94 ? _double_bytes_0_T_90 : _GEN_1502; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1504 = 8'h9b == _GEN_94 ? _double_bytes_0_T_91 : _GEN_1503; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1505 = 8'h9c == _GEN_94 ? _double_bytes_0_T_92 : _GEN_1504; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1506 = 8'h9d == _GEN_94 ? _double_bytes_0_T_93 : _GEN_1505; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1507 = 8'h9e == _GEN_94 ? _double_bytes_0_T_94 : _GEN_1506; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1508 = 8'h9f == _GEN_94 ? _double_bytes_0_T_95 : _GEN_1507; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] double_bytes_2_0 = _GEN_70 ? _GEN_1508 : 16'h0; // @[matcher_pisa.scala 145:46 matcher_pisa.scala 144:41]
  wire [15:0] _GEN_1510 = 8'h40 == _GEN_95 ? _double_bytes_0_T : 16'h0; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53 matcher_pisa.scala 144:41]
  wire [15:0] _GEN_1511 = 8'h41 == _GEN_95 ? _double_bytes_0_T_1 : _GEN_1510; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1512 = 8'h42 == _GEN_95 ? _double_bytes_0_T_2 : _GEN_1511; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1513 = 8'h43 == _GEN_95 ? _double_bytes_0_T_3 : _GEN_1512; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1514 = 8'h44 == _GEN_95 ? _double_bytes_0_T_4 : _GEN_1513; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1515 = 8'h45 == _GEN_95 ? _double_bytes_0_T_5 : _GEN_1514; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1516 = 8'h46 == _GEN_95 ? _double_bytes_0_T_6 : _GEN_1515; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1517 = 8'h47 == _GEN_95 ? _double_bytes_0_T_7 : _GEN_1516; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1518 = 8'h48 == _GEN_95 ? _double_bytes_0_T_8 : _GEN_1517; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1519 = 8'h49 == _GEN_95 ? _double_bytes_0_T_9 : _GEN_1518; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1520 = 8'h4a == _GEN_95 ? _double_bytes_0_T_10 : _GEN_1519; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1521 = 8'h4b == _GEN_95 ? _double_bytes_0_T_11 : _GEN_1520; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1522 = 8'h4c == _GEN_95 ? _double_bytes_0_T_12 : _GEN_1521; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1523 = 8'h4d == _GEN_95 ? _double_bytes_0_T_13 : _GEN_1522; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1524 = 8'h4e == _GEN_95 ? _double_bytes_0_T_14 : _GEN_1523; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1525 = 8'h4f == _GEN_95 ? _double_bytes_0_T_15 : _GEN_1524; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1526 = 8'h50 == _GEN_95 ? _double_bytes_0_T_16 : _GEN_1525; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1527 = 8'h51 == _GEN_95 ? _double_bytes_0_T_17 : _GEN_1526; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1528 = 8'h52 == _GEN_95 ? _double_bytes_0_T_18 : _GEN_1527; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1529 = 8'h53 == _GEN_95 ? _double_bytes_0_T_19 : _GEN_1528; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1530 = 8'h54 == _GEN_95 ? _double_bytes_0_T_20 : _GEN_1529; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1531 = 8'h55 == _GEN_95 ? _double_bytes_0_T_21 : _GEN_1530; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1532 = 8'h56 == _GEN_95 ? _double_bytes_0_T_22 : _GEN_1531; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1533 = 8'h57 == _GEN_95 ? _double_bytes_0_T_23 : _GEN_1532; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1534 = 8'h58 == _GEN_95 ? _double_bytes_0_T_24 : _GEN_1533; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1535 = 8'h59 == _GEN_95 ? _double_bytes_0_T_25 : _GEN_1534; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1536 = 8'h5a == _GEN_95 ? _double_bytes_0_T_26 : _GEN_1535; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1537 = 8'h5b == _GEN_95 ? _double_bytes_0_T_27 : _GEN_1536; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1538 = 8'h5c == _GEN_95 ? _double_bytes_0_T_28 : _GEN_1537; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1539 = 8'h5d == _GEN_95 ? _double_bytes_0_T_29 : _GEN_1538; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1540 = 8'h5e == _GEN_95 ? _double_bytes_0_T_30 : _GEN_1539; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1541 = 8'h5f == _GEN_95 ? _double_bytes_0_T_31 : _GEN_1540; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1542 = 8'h60 == _GEN_95 ? _double_bytes_0_T_32 : _GEN_1541; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1543 = 8'h61 == _GEN_95 ? _double_bytes_0_T_33 : _GEN_1542; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1544 = 8'h62 == _GEN_95 ? _double_bytes_0_T_34 : _GEN_1543; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1545 = 8'h63 == _GEN_95 ? _double_bytes_0_T_35 : _GEN_1544; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1546 = 8'h64 == _GEN_95 ? _double_bytes_0_T_36 : _GEN_1545; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1547 = 8'h65 == _GEN_95 ? _double_bytes_0_T_37 : _GEN_1546; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1548 = 8'h66 == _GEN_95 ? _double_bytes_0_T_38 : _GEN_1547; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1549 = 8'h67 == _GEN_95 ? _double_bytes_0_T_39 : _GEN_1548; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1550 = 8'h68 == _GEN_95 ? _double_bytes_0_T_40 : _GEN_1549; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1551 = 8'h69 == _GEN_95 ? _double_bytes_0_T_41 : _GEN_1550; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1552 = 8'h6a == _GEN_95 ? _double_bytes_0_T_42 : _GEN_1551; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1553 = 8'h6b == _GEN_95 ? _double_bytes_0_T_43 : _GEN_1552; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1554 = 8'h6c == _GEN_95 ? _double_bytes_0_T_44 : _GEN_1553; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1555 = 8'h6d == _GEN_95 ? _double_bytes_0_T_45 : _GEN_1554; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1556 = 8'h6e == _GEN_95 ? _double_bytes_0_T_46 : _GEN_1555; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1557 = 8'h6f == _GEN_95 ? _double_bytes_0_T_47 : _GEN_1556; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1558 = 8'h70 == _GEN_95 ? _double_bytes_0_T_48 : _GEN_1557; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1559 = 8'h71 == _GEN_95 ? _double_bytes_0_T_49 : _GEN_1558; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1560 = 8'h72 == _GEN_95 ? _double_bytes_0_T_50 : _GEN_1559; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1561 = 8'h73 == _GEN_95 ? _double_bytes_0_T_51 : _GEN_1560; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1562 = 8'h74 == _GEN_95 ? _double_bytes_0_T_52 : _GEN_1561; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1563 = 8'h75 == _GEN_95 ? _double_bytes_0_T_53 : _GEN_1562; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1564 = 8'h76 == _GEN_95 ? _double_bytes_0_T_54 : _GEN_1563; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1565 = 8'h77 == _GEN_95 ? _double_bytes_0_T_55 : _GEN_1564; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1566 = 8'h78 == _GEN_95 ? _double_bytes_0_T_56 : _GEN_1565; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1567 = 8'h79 == _GEN_95 ? _double_bytes_0_T_57 : _GEN_1566; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1568 = 8'h7a == _GEN_95 ? _double_bytes_0_T_58 : _GEN_1567; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1569 = 8'h7b == _GEN_95 ? _double_bytes_0_T_59 : _GEN_1568; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1570 = 8'h7c == _GEN_95 ? _double_bytes_0_T_60 : _GEN_1569; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1571 = 8'h7d == _GEN_95 ? _double_bytes_0_T_61 : _GEN_1570; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1572 = 8'h7e == _GEN_95 ? _double_bytes_0_T_62 : _GEN_1571; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1573 = 8'h7f == _GEN_95 ? _double_bytes_0_T_63 : _GEN_1572; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1574 = 8'h80 == _GEN_95 ? _double_bytes_0_T_64 : _GEN_1573; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1575 = 8'h81 == _GEN_95 ? _double_bytes_0_T_65 : _GEN_1574; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1576 = 8'h82 == _GEN_95 ? _double_bytes_0_T_66 : _GEN_1575; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1577 = 8'h83 == _GEN_95 ? _double_bytes_0_T_67 : _GEN_1576; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1578 = 8'h84 == _GEN_95 ? _double_bytes_0_T_68 : _GEN_1577; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1579 = 8'h85 == _GEN_95 ? _double_bytes_0_T_69 : _GEN_1578; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1580 = 8'h86 == _GEN_95 ? _double_bytes_0_T_70 : _GEN_1579; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1581 = 8'h87 == _GEN_95 ? _double_bytes_0_T_71 : _GEN_1580; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1582 = 8'h88 == _GEN_95 ? _double_bytes_0_T_72 : _GEN_1581; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1583 = 8'h89 == _GEN_95 ? _double_bytes_0_T_73 : _GEN_1582; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1584 = 8'h8a == _GEN_95 ? _double_bytes_0_T_74 : _GEN_1583; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1585 = 8'h8b == _GEN_95 ? _double_bytes_0_T_75 : _GEN_1584; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1586 = 8'h8c == _GEN_95 ? _double_bytes_0_T_76 : _GEN_1585; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1587 = 8'h8d == _GEN_95 ? _double_bytes_0_T_77 : _GEN_1586; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1588 = 8'h8e == _GEN_95 ? _double_bytes_0_T_78 : _GEN_1587; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1589 = 8'h8f == _GEN_95 ? _double_bytes_0_T_79 : _GEN_1588; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1590 = 8'h90 == _GEN_95 ? _double_bytes_0_T_80 : _GEN_1589; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1591 = 8'h91 == _GEN_95 ? _double_bytes_0_T_81 : _GEN_1590; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1592 = 8'h92 == _GEN_95 ? _double_bytes_0_T_82 : _GEN_1591; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1593 = 8'h93 == _GEN_95 ? _double_bytes_0_T_83 : _GEN_1592; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1594 = 8'h94 == _GEN_95 ? _double_bytes_0_T_84 : _GEN_1593; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1595 = 8'h95 == _GEN_95 ? _double_bytes_0_T_85 : _GEN_1594; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1596 = 8'h96 == _GEN_95 ? _double_bytes_0_T_86 : _GEN_1595; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1597 = 8'h97 == _GEN_95 ? _double_bytes_0_T_87 : _GEN_1596; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1598 = 8'h98 == _GEN_95 ? _double_bytes_0_T_88 : _GEN_1597; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1599 = 8'h99 == _GEN_95 ? _double_bytes_0_T_89 : _GEN_1598; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1600 = 8'h9a == _GEN_95 ? _double_bytes_0_T_90 : _GEN_1599; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1601 = 8'h9b == _GEN_95 ? _double_bytes_0_T_91 : _GEN_1600; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1602 = 8'h9c == _GEN_95 ? _double_bytes_0_T_92 : _GEN_1601; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1603 = 8'h9d == _GEN_95 ? _double_bytes_0_T_93 : _GEN_1602; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1604 = 8'h9e == _GEN_95 ? _double_bytes_0_T_94 : _GEN_1603; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1605 = 8'h9f == _GEN_95 ? _double_bytes_0_T_95 : _GEN_1604; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] double_bytes_2_1 = _GEN_71 ? _GEN_1605 : 16'h0; // @[matcher_pisa.scala 145:46 matcher_pisa.scala 144:41]
  wire [31:0] _groups_2_T_1 = {double_bytes_2_0,double_bytes_2_1}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_1607 = _GEN_58 == 2'h2 ? _groups_2_T_1 : _GEN_1412; // @[matcher_pisa.scala 139:50 matcher_pisa.scala 153:31]
  wire [31:0] _GEN_1608 = 8'ha0 == _GEN_94 ? _groups_0_T_2 : 32'h0; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39 matcher_pisa.scala 158:31]
  wire [31:0] _GEN_1609 = 8'ha1 == _GEN_94 ? _groups_0_T_3 : _GEN_1608; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1610 = 8'ha2 == _GEN_94 ? _groups_0_T_4 : _GEN_1609; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1611 = 8'ha3 == _GEN_94 ? _groups_0_T_5 : _GEN_1610; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1612 = 8'ha4 == _GEN_94 ? _groups_0_T_6 : _GEN_1611; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1613 = 8'ha5 == _GEN_94 ? _groups_0_T_7 : _GEN_1612; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1614 = 8'ha6 == _GEN_94 ? _groups_0_T_8 : _GEN_1613; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1615 = 8'ha7 == _GEN_94 ? _groups_0_T_9 : _GEN_1614; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1616 = 8'ha8 == _GEN_94 ? _groups_0_T_10 : _GEN_1615; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1617 = 8'ha9 == _GEN_94 ? _groups_0_T_11 : _GEN_1616; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1618 = 8'haa == _GEN_94 ? _groups_0_T_12 : _GEN_1617; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1619 = 8'hab == _GEN_94 ? _groups_0_T_13 : _GEN_1618; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1620 = 8'hac == _GEN_94 ? _groups_0_T_14 : _GEN_1619; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1621 = 8'had == _GEN_94 ? _groups_0_T_15 : _GEN_1620; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1622 = 8'hae == _GEN_94 ? _groups_0_T_16 : _GEN_1621; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1623 = 8'haf == _GEN_94 ? _groups_0_T_17 : _GEN_1622; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1624 = 8'hb0 == _GEN_94 ? _groups_0_T_18 : _GEN_1623; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1625 = 8'hb1 == _GEN_94 ? _groups_0_T_19 : _GEN_1624; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1626 = 8'hb2 == _GEN_94 ? _groups_0_T_20 : _GEN_1625; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1627 = 8'hb3 == _GEN_94 ? _groups_0_T_21 : _GEN_1626; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1628 = 8'hb4 == _GEN_94 ? _groups_0_T_22 : _GEN_1627; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1629 = 8'hb5 == _GEN_94 ? _groups_0_T_23 : _GEN_1628; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1630 = 8'hb6 == _GEN_94 ? _groups_0_T_24 : _GEN_1629; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1631 = 8'hb7 == _GEN_94 ? _groups_0_T_25 : _GEN_1630; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1632 = 8'hb8 == _GEN_94 ? _groups_0_T_26 : _GEN_1631; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1633 = 8'hb9 == _GEN_94 ? _groups_0_T_27 : _GEN_1632; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1634 = 8'hba == _GEN_94 ? _groups_0_T_28 : _GEN_1633; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1635 = 8'hbb == _GEN_94 ? _groups_0_T_29 : _GEN_1634; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1636 = 8'hbc == _GEN_94 ? _groups_0_T_30 : _GEN_1635; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1637 = 8'hbd == _GEN_94 ? _groups_0_T_31 : _GEN_1636; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1638 = 8'hbe == _GEN_94 ? _groups_0_T_32 : _GEN_1637; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1639 = 8'hbf == _GEN_94 ? _groups_0_T_33 : _GEN_1638; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1640 = 8'hc0 == _GEN_94 ? _groups_0_T_34 : _GEN_1639; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1641 = 8'hc1 == _GEN_94 ? _groups_0_T_35 : _GEN_1640; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1642 = 8'hc2 == _GEN_94 ? _groups_0_T_36 : _GEN_1641; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1643 = 8'hc3 == _GEN_94 ? _groups_0_T_37 : _GEN_1642; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1644 = 8'hc4 == _GEN_94 ? _groups_0_T_38 : _GEN_1643; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1645 = 8'hc5 == _GEN_94 ? _groups_0_T_39 : _GEN_1644; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1646 = 8'hc6 == _GEN_94 ? _groups_0_T_40 : _GEN_1645; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1647 = 8'hc7 == _GEN_94 ? _groups_0_T_41 : _GEN_1646; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1648 = 8'hc8 == _GEN_94 ? _groups_0_T_42 : _GEN_1647; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1649 = 8'hc9 == _GEN_94 ? _groups_0_T_43 : _GEN_1648; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1650 = 8'hca == _GEN_94 ? _groups_0_T_44 : _GEN_1649; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1651 = 8'hcb == _GEN_94 ? _groups_0_T_45 : _GEN_1650; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1652 = 8'hcc == _GEN_94 ? _groups_0_T_46 : _GEN_1651; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1653 = 8'hcd == _GEN_94 ? _groups_0_T_47 : _GEN_1652; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1654 = 8'hce == _GEN_94 ? _groups_0_T_48 : _GEN_1653; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1655 = 8'hcf == _GEN_94 ? _groups_0_T_49 : _GEN_1654; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1656 = 8'hd0 == _GEN_94 ? _groups_0_T_50 : _GEN_1655; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1657 = 8'hd1 == _GEN_94 ? _groups_0_T_51 : _GEN_1656; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1658 = 8'hd2 == _GEN_94 ? _groups_0_T_52 : _GEN_1657; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1659 = 8'hd3 == _GEN_94 ? _groups_0_T_53 : _GEN_1658; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1660 = 8'hd4 == _GEN_94 ? _groups_0_T_54 : _GEN_1659; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1661 = 8'hd5 == _GEN_94 ? _groups_0_T_55 : _GEN_1660; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1662 = 8'hd6 == _GEN_94 ? _groups_0_T_56 : _GEN_1661; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1663 = 8'hd7 == _GEN_94 ? _groups_0_T_57 : _GEN_1662; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1664 = 8'hd8 == _GEN_94 ? _groups_0_T_58 : _GEN_1663; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1665 = 8'hd9 == _GEN_94 ? _groups_0_T_59 : _GEN_1664; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1666 = 8'hda == _GEN_94 ? _groups_0_T_60 : _GEN_1665; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1667 = 8'hdb == _GEN_94 ? _groups_0_T_61 : _GEN_1666; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1668 = 8'hdc == _GEN_94 ? _groups_0_T_62 : _GEN_1667; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1669 = 8'hdd == _GEN_94 ? _groups_0_T_63 : _GEN_1668; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1670 = 8'hde == _GEN_94 ? _groups_0_T_64 : _GEN_1669; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1671 = 8'hdf == _GEN_94 ? _groups_0_T_65 : _GEN_1670; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] groups_2 = _GEN_58 == 2'h3 ? _GEN_1671 : _GEN_1607; // @[matcher_pisa.scala 155:50]
  wire [7:0] _GEN_1673 = 8'h0 == _GEN_98 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_1674 = 8'h1 == _GEN_98 ? phv_data_1 : _GEN_1673; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1675 = 8'h2 == _GEN_98 ? phv_data_2 : _GEN_1674; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1676 = 8'h3 == _GEN_98 ? phv_data_3 : _GEN_1675; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1677 = 8'h4 == _GEN_98 ? phv_data_4 : _GEN_1676; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1678 = 8'h5 == _GEN_98 ? phv_data_5 : _GEN_1677; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1679 = 8'h6 == _GEN_98 ? phv_data_6 : _GEN_1678; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1680 = 8'h7 == _GEN_98 ? phv_data_7 : _GEN_1679; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1681 = 8'h8 == _GEN_98 ? phv_data_8 : _GEN_1680; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1682 = 8'h9 == _GEN_98 ? phv_data_9 : _GEN_1681; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1683 = 8'ha == _GEN_98 ? phv_data_10 : _GEN_1682; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1684 = 8'hb == _GEN_98 ? phv_data_11 : _GEN_1683; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1685 = 8'hc == _GEN_98 ? phv_data_12 : _GEN_1684; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1686 = 8'hd == _GEN_98 ? phv_data_13 : _GEN_1685; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1687 = 8'he == _GEN_98 ? phv_data_14 : _GEN_1686; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1688 = 8'hf == _GEN_98 ? phv_data_15 : _GEN_1687; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1689 = 8'h10 == _GEN_98 ? phv_data_16 : _GEN_1688; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1690 = 8'h11 == _GEN_98 ? phv_data_17 : _GEN_1689; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1691 = 8'h12 == _GEN_98 ? phv_data_18 : _GEN_1690; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1692 = 8'h13 == _GEN_98 ? phv_data_19 : _GEN_1691; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1693 = 8'h14 == _GEN_98 ? phv_data_20 : _GEN_1692; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1694 = 8'h15 == _GEN_98 ? phv_data_21 : _GEN_1693; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1695 = 8'h16 == _GEN_98 ? phv_data_22 : _GEN_1694; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1696 = 8'h17 == _GEN_98 ? phv_data_23 : _GEN_1695; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1697 = 8'h18 == _GEN_98 ? phv_data_24 : _GEN_1696; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1698 = 8'h19 == _GEN_98 ? phv_data_25 : _GEN_1697; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1699 = 8'h1a == _GEN_98 ? phv_data_26 : _GEN_1698; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1700 = 8'h1b == _GEN_98 ? phv_data_27 : _GEN_1699; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1701 = 8'h1c == _GEN_98 ? phv_data_28 : _GEN_1700; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1702 = 8'h1d == _GEN_98 ? phv_data_29 : _GEN_1701; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1703 = 8'h1e == _GEN_98 ? phv_data_30 : _GEN_1702; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1704 = 8'h1f == _GEN_98 ? phv_data_31 : _GEN_1703; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1705 = 8'h20 == _GEN_98 ? phv_data_32 : _GEN_1704; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1706 = 8'h21 == _GEN_98 ? phv_data_33 : _GEN_1705; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1707 = 8'h22 == _GEN_98 ? phv_data_34 : _GEN_1706; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1708 = 8'h23 == _GEN_98 ? phv_data_35 : _GEN_1707; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1709 = 8'h24 == _GEN_98 ? phv_data_36 : _GEN_1708; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1710 = 8'h25 == _GEN_98 ? phv_data_37 : _GEN_1709; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1711 = 8'h26 == _GEN_98 ? phv_data_38 : _GEN_1710; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1712 = 8'h27 == _GEN_98 ? phv_data_39 : _GEN_1711; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1713 = 8'h28 == _GEN_98 ? phv_data_40 : _GEN_1712; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1714 = 8'h29 == _GEN_98 ? phv_data_41 : _GEN_1713; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1715 = 8'h2a == _GEN_98 ? phv_data_42 : _GEN_1714; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1716 = 8'h2b == _GEN_98 ? phv_data_43 : _GEN_1715; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1717 = 8'h2c == _GEN_98 ? phv_data_44 : _GEN_1716; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1718 = 8'h2d == _GEN_98 ? phv_data_45 : _GEN_1717; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1719 = 8'h2e == _GEN_98 ? phv_data_46 : _GEN_1718; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1720 = 8'h2f == _GEN_98 ? phv_data_47 : _GEN_1719; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1721 = 8'h30 == _GEN_98 ? phv_data_48 : _GEN_1720; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1722 = 8'h31 == _GEN_98 ? phv_data_49 : _GEN_1721; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1723 = 8'h32 == _GEN_98 ? phv_data_50 : _GEN_1722; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1724 = 8'h33 == _GEN_98 ? phv_data_51 : _GEN_1723; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1725 = 8'h34 == _GEN_98 ? phv_data_52 : _GEN_1724; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1726 = 8'h35 == _GEN_98 ? phv_data_53 : _GEN_1725; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1727 = 8'h36 == _GEN_98 ? phv_data_54 : _GEN_1726; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1728 = 8'h37 == _GEN_98 ? phv_data_55 : _GEN_1727; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1729 = 8'h38 == _GEN_98 ? phv_data_56 : _GEN_1728; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1730 = 8'h39 == _GEN_98 ? phv_data_57 : _GEN_1729; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1731 = 8'h3a == _GEN_98 ? phv_data_58 : _GEN_1730; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1732 = 8'h3b == _GEN_98 ? phv_data_59 : _GEN_1731; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1733 = 8'h3c == _GEN_98 ? phv_data_60 : _GEN_1732; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1734 = 8'h3d == _GEN_98 ? phv_data_61 : _GEN_1733; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1735 = 8'h3e == _GEN_98 ? phv_data_62 : _GEN_1734; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1736 = 8'h3f == _GEN_98 ? phv_data_63 : _GEN_1735; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] bytes_3_0 = _GEN_74 ? _GEN_1736 : 8'h0; // @[matcher_pisa.scala 129:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_1738 = 8'h0 == _GEN_99 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_1739 = 8'h1 == _GEN_99 ? phv_data_1 : _GEN_1738; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1740 = 8'h2 == _GEN_99 ? phv_data_2 : _GEN_1739; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1741 = 8'h3 == _GEN_99 ? phv_data_3 : _GEN_1740; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1742 = 8'h4 == _GEN_99 ? phv_data_4 : _GEN_1741; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1743 = 8'h5 == _GEN_99 ? phv_data_5 : _GEN_1742; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1744 = 8'h6 == _GEN_99 ? phv_data_6 : _GEN_1743; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1745 = 8'h7 == _GEN_99 ? phv_data_7 : _GEN_1744; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1746 = 8'h8 == _GEN_99 ? phv_data_8 : _GEN_1745; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1747 = 8'h9 == _GEN_99 ? phv_data_9 : _GEN_1746; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1748 = 8'ha == _GEN_99 ? phv_data_10 : _GEN_1747; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1749 = 8'hb == _GEN_99 ? phv_data_11 : _GEN_1748; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1750 = 8'hc == _GEN_99 ? phv_data_12 : _GEN_1749; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1751 = 8'hd == _GEN_99 ? phv_data_13 : _GEN_1750; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1752 = 8'he == _GEN_99 ? phv_data_14 : _GEN_1751; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1753 = 8'hf == _GEN_99 ? phv_data_15 : _GEN_1752; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1754 = 8'h10 == _GEN_99 ? phv_data_16 : _GEN_1753; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1755 = 8'h11 == _GEN_99 ? phv_data_17 : _GEN_1754; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1756 = 8'h12 == _GEN_99 ? phv_data_18 : _GEN_1755; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1757 = 8'h13 == _GEN_99 ? phv_data_19 : _GEN_1756; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1758 = 8'h14 == _GEN_99 ? phv_data_20 : _GEN_1757; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1759 = 8'h15 == _GEN_99 ? phv_data_21 : _GEN_1758; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1760 = 8'h16 == _GEN_99 ? phv_data_22 : _GEN_1759; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1761 = 8'h17 == _GEN_99 ? phv_data_23 : _GEN_1760; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1762 = 8'h18 == _GEN_99 ? phv_data_24 : _GEN_1761; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1763 = 8'h19 == _GEN_99 ? phv_data_25 : _GEN_1762; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1764 = 8'h1a == _GEN_99 ? phv_data_26 : _GEN_1763; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1765 = 8'h1b == _GEN_99 ? phv_data_27 : _GEN_1764; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1766 = 8'h1c == _GEN_99 ? phv_data_28 : _GEN_1765; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1767 = 8'h1d == _GEN_99 ? phv_data_29 : _GEN_1766; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1768 = 8'h1e == _GEN_99 ? phv_data_30 : _GEN_1767; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1769 = 8'h1f == _GEN_99 ? phv_data_31 : _GEN_1768; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1770 = 8'h20 == _GEN_99 ? phv_data_32 : _GEN_1769; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1771 = 8'h21 == _GEN_99 ? phv_data_33 : _GEN_1770; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1772 = 8'h22 == _GEN_99 ? phv_data_34 : _GEN_1771; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1773 = 8'h23 == _GEN_99 ? phv_data_35 : _GEN_1772; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1774 = 8'h24 == _GEN_99 ? phv_data_36 : _GEN_1773; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1775 = 8'h25 == _GEN_99 ? phv_data_37 : _GEN_1774; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1776 = 8'h26 == _GEN_99 ? phv_data_38 : _GEN_1775; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1777 = 8'h27 == _GEN_99 ? phv_data_39 : _GEN_1776; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1778 = 8'h28 == _GEN_99 ? phv_data_40 : _GEN_1777; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1779 = 8'h29 == _GEN_99 ? phv_data_41 : _GEN_1778; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1780 = 8'h2a == _GEN_99 ? phv_data_42 : _GEN_1779; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1781 = 8'h2b == _GEN_99 ? phv_data_43 : _GEN_1780; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1782 = 8'h2c == _GEN_99 ? phv_data_44 : _GEN_1781; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1783 = 8'h2d == _GEN_99 ? phv_data_45 : _GEN_1782; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1784 = 8'h2e == _GEN_99 ? phv_data_46 : _GEN_1783; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1785 = 8'h2f == _GEN_99 ? phv_data_47 : _GEN_1784; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1786 = 8'h30 == _GEN_99 ? phv_data_48 : _GEN_1785; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1787 = 8'h31 == _GEN_99 ? phv_data_49 : _GEN_1786; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1788 = 8'h32 == _GEN_99 ? phv_data_50 : _GEN_1787; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1789 = 8'h33 == _GEN_99 ? phv_data_51 : _GEN_1788; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1790 = 8'h34 == _GEN_99 ? phv_data_52 : _GEN_1789; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1791 = 8'h35 == _GEN_99 ? phv_data_53 : _GEN_1790; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1792 = 8'h36 == _GEN_99 ? phv_data_54 : _GEN_1791; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1793 = 8'h37 == _GEN_99 ? phv_data_55 : _GEN_1792; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1794 = 8'h38 == _GEN_99 ? phv_data_56 : _GEN_1793; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1795 = 8'h39 == _GEN_99 ? phv_data_57 : _GEN_1794; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1796 = 8'h3a == _GEN_99 ? phv_data_58 : _GEN_1795; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1797 = 8'h3b == _GEN_99 ? phv_data_59 : _GEN_1796; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1798 = 8'h3c == _GEN_99 ? phv_data_60 : _GEN_1797; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1799 = 8'h3d == _GEN_99 ? phv_data_61 : _GEN_1798; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1800 = 8'h3e == _GEN_99 ? phv_data_62 : _GEN_1799; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1801 = 8'h3f == _GEN_99 ? phv_data_63 : _GEN_1800; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] bytes_3_1 = _GEN_75 ? _GEN_1801 : 8'h0; // @[matcher_pisa.scala 129:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_1803 = 8'h0 == _GEN_100 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_1804 = 8'h1 == _GEN_100 ? phv_data_1 : _GEN_1803; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1805 = 8'h2 == _GEN_100 ? phv_data_2 : _GEN_1804; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1806 = 8'h3 == _GEN_100 ? phv_data_3 : _GEN_1805; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1807 = 8'h4 == _GEN_100 ? phv_data_4 : _GEN_1806; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1808 = 8'h5 == _GEN_100 ? phv_data_5 : _GEN_1807; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1809 = 8'h6 == _GEN_100 ? phv_data_6 : _GEN_1808; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1810 = 8'h7 == _GEN_100 ? phv_data_7 : _GEN_1809; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1811 = 8'h8 == _GEN_100 ? phv_data_8 : _GEN_1810; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1812 = 8'h9 == _GEN_100 ? phv_data_9 : _GEN_1811; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1813 = 8'ha == _GEN_100 ? phv_data_10 : _GEN_1812; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1814 = 8'hb == _GEN_100 ? phv_data_11 : _GEN_1813; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1815 = 8'hc == _GEN_100 ? phv_data_12 : _GEN_1814; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1816 = 8'hd == _GEN_100 ? phv_data_13 : _GEN_1815; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1817 = 8'he == _GEN_100 ? phv_data_14 : _GEN_1816; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1818 = 8'hf == _GEN_100 ? phv_data_15 : _GEN_1817; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1819 = 8'h10 == _GEN_100 ? phv_data_16 : _GEN_1818; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1820 = 8'h11 == _GEN_100 ? phv_data_17 : _GEN_1819; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1821 = 8'h12 == _GEN_100 ? phv_data_18 : _GEN_1820; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1822 = 8'h13 == _GEN_100 ? phv_data_19 : _GEN_1821; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1823 = 8'h14 == _GEN_100 ? phv_data_20 : _GEN_1822; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1824 = 8'h15 == _GEN_100 ? phv_data_21 : _GEN_1823; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1825 = 8'h16 == _GEN_100 ? phv_data_22 : _GEN_1824; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1826 = 8'h17 == _GEN_100 ? phv_data_23 : _GEN_1825; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1827 = 8'h18 == _GEN_100 ? phv_data_24 : _GEN_1826; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1828 = 8'h19 == _GEN_100 ? phv_data_25 : _GEN_1827; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1829 = 8'h1a == _GEN_100 ? phv_data_26 : _GEN_1828; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1830 = 8'h1b == _GEN_100 ? phv_data_27 : _GEN_1829; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1831 = 8'h1c == _GEN_100 ? phv_data_28 : _GEN_1830; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1832 = 8'h1d == _GEN_100 ? phv_data_29 : _GEN_1831; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1833 = 8'h1e == _GEN_100 ? phv_data_30 : _GEN_1832; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1834 = 8'h1f == _GEN_100 ? phv_data_31 : _GEN_1833; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1835 = 8'h20 == _GEN_100 ? phv_data_32 : _GEN_1834; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1836 = 8'h21 == _GEN_100 ? phv_data_33 : _GEN_1835; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1837 = 8'h22 == _GEN_100 ? phv_data_34 : _GEN_1836; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1838 = 8'h23 == _GEN_100 ? phv_data_35 : _GEN_1837; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1839 = 8'h24 == _GEN_100 ? phv_data_36 : _GEN_1838; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1840 = 8'h25 == _GEN_100 ? phv_data_37 : _GEN_1839; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1841 = 8'h26 == _GEN_100 ? phv_data_38 : _GEN_1840; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1842 = 8'h27 == _GEN_100 ? phv_data_39 : _GEN_1841; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1843 = 8'h28 == _GEN_100 ? phv_data_40 : _GEN_1842; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1844 = 8'h29 == _GEN_100 ? phv_data_41 : _GEN_1843; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1845 = 8'h2a == _GEN_100 ? phv_data_42 : _GEN_1844; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1846 = 8'h2b == _GEN_100 ? phv_data_43 : _GEN_1845; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1847 = 8'h2c == _GEN_100 ? phv_data_44 : _GEN_1846; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1848 = 8'h2d == _GEN_100 ? phv_data_45 : _GEN_1847; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1849 = 8'h2e == _GEN_100 ? phv_data_46 : _GEN_1848; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1850 = 8'h2f == _GEN_100 ? phv_data_47 : _GEN_1849; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1851 = 8'h30 == _GEN_100 ? phv_data_48 : _GEN_1850; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1852 = 8'h31 == _GEN_100 ? phv_data_49 : _GEN_1851; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1853 = 8'h32 == _GEN_100 ? phv_data_50 : _GEN_1852; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1854 = 8'h33 == _GEN_100 ? phv_data_51 : _GEN_1853; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1855 = 8'h34 == _GEN_100 ? phv_data_52 : _GEN_1854; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1856 = 8'h35 == _GEN_100 ? phv_data_53 : _GEN_1855; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1857 = 8'h36 == _GEN_100 ? phv_data_54 : _GEN_1856; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1858 = 8'h37 == _GEN_100 ? phv_data_55 : _GEN_1857; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1859 = 8'h38 == _GEN_100 ? phv_data_56 : _GEN_1858; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1860 = 8'h39 == _GEN_100 ? phv_data_57 : _GEN_1859; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1861 = 8'h3a == _GEN_100 ? phv_data_58 : _GEN_1860; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1862 = 8'h3b == _GEN_100 ? phv_data_59 : _GEN_1861; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1863 = 8'h3c == _GEN_100 ? phv_data_60 : _GEN_1862; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1864 = 8'h3d == _GEN_100 ? phv_data_61 : _GEN_1863; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1865 = 8'h3e == _GEN_100 ? phv_data_62 : _GEN_1864; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1866 = 8'h3f == _GEN_100 ? phv_data_63 : _GEN_1865; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] bytes_3_2 = _GEN_76 ? _GEN_1866 : 8'h0; // @[matcher_pisa.scala 129:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_1868 = 8'h0 == _GEN_101 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_1869 = 8'h1 == _GEN_101 ? phv_data_1 : _GEN_1868; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1870 = 8'h2 == _GEN_101 ? phv_data_2 : _GEN_1869; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1871 = 8'h3 == _GEN_101 ? phv_data_3 : _GEN_1870; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1872 = 8'h4 == _GEN_101 ? phv_data_4 : _GEN_1871; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1873 = 8'h5 == _GEN_101 ? phv_data_5 : _GEN_1872; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1874 = 8'h6 == _GEN_101 ? phv_data_6 : _GEN_1873; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1875 = 8'h7 == _GEN_101 ? phv_data_7 : _GEN_1874; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1876 = 8'h8 == _GEN_101 ? phv_data_8 : _GEN_1875; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1877 = 8'h9 == _GEN_101 ? phv_data_9 : _GEN_1876; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1878 = 8'ha == _GEN_101 ? phv_data_10 : _GEN_1877; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1879 = 8'hb == _GEN_101 ? phv_data_11 : _GEN_1878; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1880 = 8'hc == _GEN_101 ? phv_data_12 : _GEN_1879; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1881 = 8'hd == _GEN_101 ? phv_data_13 : _GEN_1880; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1882 = 8'he == _GEN_101 ? phv_data_14 : _GEN_1881; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1883 = 8'hf == _GEN_101 ? phv_data_15 : _GEN_1882; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1884 = 8'h10 == _GEN_101 ? phv_data_16 : _GEN_1883; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1885 = 8'h11 == _GEN_101 ? phv_data_17 : _GEN_1884; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1886 = 8'h12 == _GEN_101 ? phv_data_18 : _GEN_1885; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1887 = 8'h13 == _GEN_101 ? phv_data_19 : _GEN_1886; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1888 = 8'h14 == _GEN_101 ? phv_data_20 : _GEN_1887; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1889 = 8'h15 == _GEN_101 ? phv_data_21 : _GEN_1888; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1890 = 8'h16 == _GEN_101 ? phv_data_22 : _GEN_1889; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1891 = 8'h17 == _GEN_101 ? phv_data_23 : _GEN_1890; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1892 = 8'h18 == _GEN_101 ? phv_data_24 : _GEN_1891; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1893 = 8'h19 == _GEN_101 ? phv_data_25 : _GEN_1892; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1894 = 8'h1a == _GEN_101 ? phv_data_26 : _GEN_1893; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1895 = 8'h1b == _GEN_101 ? phv_data_27 : _GEN_1894; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1896 = 8'h1c == _GEN_101 ? phv_data_28 : _GEN_1895; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1897 = 8'h1d == _GEN_101 ? phv_data_29 : _GEN_1896; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1898 = 8'h1e == _GEN_101 ? phv_data_30 : _GEN_1897; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1899 = 8'h1f == _GEN_101 ? phv_data_31 : _GEN_1898; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1900 = 8'h20 == _GEN_101 ? phv_data_32 : _GEN_1899; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1901 = 8'h21 == _GEN_101 ? phv_data_33 : _GEN_1900; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1902 = 8'h22 == _GEN_101 ? phv_data_34 : _GEN_1901; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1903 = 8'h23 == _GEN_101 ? phv_data_35 : _GEN_1902; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1904 = 8'h24 == _GEN_101 ? phv_data_36 : _GEN_1903; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1905 = 8'h25 == _GEN_101 ? phv_data_37 : _GEN_1904; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1906 = 8'h26 == _GEN_101 ? phv_data_38 : _GEN_1905; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1907 = 8'h27 == _GEN_101 ? phv_data_39 : _GEN_1906; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1908 = 8'h28 == _GEN_101 ? phv_data_40 : _GEN_1907; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1909 = 8'h29 == _GEN_101 ? phv_data_41 : _GEN_1908; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1910 = 8'h2a == _GEN_101 ? phv_data_42 : _GEN_1909; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1911 = 8'h2b == _GEN_101 ? phv_data_43 : _GEN_1910; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1912 = 8'h2c == _GEN_101 ? phv_data_44 : _GEN_1911; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1913 = 8'h2d == _GEN_101 ? phv_data_45 : _GEN_1912; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1914 = 8'h2e == _GEN_101 ? phv_data_46 : _GEN_1913; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1915 = 8'h2f == _GEN_101 ? phv_data_47 : _GEN_1914; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1916 = 8'h30 == _GEN_101 ? phv_data_48 : _GEN_1915; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1917 = 8'h31 == _GEN_101 ? phv_data_49 : _GEN_1916; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1918 = 8'h32 == _GEN_101 ? phv_data_50 : _GEN_1917; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1919 = 8'h33 == _GEN_101 ? phv_data_51 : _GEN_1918; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1920 = 8'h34 == _GEN_101 ? phv_data_52 : _GEN_1919; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1921 = 8'h35 == _GEN_101 ? phv_data_53 : _GEN_1920; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1922 = 8'h36 == _GEN_101 ? phv_data_54 : _GEN_1921; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1923 = 8'h37 == _GEN_101 ? phv_data_55 : _GEN_1922; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1924 = 8'h38 == _GEN_101 ? phv_data_56 : _GEN_1923; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1925 = 8'h39 == _GEN_101 ? phv_data_57 : _GEN_1924; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1926 = 8'h3a == _GEN_101 ? phv_data_58 : _GEN_1925; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1927 = 8'h3b == _GEN_101 ? phv_data_59 : _GEN_1926; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1928 = 8'h3c == _GEN_101 ? phv_data_60 : _GEN_1927; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1929 = 8'h3d == _GEN_101 ? phv_data_61 : _GEN_1928; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1930 = 8'h3e == _GEN_101 ? phv_data_62 : _GEN_1929; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1931 = 8'h3f == _GEN_101 ? phv_data_63 : _GEN_1930; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] bytes_3_3 = _GEN_77 ? _GEN_1931 : 8'h0; // @[matcher_pisa.scala 129:46 matcher_pisa.scala 128:34]
  wire [31:0] _groups_3_T = {bytes_3_0,bytes_3_1,bytes_3_2,bytes_3_3}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_1933 = _GEN_59 == 2'h1 ? _groups_3_T : 32'h0; // @[matcher_pisa.scala 123:50 matcher_pisa.scala 137:31 matcher_pisa.scala 122:27]
  wire [15:0] _GEN_1934 = 8'h40 == _GEN_98 ? _double_bytes_0_T : 16'h0; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53 matcher_pisa.scala 144:41]
  wire [15:0] _GEN_1935 = 8'h41 == _GEN_98 ? _double_bytes_0_T_1 : _GEN_1934; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1936 = 8'h42 == _GEN_98 ? _double_bytes_0_T_2 : _GEN_1935; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1937 = 8'h43 == _GEN_98 ? _double_bytes_0_T_3 : _GEN_1936; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1938 = 8'h44 == _GEN_98 ? _double_bytes_0_T_4 : _GEN_1937; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1939 = 8'h45 == _GEN_98 ? _double_bytes_0_T_5 : _GEN_1938; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1940 = 8'h46 == _GEN_98 ? _double_bytes_0_T_6 : _GEN_1939; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1941 = 8'h47 == _GEN_98 ? _double_bytes_0_T_7 : _GEN_1940; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1942 = 8'h48 == _GEN_98 ? _double_bytes_0_T_8 : _GEN_1941; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1943 = 8'h49 == _GEN_98 ? _double_bytes_0_T_9 : _GEN_1942; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1944 = 8'h4a == _GEN_98 ? _double_bytes_0_T_10 : _GEN_1943; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1945 = 8'h4b == _GEN_98 ? _double_bytes_0_T_11 : _GEN_1944; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1946 = 8'h4c == _GEN_98 ? _double_bytes_0_T_12 : _GEN_1945; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1947 = 8'h4d == _GEN_98 ? _double_bytes_0_T_13 : _GEN_1946; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1948 = 8'h4e == _GEN_98 ? _double_bytes_0_T_14 : _GEN_1947; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1949 = 8'h4f == _GEN_98 ? _double_bytes_0_T_15 : _GEN_1948; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1950 = 8'h50 == _GEN_98 ? _double_bytes_0_T_16 : _GEN_1949; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1951 = 8'h51 == _GEN_98 ? _double_bytes_0_T_17 : _GEN_1950; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1952 = 8'h52 == _GEN_98 ? _double_bytes_0_T_18 : _GEN_1951; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1953 = 8'h53 == _GEN_98 ? _double_bytes_0_T_19 : _GEN_1952; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1954 = 8'h54 == _GEN_98 ? _double_bytes_0_T_20 : _GEN_1953; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1955 = 8'h55 == _GEN_98 ? _double_bytes_0_T_21 : _GEN_1954; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1956 = 8'h56 == _GEN_98 ? _double_bytes_0_T_22 : _GEN_1955; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1957 = 8'h57 == _GEN_98 ? _double_bytes_0_T_23 : _GEN_1956; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1958 = 8'h58 == _GEN_98 ? _double_bytes_0_T_24 : _GEN_1957; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1959 = 8'h59 == _GEN_98 ? _double_bytes_0_T_25 : _GEN_1958; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1960 = 8'h5a == _GEN_98 ? _double_bytes_0_T_26 : _GEN_1959; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1961 = 8'h5b == _GEN_98 ? _double_bytes_0_T_27 : _GEN_1960; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1962 = 8'h5c == _GEN_98 ? _double_bytes_0_T_28 : _GEN_1961; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1963 = 8'h5d == _GEN_98 ? _double_bytes_0_T_29 : _GEN_1962; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1964 = 8'h5e == _GEN_98 ? _double_bytes_0_T_30 : _GEN_1963; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1965 = 8'h5f == _GEN_98 ? _double_bytes_0_T_31 : _GEN_1964; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1966 = 8'h60 == _GEN_98 ? _double_bytes_0_T_32 : _GEN_1965; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1967 = 8'h61 == _GEN_98 ? _double_bytes_0_T_33 : _GEN_1966; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1968 = 8'h62 == _GEN_98 ? _double_bytes_0_T_34 : _GEN_1967; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1969 = 8'h63 == _GEN_98 ? _double_bytes_0_T_35 : _GEN_1968; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1970 = 8'h64 == _GEN_98 ? _double_bytes_0_T_36 : _GEN_1969; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1971 = 8'h65 == _GEN_98 ? _double_bytes_0_T_37 : _GEN_1970; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1972 = 8'h66 == _GEN_98 ? _double_bytes_0_T_38 : _GEN_1971; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1973 = 8'h67 == _GEN_98 ? _double_bytes_0_T_39 : _GEN_1972; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1974 = 8'h68 == _GEN_98 ? _double_bytes_0_T_40 : _GEN_1973; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1975 = 8'h69 == _GEN_98 ? _double_bytes_0_T_41 : _GEN_1974; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1976 = 8'h6a == _GEN_98 ? _double_bytes_0_T_42 : _GEN_1975; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1977 = 8'h6b == _GEN_98 ? _double_bytes_0_T_43 : _GEN_1976; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1978 = 8'h6c == _GEN_98 ? _double_bytes_0_T_44 : _GEN_1977; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1979 = 8'h6d == _GEN_98 ? _double_bytes_0_T_45 : _GEN_1978; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1980 = 8'h6e == _GEN_98 ? _double_bytes_0_T_46 : _GEN_1979; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1981 = 8'h6f == _GEN_98 ? _double_bytes_0_T_47 : _GEN_1980; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1982 = 8'h70 == _GEN_98 ? _double_bytes_0_T_48 : _GEN_1981; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1983 = 8'h71 == _GEN_98 ? _double_bytes_0_T_49 : _GEN_1982; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1984 = 8'h72 == _GEN_98 ? _double_bytes_0_T_50 : _GEN_1983; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1985 = 8'h73 == _GEN_98 ? _double_bytes_0_T_51 : _GEN_1984; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1986 = 8'h74 == _GEN_98 ? _double_bytes_0_T_52 : _GEN_1985; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1987 = 8'h75 == _GEN_98 ? _double_bytes_0_T_53 : _GEN_1986; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1988 = 8'h76 == _GEN_98 ? _double_bytes_0_T_54 : _GEN_1987; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1989 = 8'h77 == _GEN_98 ? _double_bytes_0_T_55 : _GEN_1988; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1990 = 8'h78 == _GEN_98 ? _double_bytes_0_T_56 : _GEN_1989; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1991 = 8'h79 == _GEN_98 ? _double_bytes_0_T_57 : _GEN_1990; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1992 = 8'h7a == _GEN_98 ? _double_bytes_0_T_58 : _GEN_1991; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1993 = 8'h7b == _GEN_98 ? _double_bytes_0_T_59 : _GEN_1992; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1994 = 8'h7c == _GEN_98 ? _double_bytes_0_T_60 : _GEN_1993; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1995 = 8'h7d == _GEN_98 ? _double_bytes_0_T_61 : _GEN_1994; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1996 = 8'h7e == _GEN_98 ? _double_bytes_0_T_62 : _GEN_1995; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1997 = 8'h7f == _GEN_98 ? _double_bytes_0_T_63 : _GEN_1996; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1998 = 8'h80 == _GEN_98 ? _double_bytes_0_T_64 : _GEN_1997; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1999 = 8'h81 == _GEN_98 ? _double_bytes_0_T_65 : _GEN_1998; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2000 = 8'h82 == _GEN_98 ? _double_bytes_0_T_66 : _GEN_1999; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2001 = 8'h83 == _GEN_98 ? _double_bytes_0_T_67 : _GEN_2000; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2002 = 8'h84 == _GEN_98 ? _double_bytes_0_T_68 : _GEN_2001; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2003 = 8'h85 == _GEN_98 ? _double_bytes_0_T_69 : _GEN_2002; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2004 = 8'h86 == _GEN_98 ? _double_bytes_0_T_70 : _GEN_2003; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2005 = 8'h87 == _GEN_98 ? _double_bytes_0_T_71 : _GEN_2004; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2006 = 8'h88 == _GEN_98 ? _double_bytes_0_T_72 : _GEN_2005; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2007 = 8'h89 == _GEN_98 ? _double_bytes_0_T_73 : _GEN_2006; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2008 = 8'h8a == _GEN_98 ? _double_bytes_0_T_74 : _GEN_2007; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2009 = 8'h8b == _GEN_98 ? _double_bytes_0_T_75 : _GEN_2008; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2010 = 8'h8c == _GEN_98 ? _double_bytes_0_T_76 : _GEN_2009; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2011 = 8'h8d == _GEN_98 ? _double_bytes_0_T_77 : _GEN_2010; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2012 = 8'h8e == _GEN_98 ? _double_bytes_0_T_78 : _GEN_2011; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2013 = 8'h8f == _GEN_98 ? _double_bytes_0_T_79 : _GEN_2012; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2014 = 8'h90 == _GEN_98 ? _double_bytes_0_T_80 : _GEN_2013; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2015 = 8'h91 == _GEN_98 ? _double_bytes_0_T_81 : _GEN_2014; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2016 = 8'h92 == _GEN_98 ? _double_bytes_0_T_82 : _GEN_2015; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2017 = 8'h93 == _GEN_98 ? _double_bytes_0_T_83 : _GEN_2016; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2018 = 8'h94 == _GEN_98 ? _double_bytes_0_T_84 : _GEN_2017; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2019 = 8'h95 == _GEN_98 ? _double_bytes_0_T_85 : _GEN_2018; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2020 = 8'h96 == _GEN_98 ? _double_bytes_0_T_86 : _GEN_2019; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2021 = 8'h97 == _GEN_98 ? _double_bytes_0_T_87 : _GEN_2020; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2022 = 8'h98 == _GEN_98 ? _double_bytes_0_T_88 : _GEN_2021; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2023 = 8'h99 == _GEN_98 ? _double_bytes_0_T_89 : _GEN_2022; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2024 = 8'h9a == _GEN_98 ? _double_bytes_0_T_90 : _GEN_2023; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2025 = 8'h9b == _GEN_98 ? _double_bytes_0_T_91 : _GEN_2024; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2026 = 8'h9c == _GEN_98 ? _double_bytes_0_T_92 : _GEN_2025; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2027 = 8'h9d == _GEN_98 ? _double_bytes_0_T_93 : _GEN_2026; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2028 = 8'h9e == _GEN_98 ? _double_bytes_0_T_94 : _GEN_2027; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2029 = 8'h9f == _GEN_98 ? _double_bytes_0_T_95 : _GEN_2028; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] double_bytes_3_0 = _GEN_74 ? _GEN_2029 : 16'h0; // @[matcher_pisa.scala 145:46 matcher_pisa.scala 144:41]
  wire [15:0] _GEN_2031 = 8'h40 == _GEN_99 ? _double_bytes_0_T : 16'h0; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53 matcher_pisa.scala 144:41]
  wire [15:0] _GEN_2032 = 8'h41 == _GEN_99 ? _double_bytes_0_T_1 : _GEN_2031; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2033 = 8'h42 == _GEN_99 ? _double_bytes_0_T_2 : _GEN_2032; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2034 = 8'h43 == _GEN_99 ? _double_bytes_0_T_3 : _GEN_2033; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2035 = 8'h44 == _GEN_99 ? _double_bytes_0_T_4 : _GEN_2034; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2036 = 8'h45 == _GEN_99 ? _double_bytes_0_T_5 : _GEN_2035; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2037 = 8'h46 == _GEN_99 ? _double_bytes_0_T_6 : _GEN_2036; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2038 = 8'h47 == _GEN_99 ? _double_bytes_0_T_7 : _GEN_2037; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2039 = 8'h48 == _GEN_99 ? _double_bytes_0_T_8 : _GEN_2038; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2040 = 8'h49 == _GEN_99 ? _double_bytes_0_T_9 : _GEN_2039; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2041 = 8'h4a == _GEN_99 ? _double_bytes_0_T_10 : _GEN_2040; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2042 = 8'h4b == _GEN_99 ? _double_bytes_0_T_11 : _GEN_2041; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2043 = 8'h4c == _GEN_99 ? _double_bytes_0_T_12 : _GEN_2042; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2044 = 8'h4d == _GEN_99 ? _double_bytes_0_T_13 : _GEN_2043; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2045 = 8'h4e == _GEN_99 ? _double_bytes_0_T_14 : _GEN_2044; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2046 = 8'h4f == _GEN_99 ? _double_bytes_0_T_15 : _GEN_2045; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2047 = 8'h50 == _GEN_99 ? _double_bytes_0_T_16 : _GEN_2046; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2048 = 8'h51 == _GEN_99 ? _double_bytes_0_T_17 : _GEN_2047; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2049 = 8'h52 == _GEN_99 ? _double_bytes_0_T_18 : _GEN_2048; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2050 = 8'h53 == _GEN_99 ? _double_bytes_0_T_19 : _GEN_2049; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2051 = 8'h54 == _GEN_99 ? _double_bytes_0_T_20 : _GEN_2050; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2052 = 8'h55 == _GEN_99 ? _double_bytes_0_T_21 : _GEN_2051; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2053 = 8'h56 == _GEN_99 ? _double_bytes_0_T_22 : _GEN_2052; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2054 = 8'h57 == _GEN_99 ? _double_bytes_0_T_23 : _GEN_2053; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2055 = 8'h58 == _GEN_99 ? _double_bytes_0_T_24 : _GEN_2054; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2056 = 8'h59 == _GEN_99 ? _double_bytes_0_T_25 : _GEN_2055; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2057 = 8'h5a == _GEN_99 ? _double_bytes_0_T_26 : _GEN_2056; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2058 = 8'h5b == _GEN_99 ? _double_bytes_0_T_27 : _GEN_2057; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2059 = 8'h5c == _GEN_99 ? _double_bytes_0_T_28 : _GEN_2058; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2060 = 8'h5d == _GEN_99 ? _double_bytes_0_T_29 : _GEN_2059; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2061 = 8'h5e == _GEN_99 ? _double_bytes_0_T_30 : _GEN_2060; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2062 = 8'h5f == _GEN_99 ? _double_bytes_0_T_31 : _GEN_2061; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2063 = 8'h60 == _GEN_99 ? _double_bytes_0_T_32 : _GEN_2062; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2064 = 8'h61 == _GEN_99 ? _double_bytes_0_T_33 : _GEN_2063; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2065 = 8'h62 == _GEN_99 ? _double_bytes_0_T_34 : _GEN_2064; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2066 = 8'h63 == _GEN_99 ? _double_bytes_0_T_35 : _GEN_2065; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2067 = 8'h64 == _GEN_99 ? _double_bytes_0_T_36 : _GEN_2066; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2068 = 8'h65 == _GEN_99 ? _double_bytes_0_T_37 : _GEN_2067; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2069 = 8'h66 == _GEN_99 ? _double_bytes_0_T_38 : _GEN_2068; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2070 = 8'h67 == _GEN_99 ? _double_bytes_0_T_39 : _GEN_2069; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2071 = 8'h68 == _GEN_99 ? _double_bytes_0_T_40 : _GEN_2070; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2072 = 8'h69 == _GEN_99 ? _double_bytes_0_T_41 : _GEN_2071; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2073 = 8'h6a == _GEN_99 ? _double_bytes_0_T_42 : _GEN_2072; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2074 = 8'h6b == _GEN_99 ? _double_bytes_0_T_43 : _GEN_2073; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2075 = 8'h6c == _GEN_99 ? _double_bytes_0_T_44 : _GEN_2074; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2076 = 8'h6d == _GEN_99 ? _double_bytes_0_T_45 : _GEN_2075; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2077 = 8'h6e == _GEN_99 ? _double_bytes_0_T_46 : _GEN_2076; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2078 = 8'h6f == _GEN_99 ? _double_bytes_0_T_47 : _GEN_2077; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2079 = 8'h70 == _GEN_99 ? _double_bytes_0_T_48 : _GEN_2078; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2080 = 8'h71 == _GEN_99 ? _double_bytes_0_T_49 : _GEN_2079; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2081 = 8'h72 == _GEN_99 ? _double_bytes_0_T_50 : _GEN_2080; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2082 = 8'h73 == _GEN_99 ? _double_bytes_0_T_51 : _GEN_2081; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2083 = 8'h74 == _GEN_99 ? _double_bytes_0_T_52 : _GEN_2082; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2084 = 8'h75 == _GEN_99 ? _double_bytes_0_T_53 : _GEN_2083; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2085 = 8'h76 == _GEN_99 ? _double_bytes_0_T_54 : _GEN_2084; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2086 = 8'h77 == _GEN_99 ? _double_bytes_0_T_55 : _GEN_2085; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2087 = 8'h78 == _GEN_99 ? _double_bytes_0_T_56 : _GEN_2086; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2088 = 8'h79 == _GEN_99 ? _double_bytes_0_T_57 : _GEN_2087; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2089 = 8'h7a == _GEN_99 ? _double_bytes_0_T_58 : _GEN_2088; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2090 = 8'h7b == _GEN_99 ? _double_bytes_0_T_59 : _GEN_2089; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2091 = 8'h7c == _GEN_99 ? _double_bytes_0_T_60 : _GEN_2090; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2092 = 8'h7d == _GEN_99 ? _double_bytes_0_T_61 : _GEN_2091; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2093 = 8'h7e == _GEN_99 ? _double_bytes_0_T_62 : _GEN_2092; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2094 = 8'h7f == _GEN_99 ? _double_bytes_0_T_63 : _GEN_2093; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2095 = 8'h80 == _GEN_99 ? _double_bytes_0_T_64 : _GEN_2094; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2096 = 8'h81 == _GEN_99 ? _double_bytes_0_T_65 : _GEN_2095; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2097 = 8'h82 == _GEN_99 ? _double_bytes_0_T_66 : _GEN_2096; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2098 = 8'h83 == _GEN_99 ? _double_bytes_0_T_67 : _GEN_2097; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2099 = 8'h84 == _GEN_99 ? _double_bytes_0_T_68 : _GEN_2098; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2100 = 8'h85 == _GEN_99 ? _double_bytes_0_T_69 : _GEN_2099; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2101 = 8'h86 == _GEN_99 ? _double_bytes_0_T_70 : _GEN_2100; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2102 = 8'h87 == _GEN_99 ? _double_bytes_0_T_71 : _GEN_2101; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2103 = 8'h88 == _GEN_99 ? _double_bytes_0_T_72 : _GEN_2102; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2104 = 8'h89 == _GEN_99 ? _double_bytes_0_T_73 : _GEN_2103; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2105 = 8'h8a == _GEN_99 ? _double_bytes_0_T_74 : _GEN_2104; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2106 = 8'h8b == _GEN_99 ? _double_bytes_0_T_75 : _GEN_2105; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2107 = 8'h8c == _GEN_99 ? _double_bytes_0_T_76 : _GEN_2106; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2108 = 8'h8d == _GEN_99 ? _double_bytes_0_T_77 : _GEN_2107; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2109 = 8'h8e == _GEN_99 ? _double_bytes_0_T_78 : _GEN_2108; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2110 = 8'h8f == _GEN_99 ? _double_bytes_0_T_79 : _GEN_2109; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2111 = 8'h90 == _GEN_99 ? _double_bytes_0_T_80 : _GEN_2110; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2112 = 8'h91 == _GEN_99 ? _double_bytes_0_T_81 : _GEN_2111; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2113 = 8'h92 == _GEN_99 ? _double_bytes_0_T_82 : _GEN_2112; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2114 = 8'h93 == _GEN_99 ? _double_bytes_0_T_83 : _GEN_2113; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2115 = 8'h94 == _GEN_99 ? _double_bytes_0_T_84 : _GEN_2114; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2116 = 8'h95 == _GEN_99 ? _double_bytes_0_T_85 : _GEN_2115; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2117 = 8'h96 == _GEN_99 ? _double_bytes_0_T_86 : _GEN_2116; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2118 = 8'h97 == _GEN_99 ? _double_bytes_0_T_87 : _GEN_2117; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2119 = 8'h98 == _GEN_99 ? _double_bytes_0_T_88 : _GEN_2118; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2120 = 8'h99 == _GEN_99 ? _double_bytes_0_T_89 : _GEN_2119; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2121 = 8'h9a == _GEN_99 ? _double_bytes_0_T_90 : _GEN_2120; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2122 = 8'h9b == _GEN_99 ? _double_bytes_0_T_91 : _GEN_2121; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2123 = 8'h9c == _GEN_99 ? _double_bytes_0_T_92 : _GEN_2122; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2124 = 8'h9d == _GEN_99 ? _double_bytes_0_T_93 : _GEN_2123; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2125 = 8'h9e == _GEN_99 ? _double_bytes_0_T_94 : _GEN_2124; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2126 = 8'h9f == _GEN_99 ? _double_bytes_0_T_95 : _GEN_2125; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] double_bytes_3_1 = _GEN_75 ? _GEN_2126 : 16'h0; // @[matcher_pisa.scala 145:46 matcher_pisa.scala 144:41]
  wire [31:0] _groups_3_T_1 = {double_bytes_3_0,double_bytes_3_1}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_2128 = _GEN_59 == 2'h2 ? _groups_3_T_1 : _GEN_1933; // @[matcher_pisa.scala 139:50 matcher_pisa.scala 153:31]
  wire [31:0] _GEN_2129 = 8'ha0 == _GEN_98 ? _groups_0_T_2 : 32'h0; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39 matcher_pisa.scala 158:31]
  wire [31:0] _GEN_2130 = 8'ha1 == _GEN_98 ? _groups_0_T_3 : _GEN_2129; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2131 = 8'ha2 == _GEN_98 ? _groups_0_T_4 : _GEN_2130; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2132 = 8'ha3 == _GEN_98 ? _groups_0_T_5 : _GEN_2131; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2133 = 8'ha4 == _GEN_98 ? _groups_0_T_6 : _GEN_2132; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2134 = 8'ha5 == _GEN_98 ? _groups_0_T_7 : _GEN_2133; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2135 = 8'ha6 == _GEN_98 ? _groups_0_T_8 : _GEN_2134; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2136 = 8'ha7 == _GEN_98 ? _groups_0_T_9 : _GEN_2135; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2137 = 8'ha8 == _GEN_98 ? _groups_0_T_10 : _GEN_2136; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2138 = 8'ha9 == _GEN_98 ? _groups_0_T_11 : _GEN_2137; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2139 = 8'haa == _GEN_98 ? _groups_0_T_12 : _GEN_2138; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2140 = 8'hab == _GEN_98 ? _groups_0_T_13 : _GEN_2139; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2141 = 8'hac == _GEN_98 ? _groups_0_T_14 : _GEN_2140; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2142 = 8'had == _GEN_98 ? _groups_0_T_15 : _GEN_2141; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2143 = 8'hae == _GEN_98 ? _groups_0_T_16 : _GEN_2142; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2144 = 8'haf == _GEN_98 ? _groups_0_T_17 : _GEN_2143; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2145 = 8'hb0 == _GEN_98 ? _groups_0_T_18 : _GEN_2144; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2146 = 8'hb1 == _GEN_98 ? _groups_0_T_19 : _GEN_2145; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2147 = 8'hb2 == _GEN_98 ? _groups_0_T_20 : _GEN_2146; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2148 = 8'hb3 == _GEN_98 ? _groups_0_T_21 : _GEN_2147; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2149 = 8'hb4 == _GEN_98 ? _groups_0_T_22 : _GEN_2148; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2150 = 8'hb5 == _GEN_98 ? _groups_0_T_23 : _GEN_2149; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2151 = 8'hb6 == _GEN_98 ? _groups_0_T_24 : _GEN_2150; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2152 = 8'hb7 == _GEN_98 ? _groups_0_T_25 : _GEN_2151; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2153 = 8'hb8 == _GEN_98 ? _groups_0_T_26 : _GEN_2152; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2154 = 8'hb9 == _GEN_98 ? _groups_0_T_27 : _GEN_2153; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2155 = 8'hba == _GEN_98 ? _groups_0_T_28 : _GEN_2154; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2156 = 8'hbb == _GEN_98 ? _groups_0_T_29 : _GEN_2155; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2157 = 8'hbc == _GEN_98 ? _groups_0_T_30 : _GEN_2156; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2158 = 8'hbd == _GEN_98 ? _groups_0_T_31 : _GEN_2157; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2159 = 8'hbe == _GEN_98 ? _groups_0_T_32 : _GEN_2158; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2160 = 8'hbf == _GEN_98 ? _groups_0_T_33 : _GEN_2159; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2161 = 8'hc0 == _GEN_98 ? _groups_0_T_34 : _GEN_2160; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2162 = 8'hc1 == _GEN_98 ? _groups_0_T_35 : _GEN_2161; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2163 = 8'hc2 == _GEN_98 ? _groups_0_T_36 : _GEN_2162; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2164 = 8'hc3 == _GEN_98 ? _groups_0_T_37 : _GEN_2163; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2165 = 8'hc4 == _GEN_98 ? _groups_0_T_38 : _GEN_2164; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2166 = 8'hc5 == _GEN_98 ? _groups_0_T_39 : _GEN_2165; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2167 = 8'hc6 == _GEN_98 ? _groups_0_T_40 : _GEN_2166; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2168 = 8'hc7 == _GEN_98 ? _groups_0_T_41 : _GEN_2167; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2169 = 8'hc8 == _GEN_98 ? _groups_0_T_42 : _GEN_2168; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2170 = 8'hc9 == _GEN_98 ? _groups_0_T_43 : _GEN_2169; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2171 = 8'hca == _GEN_98 ? _groups_0_T_44 : _GEN_2170; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2172 = 8'hcb == _GEN_98 ? _groups_0_T_45 : _GEN_2171; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2173 = 8'hcc == _GEN_98 ? _groups_0_T_46 : _GEN_2172; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2174 = 8'hcd == _GEN_98 ? _groups_0_T_47 : _GEN_2173; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2175 = 8'hce == _GEN_98 ? _groups_0_T_48 : _GEN_2174; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2176 = 8'hcf == _GEN_98 ? _groups_0_T_49 : _GEN_2175; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2177 = 8'hd0 == _GEN_98 ? _groups_0_T_50 : _GEN_2176; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2178 = 8'hd1 == _GEN_98 ? _groups_0_T_51 : _GEN_2177; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2179 = 8'hd2 == _GEN_98 ? _groups_0_T_52 : _GEN_2178; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2180 = 8'hd3 == _GEN_98 ? _groups_0_T_53 : _GEN_2179; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2181 = 8'hd4 == _GEN_98 ? _groups_0_T_54 : _GEN_2180; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2182 = 8'hd5 == _GEN_98 ? _groups_0_T_55 : _GEN_2181; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2183 = 8'hd6 == _GEN_98 ? _groups_0_T_56 : _GEN_2182; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2184 = 8'hd7 == _GEN_98 ? _groups_0_T_57 : _GEN_2183; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2185 = 8'hd8 == _GEN_98 ? _groups_0_T_58 : _GEN_2184; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2186 = 8'hd9 == _GEN_98 ? _groups_0_T_59 : _GEN_2185; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2187 = 8'hda == _GEN_98 ? _groups_0_T_60 : _GEN_2186; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2188 = 8'hdb == _GEN_98 ? _groups_0_T_61 : _GEN_2187; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2189 = 8'hdc == _GEN_98 ? _groups_0_T_62 : _GEN_2188; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2190 = 8'hdd == _GEN_98 ? _groups_0_T_63 : _GEN_2189; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2191 = 8'hde == _GEN_98 ? _groups_0_T_64 : _GEN_2190; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2192 = 8'hdf == _GEN_98 ? _groups_0_T_65 : _GEN_2191; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] groups_3 = _GEN_59 == 2'h3 ? _GEN_2192 : _GEN_2128; // @[matcher_pisa.scala 155:50]
  wire [7:0] _GEN_2194 = 8'h0 == _GEN_102 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_2195 = 8'h1 == _GEN_102 ? phv_data_1 : _GEN_2194; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2196 = 8'h2 == _GEN_102 ? phv_data_2 : _GEN_2195; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2197 = 8'h3 == _GEN_102 ? phv_data_3 : _GEN_2196; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2198 = 8'h4 == _GEN_102 ? phv_data_4 : _GEN_2197; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2199 = 8'h5 == _GEN_102 ? phv_data_5 : _GEN_2198; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2200 = 8'h6 == _GEN_102 ? phv_data_6 : _GEN_2199; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2201 = 8'h7 == _GEN_102 ? phv_data_7 : _GEN_2200; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2202 = 8'h8 == _GEN_102 ? phv_data_8 : _GEN_2201; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2203 = 8'h9 == _GEN_102 ? phv_data_9 : _GEN_2202; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2204 = 8'ha == _GEN_102 ? phv_data_10 : _GEN_2203; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2205 = 8'hb == _GEN_102 ? phv_data_11 : _GEN_2204; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2206 = 8'hc == _GEN_102 ? phv_data_12 : _GEN_2205; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2207 = 8'hd == _GEN_102 ? phv_data_13 : _GEN_2206; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2208 = 8'he == _GEN_102 ? phv_data_14 : _GEN_2207; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2209 = 8'hf == _GEN_102 ? phv_data_15 : _GEN_2208; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2210 = 8'h10 == _GEN_102 ? phv_data_16 : _GEN_2209; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2211 = 8'h11 == _GEN_102 ? phv_data_17 : _GEN_2210; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2212 = 8'h12 == _GEN_102 ? phv_data_18 : _GEN_2211; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2213 = 8'h13 == _GEN_102 ? phv_data_19 : _GEN_2212; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2214 = 8'h14 == _GEN_102 ? phv_data_20 : _GEN_2213; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2215 = 8'h15 == _GEN_102 ? phv_data_21 : _GEN_2214; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2216 = 8'h16 == _GEN_102 ? phv_data_22 : _GEN_2215; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2217 = 8'h17 == _GEN_102 ? phv_data_23 : _GEN_2216; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2218 = 8'h18 == _GEN_102 ? phv_data_24 : _GEN_2217; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2219 = 8'h19 == _GEN_102 ? phv_data_25 : _GEN_2218; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2220 = 8'h1a == _GEN_102 ? phv_data_26 : _GEN_2219; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2221 = 8'h1b == _GEN_102 ? phv_data_27 : _GEN_2220; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2222 = 8'h1c == _GEN_102 ? phv_data_28 : _GEN_2221; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2223 = 8'h1d == _GEN_102 ? phv_data_29 : _GEN_2222; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2224 = 8'h1e == _GEN_102 ? phv_data_30 : _GEN_2223; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2225 = 8'h1f == _GEN_102 ? phv_data_31 : _GEN_2224; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2226 = 8'h20 == _GEN_102 ? phv_data_32 : _GEN_2225; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2227 = 8'h21 == _GEN_102 ? phv_data_33 : _GEN_2226; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2228 = 8'h22 == _GEN_102 ? phv_data_34 : _GEN_2227; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2229 = 8'h23 == _GEN_102 ? phv_data_35 : _GEN_2228; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2230 = 8'h24 == _GEN_102 ? phv_data_36 : _GEN_2229; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2231 = 8'h25 == _GEN_102 ? phv_data_37 : _GEN_2230; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2232 = 8'h26 == _GEN_102 ? phv_data_38 : _GEN_2231; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2233 = 8'h27 == _GEN_102 ? phv_data_39 : _GEN_2232; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2234 = 8'h28 == _GEN_102 ? phv_data_40 : _GEN_2233; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2235 = 8'h29 == _GEN_102 ? phv_data_41 : _GEN_2234; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2236 = 8'h2a == _GEN_102 ? phv_data_42 : _GEN_2235; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2237 = 8'h2b == _GEN_102 ? phv_data_43 : _GEN_2236; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2238 = 8'h2c == _GEN_102 ? phv_data_44 : _GEN_2237; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2239 = 8'h2d == _GEN_102 ? phv_data_45 : _GEN_2238; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2240 = 8'h2e == _GEN_102 ? phv_data_46 : _GEN_2239; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2241 = 8'h2f == _GEN_102 ? phv_data_47 : _GEN_2240; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2242 = 8'h30 == _GEN_102 ? phv_data_48 : _GEN_2241; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2243 = 8'h31 == _GEN_102 ? phv_data_49 : _GEN_2242; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2244 = 8'h32 == _GEN_102 ? phv_data_50 : _GEN_2243; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2245 = 8'h33 == _GEN_102 ? phv_data_51 : _GEN_2244; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2246 = 8'h34 == _GEN_102 ? phv_data_52 : _GEN_2245; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2247 = 8'h35 == _GEN_102 ? phv_data_53 : _GEN_2246; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2248 = 8'h36 == _GEN_102 ? phv_data_54 : _GEN_2247; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2249 = 8'h37 == _GEN_102 ? phv_data_55 : _GEN_2248; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2250 = 8'h38 == _GEN_102 ? phv_data_56 : _GEN_2249; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2251 = 8'h39 == _GEN_102 ? phv_data_57 : _GEN_2250; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2252 = 8'h3a == _GEN_102 ? phv_data_58 : _GEN_2251; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2253 = 8'h3b == _GEN_102 ? phv_data_59 : _GEN_2252; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2254 = 8'h3c == _GEN_102 ? phv_data_60 : _GEN_2253; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2255 = 8'h3d == _GEN_102 ? phv_data_61 : _GEN_2254; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2256 = 8'h3e == _GEN_102 ? phv_data_62 : _GEN_2255; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2257 = 8'h3f == _GEN_102 ? phv_data_63 : _GEN_2256; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] bytes_4_0 = _GEN_78 ? _GEN_2257 : 8'h0; // @[matcher_pisa.scala 129:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_2259 = 8'h0 == _GEN_103 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_2260 = 8'h1 == _GEN_103 ? phv_data_1 : _GEN_2259; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2261 = 8'h2 == _GEN_103 ? phv_data_2 : _GEN_2260; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2262 = 8'h3 == _GEN_103 ? phv_data_3 : _GEN_2261; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2263 = 8'h4 == _GEN_103 ? phv_data_4 : _GEN_2262; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2264 = 8'h5 == _GEN_103 ? phv_data_5 : _GEN_2263; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2265 = 8'h6 == _GEN_103 ? phv_data_6 : _GEN_2264; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2266 = 8'h7 == _GEN_103 ? phv_data_7 : _GEN_2265; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2267 = 8'h8 == _GEN_103 ? phv_data_8 : _GEN_2266; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2268 = 8'h9 == _GEN_103 ? phv_data_9 : _GEN_2267; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2269 = 8'ha == _GEN_103 ? phv_data_10 : _GEN_2268; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2270 = 8'hb == _GEN_103 ? phv_data_11 : _GEN_2269; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2271 = 8'hc == _GEN_103 ? phv_data_12 : _GEN_2270; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2272 = 8'hd == _GEN_103 ? phv_data_13 : _GEN_2271; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2273 = 8'he == _GEN_103 ? phv_data_14 : _GEN_2272; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2274 = 8'hf == _GEN_103 ? phv_data_15 : _GEN_2273; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2275 = 8'h10 == _GEN_103 ? phv_data_16 : _GEN_2274; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2276 = 8'h11 == _GEN_103 ? phv_data_17 : _GEN_2275; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2277 = 8'h12 == _GEN_103 ? phv_data_18 : _GEN_2276; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2278 = 8'h13 == _GEN_103 ? phv_data_19 : _GEN_2277; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2279 = 8'h14 == _GEN_103 ? phv_data_20 : _GEN_2278; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2280 = 8'h15 == _GEN_103 ? phv_data_21 : _GEN_2279; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2281 = 8'h16 == _GEN_103 ? phv_data_22 : _GEN_2280; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2282 = 8'h17 == _GEN_103 ? phv_data_23 : _GEN_2281; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2283 = 8'h18 == _GEN_103 ? phv_data_24 : _GEN_2282; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2284 = 8'h19 == _GEN_103 ? phv_data_25 : _GEN_2283; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2285 = 8'h1a == _GEN_103 ? phv_data_26 : _GEN_2284; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2286 = 8'h1b == _GEN_103 ? phv_data_27 : _GEN_2285; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2287 = 8'h1c == _GEN_103 ? phv_data_28 : _GEN_2286; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2288 = 8'h1d == _GEN_103 ? phv_data_29 : _GEN_2287; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2289 = 8'h1e == _GEN_103 ? phv_data_30 : _GEN_2288; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2290 = 8'h1f == _GEN_103 ? phv_data_31 : _GEN_2289; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2291 = 8'h20 == _GEN_103 ? phv_data_32 : _GEN_2290; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2292 = 8'h21 == _GEN_103 ? phv_data_33 : _GEN_2291; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2293 = 8'h22 == _GEN_103 ? phv_data_34 : _GEN_2292; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2294 = 8'h23 == _GEN_103 ? phv_data_35 : _GEN_2293; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2295 = 8'h24 == _GEN_103 ? phv_data_36 : _GEN_2294; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2296 = 8'h25 == _GEN_103 ? phv_data_37 : _GEN_2295; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2297 = 8'h26 == _GEN_103 ? phv_data_38 : _GEN_2296; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2298 = 8'h27 == _GEN_103 ? phv_data_39 : _GEN_2297; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2299 = 8'h28 == _GEN_103 ? phv_data_40 : _GEN_2298; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2300 = 8'h29 == _GEN_103 ? phv_data_41 : _GEN_2299; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2301 = 8'h2a == _GEN_103 ? phv_data_42 : _GEN_2300; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2302 = 8'h2b == _GEN_103 ? phv_data_43 : _GEN_2301; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2303 = 8'h2c == _GEN_103 ? phv_data_44 : _GEN_2302; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2304 = 8'h2d == _GEN_103 ? phv_data_45 : _GEN_2303; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2305 = 8'h2e == _GEN_103 ? phv_data_46 : _GEN_2304; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2306 = 8'h2f == _GEN_103 ? phv_data_47 : _GEN_2305; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2307 = 8'h30 == _GEN_103 ? phv_data_48 : _GEN_2306; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2308 = 8'h31 == _GEN_103 ? phv_data_49 : _GEN_2307; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2309 = 8'h32 == _GEN_103 ? phv_data_50 : _GEN_2308; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2310 = 8'h33 == _GEN_103 ? phv_data_51 : _GEN_2309; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2311 = 8'h34 == _GEN_103 ? phv_data_52 : _GEN_2310; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2312 = 8'h35 == _GEN_103 ? phv_data_53 : _GEN_2311; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2313 = 8'h36 == _GEN_103 ? phv_data_54 : _GEN_2312; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2314 = 8'h37 == _GEN_103 ? phv_data_55 : _GEN_2313; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2315 = 8'h38 == _GEN_103 ? phv_data_56 : _GEN_2314; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2316 = 8'h39 == _GEN_103 ? phv_data_57 : _GEN_2315; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2317 = 8'h3a == _GEN_103 ? phv_data_58 : _GEN_2316; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2318 = 8'h3b == _GEN_103 ? phv_data_59 : _GEN_2317; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2319 = 8'h3c == _GEN_103 ? phv_data_60 : _GEN_2318; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2320 = 8'h3d == _GEN_103 ? phv_data_61 : _GEN_2319; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2321 = 8'h3e == _GEN_103 ? phv_data_62 : _GEN_2320; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2322 = 8'h3f == _GEN_103 ? phv_data_63 : _GEN_2321; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] bytes_4_1 = _GEN_79 ? _GEN_2322 : 8'h0; // @[matcher_pisa.scala 129:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_2324 = 8'h0 == _GEN_104 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_2325 = 8'h1 == _GEN_104 ? phv_data_1 : _GEN_2324; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2326 = 8'h2 == _GEN_104 ? phv_data_2 : _GEN_2325; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2327 = 8'h3 == _GEN_104 ? phv_data_3 : _GEN_2326; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2328 = 8'h4 == _GEN_104 ? phv_data_4 : _GEN_2327; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2329 = 8'h5 == _GEN_104 ? phv_data_5 : _GEN_2328; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2330 = 8'h6 == _GEN_104 ? phv_data_6 : _GEN_2329; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2331 = 8'h7 == _GEN_104 ? phv_data_7 : _GEN_2330; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2332 = 8'h8 == _GEN_104 ? phv_data_8 : _GEN_2331; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2333 = 8'h9 == _GEN_104 ? phv_data_9 : _GEN_2332; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2334 = 8'ha == _GEN_104 ? phv_data_10 : _GEN_2333; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2335 = 8'hb == _GEN_104 ? phv_data_11 : _GEN_2334; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2336 = 8'hc == _GEN_104 ? phv_data_12 : _GEN_2335; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2337 = 8'hd == _GEN_104 ? phv_data_13 : _GEN_2336; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2338 = 8'he == _GEN_104 ? phv_data_14 : _GEN_2337; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2339 = 8'hf == _GEN_104 ? phv_data_15 : _GEN_2338; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2340 = 8'h10 == _GEN_104 ? phv_data_16 : _GEN_2339; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2341 = 8'h11 == _GEN_104 ? phv_data_17 : _GEN_2340; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2342 = 8'h12 == _GEN_104 ? phv_data_18 : _GEN_2341; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2343 = 8'h13 == _GEN_104 ? phv_data_19 : _GEN_2342; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2344 = 8'h14 == _GEN_104 ? phv_data_20 : _GEN_2343; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2345 = 8'h15 == _GEN_104 ? phv_data_21 : _GEN_2344; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2346 = 8'h16 == _GEN_104 ? phv_data_22 : _GEN_2345; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2347 = 8'h17 == _GEN_104 ? phv_data_23 : _GEN_2346; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2348 = 8'h18 == _GEN_104 ? phv_data_24 : _GEN_2347; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2349 = 8'h19 == _GEN_104 ? phv_data_25 : _GEN_2348; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2350 = 8'h1a == _GEN_104 ? phv_data_26 : _GEN_2349; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2351 = 8'h1b == _GEN_104 ? phv_data_27 : _GEN_2350; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2352 = 8'h1c == _GEN_104 ? phv_data_28 : _GEN_2351; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2353 = 8'h1d == _GEN_104 ? phv_data_29 : _GEN_2352; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2354 = 8'h1e == _GEN_104 ? phv_data_30 : _GEN_2353; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2355 = 8'h1f == _GEN_104 ? phv_data_31 : _GEN_2354; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2356 = 8'h20 == _GEN_104 ? phv_data_32 : _GEN_2355; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2357 = 8'h21 == _GEN_104 ? phv_data_33 : _GEN_2356; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2358 = 8'h22 == _GEN_104 ? phv_data_34 : _GEN_2357; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2359 = 8'h23 == _GEN_104 ? phv_data_35 : _GEN_2358; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2360 = 8'h24 == _GEN_104 ? phv_data_36 : _GEN_2359; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2361 = 8'h25 == _GEN_104 ? phv_data_37 : _GEN_2360; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2362 = 8'h26 == _GEN_104 ? phv_data_38 : _GEN_2361; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2363 = 8'h27 == _GEN_104 ? phv_data_39 : _GEN_2362; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2364 = 8'h28 == _GEN_104 ? phv_data_40 : _GEN_2363; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2365 = 8'h29 == _GEN_104 ? phv_data_41 : _GEN_2364; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2366 = 8'h2a == _GEN_104 ? phv_data_42 : _GEN_2365; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2367 = 8'h2b == _GEN_104 ? phv_data_43 : _GEN_2366; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2368 = 8'h2c == _GEN_104 ? phv_data_44 : _GEN_2367; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2369 = 8'h2d == _GEN_104 ? phv_data_45 : _GEN_2368; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2370 = 8'h2e == _GEN_104 ? phv_data_46 : _GEN_2369; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2371 = 8'h2f == _GEN_104 ? phv_data_47 : _GEN_2370; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2372 = 8'h30 == _GEN_104 ? phv_data_48 : _GEN_2371; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2373 = 8'h31 == _GEN_104 ? phv_data_49 : _GEN_2372; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2374 = 8'h32 == _GEN_104 ? phv_data_50 : _GEN_2373; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2375 = 8'h33 == _GEN_104 ? phv_data_51 : _GEN_2374; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2376 = 8'h34 == _GEN_104 ? phv_data_52 : _GEN_2375; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2377 = 8'h35 == _GEN_104 ? phv_data_53 : _GEN_2376; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2378 = 8'h36 == _GEN_104 ? phv_data_54 : _GEN_2377; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2379 = 8'h37 == _GEN_104 ? phv_data_55 : _GEN_2378; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2380 = 8'h38 == _GEN_104 ? phv_data_56 : _GEN_2379; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2381 = 8'h39 == _GEN_104 ? phv_data_57 : _GEN_2380; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2382 = 8'h3a == _GEN_104 ? phv_data_58 : _GEN_2381; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2383 = 8'h3b == _GEN_104 ? phv_data_59 : _GEN_2382; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2384 = 8'h3c == _GEN_104 ? phv_data_60 : _GEN_2383; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2385 = 8'h3d == _GEN_104 ? phv_data_61 : _GEN_2384; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2386 = 8'h3e == _GEN_104 ? phv_data_62 : _GEN_2385; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2387 = 8'h3f == _GEN_104 ? phv_data_63 : _GEN_2386; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] bytes_4_2 = _GEN_80 ? _GEN_2387 : 8'h0; // @[matcher_pisa.scala 129:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_2389 = 8'h0 == _GEN_105 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_2390 = 8'h1 == _GEN_105 ? phv_data_1 : _GEN_2389; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2391 = 8'h2 == _GEN_105 ? phv_data_2 : _GEN_2390; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2392 = 8'h3 == _GEN_105 ? phv_data_3 : _GEN_2391; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2393 = 8'h4 == _GEN_105 ? phv_data_4 : _GEN_2392; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2394 = 8'h5 == _GEN_105 ? phv_data_5 : _GEN_2393; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2395 = 8'h6 == _GEN_105 ? phv_data_6 : _GEN_2394; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2396 = 8'h7 == _GEN_105 ? phv_data_7 : _GEN_2395; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2397 = 8'h8 == _GEN_105 ? phv_data_8 : _GEN_2396; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2398 = 8'h9 == _GEN_105 ? phv_data_9 : _GEN_2397; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2399 = 8'ha == _GEN_105 ? phv_data_10 : _GEN_2398; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2400 = 8'hb == _GEN_105 ? phv_data_11 : _GEN_2399; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2401 = 8'hc == _GEN_105 ? phv_data_12 : _GEN_2400; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2402 = 8'hd == _GEN_105 ? phv_data_13 : _GEN_2401; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2403 = 8'he == _GEN_105 ? phv_data_14 : _GEN_2402; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2404 = 8'hf == _GEN_105 ? phv_data_15 : _GEN_2403; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2405 = 8'h10 == _GEN_105 ? phv_data_16 : _GEN_2404; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2406 = 8'h11 == _GEN_105 ? phv_data_17 : _GEN_2405; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2407 = 8'h12 == _GEN_105 ? phv_data_18 : _GEN_2406; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2408 = 8'h13 == _GEN_105 ? phv_data_19 : _GEN_2407; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2409 = 8'h14 == _GEN_105 ? phv_data_20 : _GEN_2408; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2410 = 8'h15 == _GEN_105 ? phv_data_21 : _GEN_2409; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2411 = 8'h16 == _GEN_105 ? phv_data_22 : _GEN_2410; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2412 = 8'h17 == _GEN_105 ? phv_data_23 : _GEN_2411; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2413 = 8'h18 == _GEN_105 ? phv_data_24 : _GEN_2412; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2414 = 8'h19 == _GEN_105 ? phv_data_25 : _GEN_2413; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2415 = 8'h1a == _GEN_105 ? phv_data_26 : _GEN_2414; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2416 = 8'h1b == _GEN_105 ? phv_data_27 : _GEN_2415; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2417 = 8'h1c == _GEN_105 ? phv_data_28 : _GEN_2416; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2418 = 8'h1d == _GEN_105 ? phv_data_29 : _GEN_2417; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2419 = 8'h1e == _GEN_105 ? phv_data_30 : _GEN_2418; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2420 = 8'h1f == _GEN_105 ? phv_data_31 : _GEN_2419; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2421 = 8'h20 == _GEN_105 ? phv_data_32 : _GEN_2420; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2422 = 8'h21 == _GEN_105 ? phv_data_33 : _GEN_2421; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2423 = 8'h22 == _GEN_105 ? phv_data_34 : _GEN_2422; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2424 = 8'h23 == _GEN_105 ? phv_data_35 : _GEN_2423; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2425 = 8'h24 == _GEN_105 ? phv_data_36 : _GEN_2424; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2426 = 8'h25 == _GEN_105 ? phv_data_37 : _GEN_2425; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2427 = 8'h26 == _GEN_105 ? phv_data_38 : _GEN_2426; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2428 = 8'h27 == _GEN_105 ? phv_data_39 : _GEN_2427; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2429 = 8'h28 == _GEN_105 ? phv_data_40 : _GEN_2428; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2430 = 8'h29 == _GEN_105 ? phv_data_41 : _GEN_2429; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2431 = 8'h2a == _GEN_105 ? phv_data_42 : _GEN_2430; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2432 = 8'h2b == _GEN_105 ? phv_data_43 : _GEN_2431; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2433 = 8'h2c == _GEN_105 ? phv_data_44 : _GEN_2432; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2434 = 8'h2d == _GEN_105 ? phv_data_45 : _GEN_2433; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2435 = 8'h2e == _GEN_105 ? phv_data_46 : _GEN_2434; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2436 = 8'h2f == _GEN_105 ? phv_data_47 : _GEN_2435; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2437 = 8'h30 == _GEN_105 ? phv_data_48 : _GEN_2436; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2438 = 8'h31 == _GEN_105 ? phv_data_49 : _GEN_2437; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2439 = 8'h32 == _GEN_105 ? phv_data_50 : _GEN_2438; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2440 = 8'h33 == _GEN_105 ? phv_data_51 : _GEN_2439; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2441 = 8'h34 == _GEN_105 ? phv_data_52 : _GEN_2440; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2442 = 8'h35 == _GEN_105 ? phv_data_53 : _GEN_2441; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2443 = 8'h36 == _GEN_105 ? phv_data_54 : _GEN_2442; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2444 = 8'h37 == _GEN_105 ? phv_data_55 : _GEN_2443; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2445 = 8'h38 == _GEN_105 ? phv_data_56 : _GEN_2444; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2446 = 8'h39 == _GEN_105 ? phv_data_57 : _GEN_2445; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2447 = 8'h3a == _GEN_105 ? phv_data_58 : _GEN_2446; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2448 = 8'h3b == _GEN_105 ? phv_data_59 : _GEN_2447; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2449 = 8'h3c == _GEN_105 ? phv_data_60 : _GEN_2448; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2450 = 8'h3d == _GEN_105 ? phv_data_61 : _GEN_2449; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2451 = 8'h3e == _GEN_105 ? phv_data_62 : _GEN_2450; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2452 = 8'h3f == _GEN_105 ? phv_data_63 : _GEN_2451; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] bytes_4_3 = _GEN_81 ? _GEN_2452 : 8'h0; // @[matcher_pisa.scala 129:46 matcher_pisa.scala 128:34]
  wire [31:0] _groups_4_T = {bytes_4_0,bytes_4_1,bytes_4_2,bytes_4_3}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_2454 = _GEN_60 == 2'h1 ? _groups_4_T : 32'h0; // @[matcher_pisa.scala 123:50 matcher_pisa.scala 137:31 matcher_pisa.scala 122:27]
  wire [15:0] _GEN_2455 = 8'h40 == _GEN_102 ? _double_bytes_0_T : 16'h0; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53 matcher_pisa.scala 144:41]
  wire [15:0] _GEN_2456 = 8'h41 == _GEN_102 ? _double_bytes_0_T_1 : _GEN_2455; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2457 = 8'h42 == _GEN_102 ? _double_bytes_0_T_2 : _GEN_2456; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2458 = 8'h43 == _GEN_102 ? _double_bytes_0_T_3 : _GEN_2457; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2459 = 8'h44 == _GEN_102 ? _double_bytes_0_T_4 : _GEN_2458; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2460 = 8'h45 == _GEN_102 ? _double_bytes_0_T_5 : _GEN_2459; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2461 = 8'h46 == _GEN_102 ? _double_bytes_0_T_6 : _GEN_2460; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2462 = 8'h47 == _GEN_102 ? _double_bytes_0_T_7 : _GEN_2461; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2463 = 8'h48 == _GEN_102 ? _double_bytes_0_T_8 : _GEN_2462; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2464 = 8'h49 == _GEN_102 ? _double_bytes_0_T_9 : _GEN_2463; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2465 = 8'h4a == _GEN_102 ? _double_bytes_0_T_10 : _GEN_2464; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2466 = 8'h4b == _GEN_102 ? _double_bytes_0_T_11 : _GEN_2465; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2467 = 8'h4c == _GEN_102 ? _double_bytes_0_T_12 : _GEN_2466; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2468 = 8'h4d == _GEN_102 ? _double_bytes_0_T_13 : _GEN_2467; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2469 = 8'h4e == _GEN_102 ? _double_bytes_0_T_14 : _GEN_2468; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2470 = 8'h4f == _GEN_102 ? _double_bytes_0_T_15 : _GEN_2469; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2471 = 8'h50 == _GEN_102 ? _double_bytes_0_T_16 : _GEN_2470; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2472 = 8'h51 == _GEN_102 ? _double_bytes_0_T_17 : _GEN_2471; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2473 = 8'h52 == _GEN_102 ? _double_bytes_0_T_18 : _GEN_2472; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2474 = 8'h53 == _GEN_102 ? _double_bytes_0_T_19 : _GEN_2473; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2475 = 8'h54 == _GEN_102 ? _double_bytes_0_T_20 : _GEN_2474; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2476 = 8'h55 == _GEN_102 ? _double_bytes_0_T_21 : _GEN_2475; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2477 = 8'h56 == _GEN_102 ? _double_bytes_0_T_22 : _GEN_2476; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2478 = 8'h57 == _GEN_102 ? _double_bytes_0_T_23 : _GEN_2477; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2479 = 8'h58 == _GEN_102 ? _double_bytes_0_T_24 : _GEN_2478; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2480 = 8'h59 == _GEN_102 ? _double_bytes_0_T_25 : _GEN_2479; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2481 = 8'h5a == _GEN_102 ? _double_bytes_0_T_26 : _GEN_2480; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2482 = 8'h5b == _GEN_102 ? _double_bytes_0_T_27 : _GEN_2481; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2483 = 8'h5c == _GEN_102 ? _double_bytes_0_T_28 : _GEN_2482; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2484 = 8'h5d == _GEN_102 ? _double_bytes_0_T_29 : _GEN_2483; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2485 = 8'h5e == _GEN_102 ? _double_bytes_0_T_30 : _GEN_2484; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2486 = 8'h5f == _GEN_102 ? _double_bytes_0_T_31 : _GEN_2485; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2487 = 8'h60 == _GEN_102 ? _double_bytes_0_T_32 : _GEN_2486; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2488 = 8'h61 == _GEN_102 ? _double_bytes_0_T_33 : _GEN_2487; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2489 = 8'h62 == _GEN_102 ? _double_bytes_0_T_34 : _GEN_2488; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2490 = 8'h63 == _GEN_102 ? _double_bytes_0_T_35 : _GEN_2489; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2491 = 8'h64 == _GEN_102 ? _double_bytes_0_T_36 : _GEN_2490; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2492 = 8'h65 == _GEN_102 ? _double_bytes_0_T_37 : _GEN_2491; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2493 = 8'h66 == _GEN_102 ? _double_bytes_0_T_38 : _GEN_2492; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2494 = 8'h67 == _GEN_102 ? _double_bytes_0_T_39 : _GEN_2493; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2495 = 8'h68 == _GEN_102 ? _double_bytes_0_T_40 : _GEN_2494; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2496 = 8'h69 == _GEN_102 ? _double_bytes_0_T_41 : _GEN_2495; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2497 = 8'h6a == _GEN_102 ? _double_bytes_0_T_42 : _GEN_2496; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2498 = 8'h6b == _GEN_102 ? _double_bytes_0_T_43 : _GEN_2497; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2499 = 8'h6c == _GEN_102 ? _double_bytes_0_T_44 : _GEN_2498; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2500 = 8'h6d == _GEN_102 ? _double_bytes_0_T_45 : _GEN_2499; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2501 = 8'h6e == _GEN_102 ? _double_bytes_0_T_46 : _GEN_2500; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2502 = 8'h6f == _GEN_102 ? _double_bytes_0_T_47 : _GEN_2501; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2503 = 8'h70 == _GEN_102 ? _double_bytes_0_T_48 : _GEN_2502; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2504 = 8'h71 == _GEN_102 ? _double_bytes_0_T_49 : _GEN_2503; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2505 = 8'h72 == _GEN_102 ? _double_bytes_0_T_50 : _GEN_2504; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2506 = 8'h73 == _GEN_102 ? _double_bytes_0_T_51 : _GEN_2505; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2507 = 8'h74 == _GEN_102 ? _double_bytes_0_T_52 : _GEN_2506; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2508 = 8'h75 == _GEN_102 ? _double_bytes_0_T_53 : _GEN_2507; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2509 = 8'h76 == _GEN_102 ? _double_bytes_0_T_54 : _GEN_2508; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2510 = 8'h77 == _GEN_102 ? _double_bytes_0_T_55 : _GEN_2509; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2511 = 8'h78 == _GEN_102 ? _double_bytes_0_T_56 : _GEN_2510; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2512 = 8'h79 == _GEN_102 ? _double_bytes_0_T_57 : _GEN_2511; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2513 = 8'h7a == _GEN_102 ? _double_bytes_0_T_58 : _GEN_2512; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2514 = 8'h7b == _GEN_102 ? _double_bytes_0_T_59 : _GEN_2513; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2515 = 8'h7c == _GEN_102 ? _double_bytes_0_T_60 : _GEN_2514; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2516 = 8'h7d == _GEN_102 ? _double_bytes_0_T_61 : _GEN_2515; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2517 = 8'h7e == _GEN_102 ? _double_bytes_0_T_62 : _GEN_2516; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2518 = 8'h7f == _GEN_102 ? _double_bytes_0_T_63 : _GEN_2517; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2519 = 8'h80 == _GEN_102 ? _double_bytes_0_T_64 : _GEN_2518; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2520 = 8'h81 == _GEN_102 ? _double_bytes_0_T_65 : _GEN_2519; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2521 = 8'h82 == _GEN_102 ? _double_bytes_0_T_66 : _GEN_2520; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2522 = 8'h83 == _GEN_102 ? _double_bytes_0_T_67 : _GEN_2521; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2523 = 8'h84 == _GEN_102 ? _double_bytes_0_T_68 : _GEN_2522; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2524 = 8'h85 == _GEN_102 ? _double_bytes_0_T_69 : _GEN_2523; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2525 = 8'h86 == _GEN_102 ? _double_bytes_0_T_70 : _GEN_2524; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2526 = 8'h87 == _GEN_102 ? _double_bytes_0_T_71 : _GEN_2525; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2527 = 8'h88 == _GEN_102 ? _double_bytes_0_T_72 : _GEN_2526; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2528 = 8'h89 == _GEN_102 ? _double_bytes_0_T_73 : _GEN_2527; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2529 = 8'h8a == _GEN_102 ? _double_bytes_0_T_74 : _GEN_2528; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2530 = 8'h8b == _GEN_102 ? _double_bytes_0_T_75 : _GEN_2529; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2531 = 8'h8c == _GEN_102 ? _double_bytes_0_T_76 : _GEN_2530; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2532 = 8'h8d == _GEN_102 ? _double_bytes_0_T_77 : _GEN_2531; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2533 = 8'h8e == _GEN_102 ? _double_bytes_0_T_78 : _GEN_2532; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2534 = 8'h8f == _GEN_102 ? _double_bytes_0_T_79 : _GEN_2533; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2535 = 8'h90 == _GEN_102 ? _double_bytes_0_T_80 : _GEN_2534; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2536 = 8'h91 == _GEN_102 ? _double_bytes_0_T_81 : _GEN_2535; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2537 = 8'h92 == _GEN_102 ? _double_bytes_0_T_82 : _GEN_2536; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2538 = 8'h93 == _GEN_102 ? _double_bytes_0_T_83 : _GEN_2537; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2539 = 8'h94 == _GEN_102 ? _double_bytes_0_T_84 : _GEN_2538; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2540 = 8'h95 == _GEN_102 ? _double_bytes_0_T_85 : _GEN_2539; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2541 = 8'h96 == _GEN_102 ? _double_bytes_0_T_86 : _GEN_2540; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2542 = 8'h97 == _GEN_102 ? _double_bytes_0_T_87 : _GEN_2541; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2543 = 8'h98 == _GEN_102 ? _double_bytes_0_T_88 : _GEN_2542; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2544 = 8'h99 == _GEN_102 ? _double_bytes_0_T_89 : _GEN_2543; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2545 = 8'h9a == _GEN_102 ? _double_bytes_0_T_90 : _GEN_2544; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2546 = 8'h9b == _GEN_102 ? _double_bytes_0_T_91 : _GEN_2545; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2547 = 8'h9c == _GEN_102 ? _double_bytes_0_T_92 : _GEN_2546; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2548 = 8'h9d == _GEN_102 ? _double_bytes_0_T_93 : _GEN_2547; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2549 = 8'h9e == _GEN_102 ? _double_bytes_0_T_94 : _GEN_2548; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2550 = 8'h9f == _GEN_102 ? _double_bytes_0_T_95 : _GEN_2549; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] double_bytes_4_0 = _GEN_78 ? _GEN_2550 : 16'h0; // @[matcher_pisa.scala 145:46 matcher_pisa.scala 144:41]
  wire [15:0] _GEN_2552 = 8'h40 == _GEN_103 ? _double_bytes_0_T : 16'h0; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53 matcher_pisa.scala 144:41]
  wire [15:0] _GEN_2553 = 8'h41 == _GEN_103 ? _double_bytes_0_T_1 : _GEN_2552; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2554 = 8'h42 == _GEN_103 ? _double_bytes_0_T_2 : _GEN_2553; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2555 = 8'h43 == _GEN_103 ? _double_bytes_0_T_3 : _GEN_2554; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2556 = 8'h44 == _GEN_103 ? _double_bytes_0_T_4 : _GEN_2555; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2557 = 8'h45 == _GEN_103 ? _double_bytes_0_T_5 : _GEN_2556; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2558 = 8'h46 == _GEN_103 ? _double_bytes_0_T_6 : _GEN_2557; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2559 = 8'h47 == _GEN_103 ? _double_bytes_0_T_7 : _GEN_2558; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2560 = 8'h48 == _GEN_103 ? _double_bytes_0_T_8 : _GEN_2559; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2561 = 8'h49 == _GEN_103 ? _double_bytes_0_T_9 : _GEN_2560; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2562 = 8'h4a == _GEN_103 ? _double_bytes_0_T_10 : _GEN_2561; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2563 = 8'h4b == _GEN_103 ? _double_bytes_0_T_11 : _GEN_2562; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2564 = 8'h4c == _GEN_103 ? _double_bytes_0_T_12 : _GEN_2563; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2565 = 8'h4d == _GEN_103 ? _double_bytes_0_T_13 : _GEN_2564; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2566 = 8'h4e == _GEN_103 ? _double_bytes_0_T_14 : _GEN_2565; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2567 = 8'h4f == _GEN_103 ? _double_bytes_0_T_15 : _GEN_2566; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2568 = 8'h50 == _GEN_103 ? _double_bytes_0_T_16 : _GEN_2567; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2569 = 8'h51 == _GEN_103 ? _double_bytes_0_T_17 : _GEN_2568; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2570 = 8'h52 == _GEN_103 ? _double_bytes_0_T_18 : _GEN_2569; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2571 = 8'h53 == _GEN_103 ? _double_bytes_0_T_19 : _GEN_2570; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2572 = 8'h54 == _GEN_103 ? _double_bytes_0_T_20 : _GEN_2571; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2573 = 8'h55 == _GEN_103 ? _double_bytes_0_T_21 : _GEN_2572; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2574 = 8'h56 == _GEN_103 ? _double_bytes_0_T_22 : _GEN_2573; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2575 = 8'h57 == _GEN_103 ? _double_bytes_0_T_23 : _GEN_2574; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2576 = 8'h58 == _GEN_103 ? _double_bytes_0_T_24 : _GEN_2575; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2577 = 8'h59 == _GEN_103 ? _double_bytes_0_T_25 : _GEN_2576; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2578 = 8'h5a == _GEN_103 ? _double_bytes_0_T_26 : _GEN_2577; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2579 = 8'h5b == _GEN_103 ? _double_bytes_0_T_27 : _GEN_2578; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2580 = 8'h5c == _GEN_103 ? _double_bytes_0_T_28 : _GEN_2579; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2581 = 8'h5d == _GEN_103 ? _double_bytes_0_T_29 : _GEN_2580; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2582 = 8'h5e == _GEN_103 ? _double_bytes_0_T_30 : _GEN_2581; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2583 = 8'h5f == _GEN_103 ? _double_bytes_0_T_31 : _GEN_2582; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2584 = 8'h60 == _GEN_103 ? _double_bytes_0_T_32 : _GEN_2583; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2585 = 8'h61 == _GEN_103 ? _double_bytes_0_T_33 : _GEN_2584; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2586 = 8'h62 == _GEN_103 ? _double_bytes_0_T_34 : _GEN_2585; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2587 = 8'h63 == _GEN_103 ? _double_bytes_0_T_35 : _GEN_2586; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2588 = 8'h64 == _GEN_103 ? _double_bytes_0_T_36 : _GEN_2587; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2589 = 8'h65 == _GEN_103 ? _double_bytes_0_T_37 : _GEN_2588; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2590 = 8'h66 == _GEN_103 ? _double_bytes_0_T_38 : _GEN_2589; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2591 = 8'h67 == _GEN_103 ? _double_bytes_0_T_39 : _GEN_2590; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2592 = 8'h68 == _GEN_103 ? _double_bytes_0_T_40 : _GEN_2591; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2593 = 8'h69 == _GEN_103 ? _double_bytes_0_T_41 : _GEN_2592; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2594 = 8'h6a == _GEN_103 ? _double_bytes_0_T_42 : _GEN_2593; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2595 = 8'h6b == _GEN_103 ? _double_bytes_0_T_43 : _GEN_2594; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2596 = 8'h6c == _GEN_103 ? _double_bytes_0_T_44 : _GEN_2595; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2597 = 8'h6d == _GEN_103 ? _double_bytes_0_T_45 : _GEN_2596; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2598 = 8'h6e == _GEN_103 ? _double_bytes_0_T_46 : _GEN_2597; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2599 = 8'h6f == _GEN_103 ? _double_bytes_0_T_47 : _GEN_2598; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2600 = 8'h70 == _GEN_103 ? _double_bytes_0_T_48 : _GEN_2599; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2601 = 8'h71 == _GEN_103 ? _double_bytes_0_T_49 : _GEN_2600; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2602 = 8'h72 == _GEN_103 ? _double_bytes_0_T_50 : _GEN_2601; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2603 = 8'h73 == _GEN_103 ? _double_bytes_0_T_51 : _GEN_2602; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2604 = 8'h74 == _GEN_103 ? _double_bytes_0_T_52 : _GEN_2603; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2605 = 8'h75 == _GEN_103 ? _double_bytes_0_T_53 : _GEN_2604; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2606 = 8'h76 == _GEN_103 ? _double_bytes_0_T_54 : _GEN_2605; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2607 = 8'h77 == _GEN_103 ? _double_bytes_0_T_55 : _GEN_2606; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2608 = 8'h78 == _GEN_103 ? _double_bytes_0_T_56 : _GEN_2607; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2609 = 8'h79 == _GEN_103 ? _double_bytes_0_T_57 : _GEN_2608; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2610 = 8'h7a == _GEN_103 ? _double_bytes_0_T_58 : _GEN_2609; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2611 = 8'h7b == _GEN_103 ? _double_bytes_0_T_59 : _GEN_2610; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2612 = 8'h7c == _GEN_103 ? _double_bytes_0_T_60 : _GEN_2611; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2613 = 8'h7d == _GEN_103 ? _double_bytes_0_T_61 : _GEN_2612; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2614 = 8'h7e == _GEN_103 ? _double_bytes_0_T_62 : _GEN_2613; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2615 = 8'h7f == _GEN_103 ? _double_bytes_0_T_63 : _GEN_2614; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2616 = 8'h80 == _GEN_103 ? _double_bytes_0_T_64 : _GEN_2615; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2617 = 8'h81 == _GEN_103 ? _double_bytes_0_T_65 : _GEN_2616; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2618 = 8'h82 == _GEN_103 ? _double_bytes_0_T_66 : _GEN_2617; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2619 = 8'h83 == _GEN_103 ? _double_bytes_0_T_67 : _GEN_2618; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2620 = 8'h84 == _GEN_103 ? _double_bytes_0_T_68 : _GEN_2619; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2621 = 8'h85 == _GEN_103 ? _double_bytes_0_T_69 : _GEN_2620; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2622 = 8'h86 == _GEN_103 ? _double_bytes_0_T_70 : _GEN_2621; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2623 = 8'h87 == _GEN_103 ? _double_bytes_0_T_71 : _GEN_2622; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2624 = 8'h88 == _GEN_103 ? _double_bytes_0_T_72 : _GEN_2623; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2625 = 8'h89 == _GEN_103 ? _double_bytes_0_T_73 : _GEN_2624; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2626 = 8'h8a == _GEN_103 ? _double_bytes_0_T_74 : _GEN_2625; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2627 = 8'h8b == _GEN_103 ? _double_bytes_0_T_75 : _GEN_2626; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2628 = 8'h8c == _GEN_103 ? _double_bytes_0_T_76 : _GEN_2627; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2629 = 8'h8d == _GEN_103 ? _double_bytes_0_T_77 : _GEN_2628; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2630 = 8'h8e == _GEN_103 ? _double_bytes_0_T_78 : _GEN_2629; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2631 = 8'h8f == _GEN_103 ? _double_bytes_0_T_79 : _GEN_2630; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2632 = 8'h90 == _GEN_103 ? _double_bytes_0_T_80 : _GEN_2631; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2633 = 8'h91 == _GEN_103 ? _double_bytes_0_T_81 : _GEN_2632; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2634 = 8'h92 == _GEN_103 ? _double_bytes_0_T_82 : _GEN_2633; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2635 = 8'h93 == _GEN_103 ? _double_bytes_0_T_83 : _GEN_2634; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2636 = 8'h94 == _GEN_103 ? _double_bytes_0_T_84 : _GEN_2635; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2637 = 8'h95 == _GEN_103 ? _double_bytes_0_T_85 : _GEN_2636; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2638 = 8'h96 == _GEN_103 ? _double_bytes_0_T_86 : _GEN_2637; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2639 = 8'h97 == _GEN_103 ? _double_bytes_0_T_87 : _GEN_2638; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2640 = 8'h98 == _GEN_103 ? _double_bytes_0_T_88 : _GEN_2639; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2641 = 8'h99 == _GEN_103 ? _double_bytes_0_T_89 : _GEN_2640; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2642 = 8'h9a == _GEN_103 ? _double_bytes_0_T_90 : _GEN_2641; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2643 = 8'h9b == _GEN_103 ? _double_bytes_0_T_91 : _GEN_2642; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2644 = 8'h9c == _GEN_103 ? _double_bytes_0_T_92 : _GEN_2643; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2645 = 8'h9d == _GEN_103 ? _double_bytes_0_T_93 : _GEN_2644; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2646 = 8'h9e == _GEN_103 ? _double_bytes_0_T_94 : _GEN_2645; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2647 = 8'h9f == _GEN_103 ? _double_bytes_0_T_95 : _GEN_2646; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] double_bytes_4_1 = _GEN_79 ? _GEN_2647 : 16'h0; // @[matcher_pisa.scala 145:46 matcher_pisa.scala 144:41]
  wire [31:0] _groups_4_T_1 = {double_bytes_4_0,double_bytes_4_1}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_2649 = _GEN_60 == 2'h2 ? _groups_4_T_1 : _GEN_2454; // @[matcher_pisa.scala 139:50 matcher_pisa.scala 153:31]
  wire [31:0] _GEN_2650 = 8'ha0 == _GEN_102 ? _groups_0_T_2 : 32'h0; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39 matcher_pisa.scala 158:31]
  wire [31:0] _GEN_2651 = 8'ha1 == _GEN_102 ? _groups_0_T_3 : _GEN_2650; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2652 = 8'ha2 == _GEN_102 ? _groups_0_T_4 : _GEN_2651; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2653 = 8'ha3 == _GEN_102 ? _groups_0_T_5 : _GEN_2652; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2654 = 8'ha4 == _GEN_102 ? _groups_0_T_6 : _GEN_2653; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2655 = 8'ha5 == _GEN_102 ? _groups_0_T_7 : _GEN_2654; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2656 = 8'ha6 == _GEN_102 ? _groups_0_T_8 : _GEN_2655; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2657 = 8'ha7 == _GEN_102 ? _groups_0_T_9 : _GEN_2656; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2658 = 8'ha8 == _GEN_102 ? _groups_0_T_10 : _GEN_2657; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2659 = 8'ha9 == _GEN_102 ? _groups_0_T_11 : _GEN_2658; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2660 = 8'haa == _GEN_102 ? _groups_0_T_12 : _GEN_2659; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2661 = 8'hab == _GEN_102 ? _groups_0_T_13 : _GEN_2660; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2662 = 8'hac == _GEN_102 ? _groups_0_T_14 : _GEN_2661; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2663 = 8'had == _GEN_102 ? _groups_0_T_15 : _GEN_2662; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2664 = 8'hae == _GEN_102 ? _groups_0_T_16 : _GEN_2663; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2665 = 8'haf == _GEN_102 ? _groups_0_T_17 : _GEN_2664; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2666 = 8'hb0 == _GEN_102 ? _groups_0_T_18 : _GEN_2665; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2667 = 8'hb1 == _GEN_102 ? _groups_0_T_19 : _GEN_2666; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2668 = 8'hb2 == _GEN_102 ? _groups_0_T_20 : _GEN_2667; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2669 = 8'hb3 == _GEN_102 ? _groups_0_T_21 : _GEN_2668; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2670 = 8'hb4 == _GEN_102 ? _groups_0_T_22 : _GEN_2669; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2671 = 8'hb5 == _GEN_102 ? _groups_0_T_23 : _GEN_2670; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2672 = 8'hb6 == _GEN_102 ? _groups_0_T_24 : _GEN_2671; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2673 = 8'hb7 == _GEN_102 ? _groups_0_T_25 : _GEN_2672; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2674 = 8'hb8 == _GEN_102 ? _groups_0_T_26 : _GEN_2673; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2675 = 8'hb9 == _GEN_102 ? _groups_0_T_27 : _GEN_2674; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2676 = 8'hba == _GEN_102 ? _groups_0_T_28 : _GEN_2675; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2677 = 8'hbb == _GEN_102 ? _groups_0_T_29 : _GEN_2676; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2678 = 8'hbc == _GEN_102 ? _groups_0_T_30 : _GEN_2677; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2679 = 8'hbd == _GEN_102 ? _groups_0_T_31 : _GEN_2678; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2680 = 8'hbe == _GEN_102 ? _groups_0_T_32 : _GEN_2679; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2681 = 8'hbf == _GEN_102 ? _groups_0_T_33 : _GEN_2680; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2682 = 8'hc0 == _GEN_102 ? _groups_0_T_34 : _GEN_2681; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2683 = 8'hc1 == _GEN_102 ? _groups_0_T_35 : _GEN_2682; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2684 = 8'hc2 == _GEN_102 ? _groups_0_T_36 : _GEN_2683; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2685 = 8'hc3 == _GEN_102 ? _groups_0_T_37 : _GEN_2684; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2686 = 8'hc4 == _GEN_102 ? _groups_0_T_38 : _GEN_2685; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2687 = 8'hc5 == _GEN_102 ? _groups_0_T_39 : _GEN_2686; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2688 = 8'hc6 == _GEN_102 ? _groups_0_T_40 : _GEN_2687; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2689 = 8'hc7 == _GEN_102 ? _groups_0_T_41 : _GEN_2688; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2690 = 8'hc8 == _GEN_102 ? _groups_0_T_42 : _GEN_2689; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2691 = 8'hc9 == _GEN_102 ? _groups_0_T_43 : _GEN_2690; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2692 = 8'hca == _GEN_102 ? _groups_0_T_44 : _GEN_2691; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2693 = 8'hcb == _GEN_102 ? _groups_0_T_45 : _GEN_2692; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2694 = 8'hcc == _GEN_102 ? _groups_0_T_46 : _GEN_2693; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2695 = 8'hcd == _GEN_102 ? _groups_0_T_47 : _GEN_2694; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2696 = 8'hce == _GEN_102 ? _groups_0_T_48 : _GEN_2695; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2697 = 8'hcf == _GEN_102 ? _groups_0_T_49 : _GEN_2696; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2698 = 8'hd0 == _GEN_102 ? _groups_0_T_50 : _GEN_2697; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2699 = 8'hd1 == _GEN_102 ? _groups_0_T_51 : _GEN_2698; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2700 = 8'hd2 == _GEN_102 ? _groups_0_T_52 : _GEN_2699; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2701 = 8'hd3 == _GEN_102 ? _groups_0_T_53 : _GEN_2700; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2702 = 8'hd4 == _GEN_102 ? _groups_0_T_54 : _GEN_2701; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2703 = 8'hd5 == _GEN_102 ? _groups_0_T_55 : _GEN_2702; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2704 = 8'hd6 == _GEN_102 ? _groups_0_T_56 : _GEN_2703; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2705 = 8'hd7 == _GEN_102 ? _groups_0_T_57 : _GEN_2704; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2706 = 8'hd8 == _GEN_102 ? _groups_0_T_58 : _GEN_2705; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2707 = 8'hd9 == _GEN_102 ? _groups_0_T_59 : _GEN_2706; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2708 = 8'hda == _GEN_102 ? _groups_0_T_60 : _GEN_2707; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2709 = 8'hdb == _GEN_102 ? _groups_0_T_61 : _GEN_2708; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2710 = 8'hdc == _GEN_102 ? _groups_0_T_62 : _GEN_2709; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2711 = 8'hdd == _GEN_102 ? _groups_0_T_63 : _GEN_2710; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2712 = 8'hde == _GEN_102 ? _groups_0_T_64 : _GEN_2711; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_2713 = 8'hdf == _GEN_102 ? _groups_0_T_65 : _GEN_2712; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] groups_4 = _GEN_60 == 2'h3 ? _GEN_2713 : _GEN_2649; // @[matcher_pisa.scala 155:50]
  wire [7:0] _GEN_2715 = 8'h0 == _GEN_106 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_2716 = 8'h1 == _GEN_106 ? phv_data_1 : _GEN_2715; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2717 = 8'h2 == _GEN_106 ? phv_data_2 : _GEN_2716; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2718 = 8'h3 == _GEN_106 ? phv_data_3 : _GEN_2717; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2719 = 8'h4 == _GEN_106 ? phv_data_4 : _GEN_2718; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2720 = 8'h5 == _GEN_106 ? phv_data_5 : _GEN_2719; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2721 = 8'h6 == _GEN_106 ? phv_data_6 : _GEN_2720; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2722 = 8'h7 == _GEN_106 ? phv_data_7 : _GEN_2721; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2723 = 8'h8 == _GEN_106 ? phv_data_8 : _GEN_2722; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2724 = 8'h9 == _GEN_106 ? phv_data_9 : _GEN_2723; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2725 = 8'ha == _GEN_106 ? phv_data_10 : _GEN_2724; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2726 = 8'hb == _GEN_106 ? phv_data_11 : _GEN_2725; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2727 = 8'hc == _GEN_106 ? phv_data_12 : _GEN_2726; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2728 = 8'hd == _GEN_106 ? phv_data_13 : _GEN_2727; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2729 = 8'he == _GEN_106 ? phv_data_14 : _GEN_2728; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2730 = 8'hf == _GEN_106 ? phv_data_15 : _GEN_2729; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2731 = 8'h10 == _GEN_106 ? phv_data_16 : _GEN_2730; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2732 = 8'h11 == _GEN_106 ? phv_data_17 : _GEN_2731; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2733 = 8'h12 == _GEN_106 ? phv_data_18 : _GEN_2732; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2734 = 8'h13 == _GEN_106 ? phv_data_19 : _GEN_2733; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2735 = 8'h14 == _GEN_106 ? phv_data_20 : _GEN_2734; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2736 = 8'h15 == _GEN_106 ? phv_data_21 : _GEN_2735; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2737 = 8'h16 == _GEN_106 ? phv_data_22 : _GEN_2736; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2738 = 8'h17 == _GEN_106 ? phv_data_23 : _GEN_2737; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2739 = 8'h18 == _GEN_106 ? phv_data_24 : _GEN_2738; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2740 = 8'h19 == _GEN_106 ? phv_data_25 : _GEN_2739; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2741 = 8'h1a == _GEN_106 ? phv_data_26 : _GEN_2740; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2742 = 8'h1b == _GEN_106 ? phv_data_27 : _GEN_2741; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2743 = 8'h1c == _GEN_106 ? phv_data_28 : _GEN_2742; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2744 = 8'h1d == _GEN_106 ? phv_data_29 : _GEN_2743; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2745 = 8'h1e == _GEN_106 ? phv_data_30 : _GEN_2744; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2746 = 8'h1f == _GEN_106 ? phv_data_31 : _GEN_2745; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2747 = 8'h20 == _GEN_106 ? phv_data_32 : _GEN_2746; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2748 = 8'h21 == _GEN_106 ? phv_data_33 : _GEN_2747; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2749 = 8'h22 == _GEN_106 ? phv_data_34 : _GEN_2748; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2750 = 8'h23 == _GEN_106 ? phv_data_35 : _GEN_2749; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2751 = 8'h24 == _GEN_106 ? phv_data_36 : _GEN_2750; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2752 = 8'h25 == _GEN_106 ? phv_data_37 : _GEN_2751; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2753 = 8'h26 == _GEN_106 ? phv_data_38 : _GEN_2752; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2754 = 8'h27 == _GEN_106 ? phv_data_39 : _GEN_2753; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2755 = 8'h28 == _GEN_106 ? phv_data_40 : _GEN_2754; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2756 = 8'h29 == _GEN_106 ? phv_data_41 : _GEN_2755; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2757 = 8'h2a == _GEN_106 ? phv_data_42 : _GEN_2756; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2758 = 8'h2b == _GEN_106 ? phv_data_43 : _GEN_2757; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2759 = 8'h2c == _GEN_106 ? phv_data_44 : _GEN_2758; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2760 = 8'h2d == _GEN_106 ? phv_data_45 : _GEN_2759; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2761 = 8'h2e == _GEN_106 ? phv_data_46 : _GEN_2760; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2762 = 8'h2f == _GEN_106 ? phv_data_47 : _GEN_2761; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2763 = 8'h30 == _GEN_106 ? phv_data_48 : _GEN_2762; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2764 = 8'h31 == _GEN_106 ? phv_data_49 : _GEN_2763; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2765 = 8'h32 == _GEN_106 ? phv_data_50 : _GEN_2764; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2766 = 8'h33 == _GEN_106 ? phv_data_51 : _GEN_2765; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2767 = 8'h34 == _GEN_106 ? phv_data_52 : _GEN_2766; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2768 = 8'h35 == _GEN_106 ? phv_data_53 : _GEN_2767; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2769 = 8'h36 == _GEN_106 ? phv_data_54 : _GEN_2768; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2770 = 8'h37 == _GEN_106 ? phv_data_55 : _GEN_2769; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2771 = 8'h38 == _GEN_106 ? phv_data_56 : _GEN_2770; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2772 = 8'h39 == _GEN_106 ? phv_data_57 : _GEN_2771; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2773 = 8'h3a == _GEN_106 ? phv_data_58 : _GEN_2772; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2774 = 8'h3b == _GEN_106 ? phv_data_59 : _GEN_2773; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2775 = 8'h3c == _GEN_106 ? phv_data_60 : _GEN_2774; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2776 = 8'h3d == _GEN_106 ? phv_data_61 : _GEN_2775; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2777 = 8'h3e == _GEN_106 ? phv_data_62 : _GEN_2776; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2778 = 8'h3f == _GEN_106 ? phv_data_63 : _GEN_2777; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] bytes_5_0 = _GEN_82 ? _GEN_2778 : 8'h0; // @[matcher_pisa.scala 129:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_2780 = 8'h0 == _GEN_107 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_2781 = 8'h1 == _GEN_107 ? phv_data_1 : _GEN_2780; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2782 = 8'h2 == _GEN_107 ? phv_data_2 : _GEN_2781; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2783 = 8'h3 == _GEN_107 ? phv_data_3 : _GEN_2782; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2784 = 8'h4 == _GEN_107 ? phv_data_4 : _GEN_2783; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2785 = 8'h5 == _GEN_107 ? phv_data_5 : _GEN_2784; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2786 = 8'h6 == _GEN_107 ? phv_data_6 : _GEN_2785; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2787 = 8'h7 == _GEN_107 ? phv_data_7 : _GEN_2786; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2788 = 8'h8 == _GEN_107 ? phv_data_8 : _GEN_2787; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2789 = 8'h9 == _GEN_107 ? phv_data_9 : _GEN_2788; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2790 = 8'ha == _GEN_107 ? phv_data_10 : _GEN_2789; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2791 = 8'hb == _GEN_107 ? phv_data_11 : _GEN_2790; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2792 = 8'hc == _GEN_107 ? phv_data_12 : _GEN_2791; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2793 = 8'hd == _GEN_107 ? phv_data_13 : _GEN_2792; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2794 = 8'he == _GEN_107 ? phv_data_14 : _GEN_2793; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2795 = 8'hf == _GEN_107 ? phv_data_15 : _GEN_2794; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2796 = 8'h10 == _GEN_107 ? phv_data_16 : _GEN_2795; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2797 = 8'h11 == _GEN_107 ? phv_data_17 : _GEN_2796; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2798 = 8'h12 == _GEN_107 ? phv_data_18 : _GEN_2797; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2799 = 8'h13 == _GEN_107 ? phv_data_19 : _GEN_2798; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2800 = 8'h14 == _GEN_107 ? phv_data_20 : _GEN_2799; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2801 = 8'h15 == _GEN_107 ? phv_data_21 : _GEN_2800; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2802 = 8'h16 == _GEN_107 ? phv_data_22 : _GEN_2801; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2803 = 8'h17 == _GEN_107 ? phv_data_23 : _GEN_2802; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2804 = 8'h18 == _GEN_107 ? phv_data_24 : _GEN_2803; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2805 = 8'h19 == _GEN_107 ? phv_data_25 : _GEN_2804; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2806 = 8'h1a == _GEN_107 ? phv_data_26 : _GEN_2805; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2807 = 8'h1b == _GEN_107 ? phv_data_27 : _GEN_2806; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2808 = 8'h1c == _GEN_107 ? phv_data_28 : _GEN_2807; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2809 = 8'h1d == _GEN_107 ? phv_data_29 : _GEN_2808; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2810 = 8'h1e == _GEN_107 ? phv_data_30 : _GEN_2809; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2811 = 8'h1f == _GEN_107 ? phv_data_31 : _GEN_2810; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2812 = 8'h20 == _GEN_107 ? phv_data_32 : _GEN_2811; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2813 = 8'h21 == _GEN_107 ? phv_data_33 : _GEN_2812; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2814 = 8'h22 == _GEN_107 ? phv_data_34 : _GEN_2813; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2815 = 8'h23 == _GEN_107 ? phv_data_35 : _GEN_2814; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2816 = 8'h24 == _GEN_107 ? phv_data_36 : _GEN_2815; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2817 = 8'h25 == _GEN_107 ? phv_data_37 : _GEN_2816; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2818 = 8'h26 == _GEN_107 ? phv_data_38 : _GEN_2817; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2819 = 8'h27 == _GEN_107 ? phv_data_39 : _GEN_2818; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2820 = 8'h28 == _GEN_107 ? phv_data_40 : _GEN_2819; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2821 = 8'h29 == _GEN_107 ? phv_data_41 : _GEN_2820; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2822 = 8'h2a == _GEN_107 ? phv_data_42 : _GEN_2821; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2823 = 8'h2b == _GEN_107 ? phv_data_43 : _GEN_2822; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2824 = 8'h2c == _GEN_107 ? phv_data_44 : _GEN_2823; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2825 = 8'h2d == _GEN_107 ? phv_data_45 : _GEN_2824; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2826 = 8'h2e == _GEN_107 ? phv_data_46 : _GEN_2825; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2827 = 8'h2f == _GEN_107 ? phv_data_47 : _GEN_2826; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2828 = 8'h30 == _GEN_107 ? phv_data_48 : _GEN_2827; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2829 = 8'h31 == _GEN_107 ? phv_data_49 : _GEN_2828; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2830 = 8'h32 == _GEN_107 ? phv_data_50 : _GEN_2829; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2831 = 8'h33 == _GEN_107 ? phv_data_51 : _GEN_2830; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2832 = 8'h34 == _GEN_107 ? phv_data_52 : _GEN_2831; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2833 = 8'h35 == _GEN_107 ? phv_data_53 : _GEN_2832; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2834 = 8'h36 == _GEN_107 ? phv_data_54 : _GEN_2833; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2835 = 8'h37 == _GEN_107 ? phv_data_55 : _GEN_2834; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2836 = 8'h38 == _GEN_107 ? phv_data_56 : _GEN_2835; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2837 = 8'h39 == _GEN_107 ? phv_data_57 : _GEN_2836; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2838 = 8'h3a == _GEN_107 ? phv_data_58 : _GEN_2837; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2839 = 8'h3b == _GEN_107 ? phv_data_59 : _GEN_2838; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2840 = 8'h3c == _GEN_107 ? phv_data_60 : _GEN_2839; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2841 = 8'h3d == _GEN_107 ? phv_data_61 : _GEN_2840; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2842 = 8'h3e == _GEN_107 ? phv_data_62 : _GEN_2841; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2843 = 8'h3f == _GEN_107 ? phv_data_63 : _GEN_2842; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] bytes_5_1 = _GEN_83 ? _GEN_2843 : 8'h0; // @[matcher_pisa.scala 129:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_2845 = 8'h0 == _GEN_108 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_2846 = 8'h1 == _GEN_108 ? phv_data_1 : _GEN_2845; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2847 = 8'h2 == _GEN_108 ? phv_data_2 : _GEN_2846; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2848 = 8'h3 == _GEN_108 ? phv_data_3 : _GEN_2847; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2849 = 8'h4 == _GEN_108 ? phv_data_4 : _GEN_2848; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2850 = 8'h5 == _GEN_108 ? phv_data_5 : _GEN_2849; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2851 = 8'h6 == _GEN_108 ? phv_data_6 : _GEN_2850; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2852 = 8'h7 == _GEN_108 ? phv_data_7 : _GEN_2851; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2853 = 8'h8 == _GEN_108 ? phv_data_8 : _GEN_2852; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2854 = 8'h9 == _GEN_108 ? phv_data_9 : _GEN_2853; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2855 = 8'ha == _GEN_108 ? phv_data_10 : _GEN_2854; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2856 = 8'hb == _GEN_108 ? phv_data_11 : _GEN_2855; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2857 = 8'hc == _GEN_108 ? phv_data_12 : _GEN_2856; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2858 = 8'hd == _GEN_108 ? phv_data_13 : _GEN_2857; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2859 = 8'he == _GEN_108 ? phv_data_14 : _GEN_2858; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2860 = 8'hf == _GEN_108 ? phv_data_15 : _GEN_2859; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2861 = 8'h10 == _GEN_108 ? phv_data_16 : _GEN_2860; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2862 = 8'h11 == _GEN_108 ? phv_data_17 : _GEN_2861; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2863 = 8'h12 == _GEN_108 ? phv_data_18 : _GEN_2862; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2864 = 8'h13 == _GEN_108 ? phv_data_19 : _GEN_2863; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2865 = 8'h14 == _GEN_108 ? phv_data_20 : _GEN_2864; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2866 = 8'h15 == _GEN_108 ? phv_data_21 : _GEN_2865; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2867 = 8'h16 == _GEN_108 ? phv_data_22 : _GEN_2866; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2868 = 8'h17 == _GEN_108 ? phv_data_23 : _GEN_2867; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2869 = 8'h18 == _GEN_108 ? phv_data_24 : _GEN_2868; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2870 = 8'h19 == _GEN_108 ? phv_data_25 : _GEN_2869; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2871 = 8'h1a == _GEN_108 ? phv_data_26 : _GEN_2870; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2872 = 8'h1b == _GEN_108 ? phv_data_27 : _GEN_2871; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2873 = 8'h1c == _GEN_108 ? phv_data_28 : _GEN_2872; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2874 = 8'h1d == _GEN_108 ? phv_data_29 : _GEN_2873; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2875 = 8'h1e == _GEN_108 ? phv_data_30 : _GEN_2874; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2876 = 8'h1f == _GEN_108 ? phv_data_31 : _GEN_2875; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2877 = 8'h20 == _GEN_108 ? phv_data_32 : _GEN_2876; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2878 = 8'h21 == _GEN_108 ? phv_data_33 : _GEN_2877; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2879 = 8'h22 == _GEN_108 ? phv_data_34 : _GEN_2878; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2880 = 8'h23 == _GEN_108 ? phv_data_35 : _GEN_2879; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2881 = 8'h24 == _GEN_108 ? phv_data_36 : _GEN_2880; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2882 = 8'h25 == _GEN_108 ? phv_data_37 : _GEN_2881; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2883 = 8'h26 == _GEN_108 ? phv_data_38 : _GEN_2882; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2884 = 8'h27 == _GEN_108 ? phv_data_39 : _GEN_2883; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2885 = 8'h28 == _GEN_108 ? phv_data_40 : _GEN_2884; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2886 = 8'h29 == _GEN_108 ? phv_data_41 : _GEN_2885; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2887 = 8'h2a == _GEN_108 ? phv_data_42 : _GEN_2886; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2888 = 8'h2b == _GEN_108 ? phv_data_43 : _GEN_2887; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2889 = 8'h2c == _GEN_108 ? phv_data_44 : _GEN_2888; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2890 = 8'h2d == _GEN_108 ? phv_data_45 : _GEN_2889; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2891 = 8'h2e == _GEN_108 ? phv_data_46 : _GEN_2890; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2892 = 8'h2f == _GEN_108 ? phv_data_47 : _GEN_2891; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2893 = 8'h30 == _GEN_108 ? phv_data_48 : _GEN_2892; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2894 = 8'h31 == _GEN_108 ? phv_data_49 : _GEN_2893; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2895 = 8'h32 == _GEN_108 ? phv_data_50 : _GEN_2894; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2896 = 8'h33 == _GEN_108 ? phv_data_51 : _GEN_2895; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2897 = 8'h34 == _GEN_108 ? phv_data_52 : _GEN_2896; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2898 = 8'h35 == _GEN_108 ? phv_data_53 : _GEN_2897; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2899 = 8'h36 == _GEN_108 ? phv_data_54 : _GEN_2898; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2900 = 8'h37 == _GEN_108 ? phv_data_55 : _GEN_2899; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2901 = 8'h38 == _GEN_108 ? phv_data_56 : _GEN_2900; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2902 = 8'h39 == _GEN_108 ? phv_data_57 : _GEN_2901; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2903 = 8'h3a == _GEN_108 ? phv_data_58 : _GEN_2902; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2904 = 8'h3b == _GEN_108 ? phv_data_59 : _GEN_2903; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2905 = 8'h3c == _GEN_108 ? phv_data_60 : _GEN_2904; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2906 = 8'h3d == _GEN_108 ? phv_data_61 : _GEN_2905; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2907 = 8'h3e == _GEN_108 ? phv_data_62 : _GEN_2906; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2908 = 8'h3f == _GEN_108 ? phv_data_63 : _GEN_2907; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] bytes_5_2 = _GEN_84 ? _GEN_2908 : 8'h0; // @[matcher_pisa.scala 129:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_2910 = 8'h0 == _GEN_109 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_2911 = 8'h1 == _GEN_109 ? phv_data_1 : _GEN_2910; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2912 = 8'h2 == _GEN_109 ? phv_data_2 : _GEN_2911; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2913 = 8'h3 == _GEN_109 ? phv_data_3 : _GEN_2912; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2914 = 8'h4 == _GEN_109 ? phv_data_4 : _GEN_2913; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2915 = 8'h5 == _GEN_109 ? phv_data_5 : _GEN_2914; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2916 = 8'h6 == _GEN_109 ? phv_data_6 : _GEN_2915; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2917 = 8'h7 == _GEN_109 ? phv_data_7 : _GEN_2916; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2918 = 8'h8 == _GEN_109 ? phv_data_8 : _GEN_2917; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2919 = 8'h9 == _GEN_109 ? phv_data_9 : _GEN_2918; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2920 = 8'ha == _GEN_109 ? phv_data_10 : _GEN_2919; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2921 = 8'hb == _GEN_109 ? phv_data_11 : _GEN_2920; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2922 = 8'hc == _GEN_109 ? phv_data_12 : _GEN_2921; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2923 = 8'hd == _GEN_109 ? phv_data_13 : _GEN_2922; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2924 = 8'he == _GEN_109 ? phv_data_14 : _GEN_2923; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2925 = 8'hf == _GEN_109 ? phv_data_15 : _GEN_2924; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2926 = 8'h10 == _GEN_109 ? phv_data_16 : _GEN_2925; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2927 = 8'h11 == _GEN_109 ? phv_data_17 : _GEN_2926; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2928 = 8'h12 == _GEN_109 ? phv_data_18 : _GEN_2927; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2929 = 8'h13 == _GEN_109 ? phv_data_19 : _GEN_2928; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2930 = 8'h14 == _GEN_109 ? phv_data_20 : _GEN_2929; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2931 = 8'h15 == _GEN_109 ? phv_data_21 : _GEN_2930; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2932 = 8'h16 == _GEN_109 ? phv_data_22 : _GEN_2931; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2933 = 8'h17 == _GEN_109 ? phv_data_23 : _GEN_2932; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2934 = 8'h18 == _GEN_109 ? phv_data_24 : _GEN_2933; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2935 = 8'h19 == _GEN_109 ? phv_data_25 : _GEN_2934; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2936 = 8'h1a == _GEN_109 ? phv_data_26 : _GEN_2935; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2937 = 8'h1b == _GEN_109 ? phv_data_27 : _GEN_2936; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2938 = 8'h1c == _GEN_109 ? phv_data_28 : _GEN_2937; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2939 = 8'h1d == _GEN_109 ? phv_data_29 : _GEN_2938; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2940 = 8'h1e == _GEN_109 ? phv_data_30 : _GEN_2939; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2941 = 8'h1f == _GEN_109 ? phv_data_31 : _GEN_2940; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2942 = 8'h20 == _GEN_109 ? phv_data_32 : _GEN_2941; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2943 = 8'h21 == _GEN_109 ? phv_data_33 : _GEN_2942; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2944 = 8'h22 == _GEN_109 ? phv_data_34 : _GEN_2943; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2945 = 8'h23 == _GEN_109 ? phv_data_35 : _GEN_2944; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2946 = 8'h24 == _GEN_109 ? phv_data_36 : _GEN_2945; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2947 = 8'h25 == _GEN_109 ? phv_data_37 : _GEN_2946; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2948 = 8'h26 == _GEN_109 ? phv_data_38 : _GEN_2947; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2949 = 8'h27 == _GEN_109 ? phv_data_39 : _GEN_2948; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2950 = 8'h28 == _GEN_109 ? phv_data_40 : _GEN_2949; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2951 = 8'h29 == _GEN_109 ? phv_data_41 : _GEN_2950; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2952 = 8'h2a == _GEN_109 ? phv_data_42 : _GEN_2951; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2953 = 8'h2b == _GEN_109 ? phv_data_43 : _GEN_2952; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2954 = 8'h2c == _GEN_109 ? phv_data_44 : _GEN_2953; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2955 = 8'h2d == _GEN_109 ? phv_data_45 : _GEN_2954; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2956 = 8'h2e == _GEN_109 ? phv_data_46 : _GEN_2955; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2957 = 8'h2f == _GEN_109 ? phv_data_47 : _GEN_2956; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2958 = 8'h30 == _GEN_109 ? phv_data_48 : _GEN_2957; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2959 = 8'h31 == _GEN_109 ? phv_data_49 : _GEN_2958; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2960 = 8'h32 == _GEN_109 ? phv_data_50 : _GEN_2959; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2961 = 8'h33 == _GEN_109 ? phv_data_51 : _GEN_2960; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2962 = 8'h34 == _GEN_109 ? phv_data_52 : _GEN_2961; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2963 = 8'h35 == _GEN_109 ? phv_data_53 : _GEN_2962; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2964 = 8'h36 == _GEN_109 ? phv_data_54 : _GEN_2963; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2965 = 8'h37 == _GEN_109 ? phv_data_55 : _GEN_2964; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2966 = 8'h38 == _GEN_109 ? phv_data_56 : _GEN_2965; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2967 = 8'h39 == _GEN_109 ? phv_data_57 : _GEN_2966; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2968 = 8'h3a == _GEN_109 ? phv_data_58 : _GEN_2967; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2969 = 8'h3b == _GEN_109 ? phv_data_59 : _GEN_2968; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2970 = 8'h3c == _GEN_109 ? phv_data_60 : _GEN_2969; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2971 = 8'h3d == _GEN_109 ? phv_data_61 : _GEN_2970; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2972 = 8'h3e == _GEN_109 ? phv_data_62 : _GEN_2971; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_2973 = 8'h3f == _GEN_109 ? phv_data_63 : _GEN_2972; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] bytes_5_3 = _GEN_85 ? _GEN_2973 : 8'h0; // @[matcher_pisa.scala 129:46 matcher_pisa.scala 128:34]
  wire [31:0] _groups_5_T = {bytes_5_0,bytes_5_1,bytes_5_2,bytes_5_3}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_2975 = _GEN_61 == 2'h1 ? _groups_5_T : 32'h0; // @[matcher_pisa.scala 123:50 matcher_pisa.scala 137:31 matcher_pisa.scala 122:27]
  wire [15:0] _GEN_2976 = 8'h40 == _GEN_106 ? _double_bytes_0_T : 16'h0; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53 matcher_pisa.scala 144:41]
  wire [15:0] _GEN_2977 = 8'h41 == _GEN_106 ? _double_bytes_0_T_1 : _GEN_2976; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2978 = 8'h42 == _GEN_106 ? _double_bytes_0_T_2 : _GEN_2977; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2979 = 8'h43 == _GEN_106 ? _double_bytes_0_T_3 : _GEN_2978; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2980 = 8'h44 == _GEN_106 ? _double_bytes_0_T_4 : _GEN_2979; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2981 = 8'h45 == _GEN_106 ? _double_bytes_0_T_5 : _GEN_2980; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2982 = 8'h46 == _GEN_106 ? _double_bytes_0_T_6 : _GEN_2981; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2983 = 8'h47 == _GEN_106 ? _double_bytes_0_T_7 : _GEN_2982; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2984 = 8'h48 == _GEN_106 ? _double_bytes_0_T_8 : _GEN_2983; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2985 = 8'h49 == _GEN_106 ? _double_bytes_0_T_9 : _GEN_2984; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2986 = 8'h4a == _GEN_106 ? _double_bytes_0_T_10 : _GEN_2985; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2987 = 8'h4b == _GEN_106 ? _double_bytes_0_T_11 : _GEN_2986; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2988 = 8'h4c == _GEN_106 ? _double_bytes_0_T_12 : _GEN_2987; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2989 = 8'h4d == _GEN_106 ? _double_bytes_0_T_13 : _GEN_2988; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2990 = 8'h4e == _GEN_106 ? _double_bytes_0_T_14 : _GEN_2989; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2991 = 8'h4f == _GEN_106 ? _double_bytes_0_T_15 : _GEN_2990; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2992 = 8'h50 == _GEN_106 ? _double_bytes_0_T_16 : _GEN_2991; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2993 = 8'h51 == _GEN_106 ? _double_bytes_0_T_17 : _GEN_2992; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2994 = 8'h52 == _GEN_106 ? _double_bytes_0_T_18 : _GEN_2993; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2995 = 8'h53 == _GEN_106 ? _double_bytes_0_T_19 : _GEN_2994; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2996 = 8'h54 == _GEN_106 ? _double_bytes_0_T_20 : _GEN_2995; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2997 = 8'h55 == _GEN_106 ? _double_bytes_0_T_21 : _GEN_2996; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2998 = 8'h56 == _GEN_106 ? _double_bytes_0_T_22 : _GEN_2997; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_2999 = 8'h57 == _GEN_106 ? _double_bytes_0_T_23 : _GEN_2998; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3000 = 8'h58 == _GEN_106 ? _double_bytes_0_T_24 : _GEN_2999; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3001 = 8'h59 == _GEN_106 ? _double_bytes_0_T_25 : _GEN_3000; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3002 = 8'h5a == _GEN_106 ? _double_bytes_0_T_26 : _GEN_3001; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3003 = 8'h5b == _GEN_106 ? _double_bytes_0_T_27 : _GEN_3002; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3004 = 8'h5c == _GEN_106 ? _double_bytes_0_T_28 : _GEN_3003; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3005 = 8'h5d == _GEN_106 ? _double_bytes_0_T_29 : _GEN_3004; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3006 = 8'h5e == _GEN_106 ? _double_bytes_0_T_30 : _GEN_3005; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3007 = 8'h5f == _GEN_106 ? _double_bytes_0_T_31 : _GEN_3006; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3008 = 8'h60 == _GEN_106 ? _double_bytes_0_T_32 : _GEN_3007; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3009 = 8'h61 == _GEN_106 ? _double_bytes_0_T_33 : _GEN_3008; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3010 = 8'h62 == _GEN_106 ? _double_bytes_0_T_34 : _GEN_3009; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3011 = 8'h63 == _GEN_106 ? _double_bytes_0_T_35 : _GEN_3010; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3012 = 8'h64 == _GEN_106 ? _double_bytes_0_T_36 : _GEN_3011; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3013 = 8'h65 == _GEN_106 ? _double_bytes_0_T_37 : _GEN_3012; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3014 = 8'h66 == _GEN_106 ? _double_bytes_0_T_38 : _GEN_3013; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3015 = 8'h67 == _GEN_106 ? _double_bytes_0_T_39 : _GEN_3014; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3016 = 8'h68 == _GEN_106 ? _double_bytes_0_T_40 : _GEN_3015; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3017 = 8'h69 == _GEN_106 ? _double_bytes_0_T_41 : _GEN_3016; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3018 = 8'h6a == _GEN_106 ? _double_bytes_0_T_42 : _GEN_3017; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3019 = 8'h6b == _GEN_106 ? _double_bytes_0_T_43 : _GEN_3018; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3020 = 8'h6c == _GEN_106 ? _double_bytes_0_T_44 : _GEN_3019; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3021 = 8'h6d == _GEN_106 ? _double_bytes_0_T_45 : _GEN_3020; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3022 = 8'h6e == _GEN_106 ? _double_bytes_0_T_46 : _GEN_3021; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3023 = 8'h6f == _GEN_106 ? _double_bytes_0_T_47 : _GEN_3022; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3024 = 8'h70 == _GEN_106 ? _double_bytes_0_T_48 : _GEN_3023; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3025 = 8'h71 == _GEN_106 ? _double_bytes_0_T_49 : _GEN_3024; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3026 = 8'h72 == _GEN_106 ? _double_bytes_0_T_50 : _GEN_3025; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3027 = 8'h73 == _GEN_106 ? _double_bytes_0_T_51 : _GEN_3026; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3028 = 8'h74 == _GEN_106 ? _double_bytes_0_T_52 : _GEN_3027; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3029 = 8'h75 == _GEN_106 ? _double_bytes_0_T_53 : _GEN_3028; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3030 = 8'h76 == _GEN_106 ? _double_bytes_0_T_54 : _GEN_3029; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3031 = 8'h77 == _GEN_106 ? _double_bytes_0_T_55 : _GEN_3030; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3032 = 8'h78 == _GEN_106 ? _double_bytes_0_T_56 : _GEN_3031; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3033 = 8'h79 == _GEN_106 ? _double_bytes_0_T_57 : _GEN_3032; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3034 = 8'h7a == _GEN_106 ? _double_bytes_0_T_58 : _GEN_3033; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3035 = 8'h7b == _GEN_106 ? _double_bytes_0_T_59 : _GEN_3034; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3036 = 8'h7c == _GEN_106 ? _double_bytes_0_T_60 : _GEN_3035; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3037 = 8'h7d == _GEN_106 ? _double_bytes_0_T_61 : _GEN_3036; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3038 = 8'h7e == _GEN_106 ? _double_bytes_0_T_62 : _GEN_3037; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3039 = 8'h7f == _GEN_106 ? _double_bytes_0_T_63 : _GEN_3038; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3040 = 8'h80 == _GEN_106 ? _double_bytes_0_T_64 : _GEN_3039; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3041 = 8'h81 == _GEN_106 ? _double_bytes_0_T_65 : _GEN_3040; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3042 = 8'h82 == _GEN_106 ? _double_bytes_0_T_66 : _GEN_3041; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3043 = 8'h83 == _GEN_106 ? _double_bytes_0_T_67 : _GEN_3042; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3044 = 8'h84 == _GEN_106 ? _double_bytes_0_T_68 : _GEN_3043; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3045 = 8'h85 == _GEN_106 ? _double_bytes_0_T_69 : _GEN_3044; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3046 = 8'h86 == _GEN_106 ? _double_bytes_0_T_70 : _GEN_3045; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3047 = 8'h87 == _GEN_106 ? _double_bytes_0_T_71 : _GEN_3046; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3048 = 8'h88 == _GEN_106 ? _double_bytes_0_T_72 : _GEN_3047; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3049 = 8'h89 == _GEN_106 ? _double_bytes_0_T_73 : _GEN_3048; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3050 = 8'h8a == _GEN_106 ? _double_bytes_0_T_74 : _GEN_3049; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3051 = 8'h8b == _GEN_106 ? _double_bytes_0_T_75 : _GEN_3050; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3052 = 8'h8c == _GEN_106 ? _double_bytes_0_T_76 : _GEN_3051; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3053 = 8'h8d == _GEN_106 ? _double_bytes_0_T_77 : _GEN_3052; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3054 = 8'h8e == _GEN_106 ? _double_bytes_0_T_78 : _GEN_3053; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3055 = 8'h8f == _GEN_106 ? _double_bytes_0_T_79 : _GEN_3054; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3056 = 8'h90 == _GEN_106 ? _double_bytes_0_T_80 : _GEN_3055; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3057 = 8'h91 == _GEN_106 ? _double_bytes_0_T_81 : _GEN_3056; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3058 = 8'h92 == _GEN_106 ? _double_bytes_0_T_82 : _GEN_3057; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3059 = 8'h93 == _GEN_106 ? _double_bytes_0_T_83 : _GEN_3058; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3060 = 8'h94 == _GEN_106 ? _double_bytes_0_T_84 : _GEN_3059; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3061 = 8'h95 == _GEN_106 ? _double_bytes_0_T_85 : _GEN_3060; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3062 = 8'h96 == _GEN_106 ? _double_bytes_0_T_86 : _GEN_3061; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3063 = 8'h97 == _GEN_106 ? _double_bytes_0_T_87 : _GEN_3062; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3064 = 8'h98 == _GEN_106 ? _double_bytes_0_T_88 : _GEN_3063; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3065 = 8'h99 == _GEN_106 ? _double_bytes_0_T_89 : _GEN_3064; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3066 = 8'h9a == _GEN_106 ? _double_bytes_0_T_90 : _GEN_3065; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3067 = 8'h9b == _GEN_106 ? _double_bytes_0_T_91 : _GEN_3066; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3068 = 8'h9c == _GEN_106 ? _double_bytes_0_T_92 : _GEN_3067; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3069 = 8'h9d == _GEN_106 ? _double_bytes_0_T_93 : _GEN_3068; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3070 = 8'h9e == _GEN_106 ? _double_bytes_0_T_94 : _GEN_3069; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3071 = 8'h9f == _GEN_106 ? _double_bytes_0_T_95 : _GEN_3070; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] double_bytes_5_0 = _GEN_82 ? _GEN_3071 : 16'h0; // @[matcher_pisa.scala 145:46 matcher_pisa.scala 144:41]
  wire [15:0] _GEN_3073 = 8'h40 == _GEN_107 ? _double_bytes_0_T : 16'h0; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53 matcher_pisa.scala 144:41]
  wire [15:0] _GEN_3074 = 8'h41 == _GEN_107 ? _double_bytes_0_T_1 : _GEN_3073; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3075 = 8'h42 == _GEN_107 ? _double_bytes_0_T_2 : _GEN_3074; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3076 = 8'h43 == _GEN_107 ? _double_bytes_0_T_3 : _GEN_3075; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3077 = 8'h44 == _GEN_107 ? _double_bytes_0_T_4 : _GEN_3076; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3078 = 8'h45 == _GEN_107 ? _double_bytes_0_T_5 : _GEN_3077; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3079 = 8'h46 == _GEN_107 ? _double_bytes_0_T_6 : _GEN_3078; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3080 = 8'h47 == _GEN_107 ? _double_bytes_0_T_7 : _GEN_3079; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3081 = 8'h48 == _GEN_107 ? _double_bytes_0_T_8 : _GEN_3080; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3082 = 8'h49 == _GEN_107 ? _double_bytes_0_T_9 : _GEN_3081; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3083 = 8'h4a == _GEN_107 ? _double_bytes_0_T_10 : _GEN_3082; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3084 = 8'h4b == _GEN_107 ? _double_bytes_0_T_11 : _GEN_3083; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3085 = 8'h4c == _GEN_107 ? _double_bytes_0_T_12 : _GEN_3084; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3086 = 8'h4d == _GEN_107 ? _double_bytes_0_T_13 : _GEN_3085; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3087 = 8'h4e == _GEN_107 ? _double_bytes_0_T_14 : _GEN_3086; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3088 = 8'h4f == _GEN_107 ? _double_bytes_0_T_15 : _GEN_3087; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3089 = 8'h50 == _GEN_107 ? _double_bytes_0_T_16 : _GEN_3088; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3090 = 8'h51 == _GEN_107 ? _double_bytes_0_T_17 : _GEN_3089; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3091 = 8'h52 == _GEN_107 ? _double_bytes_0_T_18 : _GEN_3090; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3092 = 8'h53 == _GEN_107 ? _double_bytes_0_T_19 : _GEN_3091; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3093 = 8'h54 == _GEN_107 ? _double_bytes_0_T_20 : _GEN_3092; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3094 = 8'h55 == _GEN_107 ? _double_bytes_0_T_21 : _GEN_3093; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3095 = 8'h56 == _GEN_107 ? _double_bytes_0_T_22 : _GEN_3094; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3096 = 8'h57 == _GEN_107 ? _double_bytes_0_T_23 : _GEN_3095; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3097 = 8'h58 == _GEN_107 ? _double_bytes_0_T_24 : _GEN_3096; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3098 = 8'h59 == _GEN_107 ? _double_bytes_0_T_25 : _GEN_3097; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3099 = 8'h5a == _GEN_107 ? _double_bytes_0_T_26 : _GEN_3098; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3100 = 8'h5b == _GEN_107 ? _double_bytes_0_T_27 : _GEN_3099; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3101 = 8'h5c == _GEN_107 ? _double_bytes_0_T_28 : _GEN_3100; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3102 = 8'h5d == _GEN_107 ? _double_bytes_0_T_29 : _GEN_3101; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3103 = 8'h5e == _GEN_107 ? _double_bytes_0_T_30 : _GEN_3102; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3104 = 8'h5f == _GEN_107 ? _double_bytes_0_T_31 : _GEN_3103; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3105 = 8'h60 == _GEN_107 ? _double_bytes_0_T_32 : _GEN_3104; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3106 = 8'h61 == _GEN_107 ? _double_bytes_0_T_33 : _GEN_3105; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3107 = 8'h62 == _GEN_107 ? _double_bytes_0_T_34 : _GEN_3106; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3108 = 8'h63 == _GEN_107 ? _double_bytes_0_T_35 : _GEN_3107; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3109 = 8'h64 == _GEN_107 ? _double_bytes_0_T_36 : _GEN_3108; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3110 = 8'h65 == _GEN_107 ? _double_bytes_0_T_37 : _GEN_3109; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3111 = 8'h66 == _GEN_107 ? _double_bytes_0_T_38 : _GEN_3110; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3112 = 8'h67 == _GEN_107 ? _double_bytes_0_T_39 : _GEN_3111; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3113 = 8'h68 == _GEN_107 ? _double_bytes_0_T_40 : _GEN_3112; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3114 = 8'h69 == _GEN_107 ? _double_bytes_0_T_41 : _GEN_3113; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3115 = 8'h6a == _GEN_107 ? _double_bytes_0_T_42 : _GEN_3114; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3116 = 8'h6b == _GEN_107 ? _double_bytes_0_T_43 : _GEN_3115; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3117 = 8'h6c == _GEN_107 ? _double_bytes_0_T_44 : _GEN_3116; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3118 = 8'h6d == _GEN_107 ? _double_bytes_0_T_45 : _GEN_3117; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3119 = 8'h6e == _GEN_107 ? _double_bytes_0_T_46 : _GEN_3118; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3120 = 8'h6f == _GEN_107 ? _double_bytes_0_T_47 : _GEN_3119; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3121 = 8'h70 == _GEN_107 ? _double_bytes_0_T_48 : _GEN_3120; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3122 = 8'h71 == _GEN_107 ? _double_bytes_0_T_49 : _GEN_3121; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3123 = 8'h72 == _GEN_107 ? _double_bytes_0_T_50 : _GEN_3122; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3124 = 8'h73 == _GEN_107 ? _double_bytes_0_T_51 : _GEN_3123; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3125 = 8'h74 == _GEN_107 ? _double_bytes_0_T_52 : _GEN_3124; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3126 = 8'h75 == _GEN_107 ? _double_bytes_0_T_53 : _GEN_3125; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3127 = 8'h76 == _GEN_107 ? _double_bytes_0_T_54 : _GEN_3126; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3128 = 8'h77 == _GEN_107 ? _double_bytes_0_T_55 : _GEN_3127; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3129 = 8'h78 == _GEN_107 ? _double_bytes_0_T_56 : _GEN_3128; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3130 = 8'h79 == _GEN_107 ? _double_bytes_0_T_57 : _GEN_3129; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3131 = 8'h7a == _GEN_107 ? _double_bytes_0_T_58 : _GEN_3130; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3132 = 8'h7b == _GEN_107 ? _double_bytes_0_T_59 : _GEN_3131; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3133 = 8'h7c == _GEN_107 ? _double_bytes_0_T_60 : _GEN_3132; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3134 = 8'h7d == _GEN_107 ? _double_bytes_0_T_61 : _GEN_3133; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3135 = 8'h7e == _GEN_107 ? _double_bytes_0_T_62 : _GEN_3134; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3136 = 8'h7f == _GEN_107 ? _double_bytes_0_T_63 : _GEN_3135; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3137 = 8'h80 == _GEN_107 ? _double_bytes_0_T_64 : _GEN_3136; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3138 = 8'h81 == _GEN_107 ? _double_bytes_0_T_65 : _GEN_3137; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3139 = 8'h82 == _GEN_107 ? _double_bytes_0_T_66 : _GEN_3138; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3140 = 8'h83 == _GEN_107 ? _double_bytes_0_T_67 : _GEN_3139; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3141 = 8'h84 == _GEN_107 ? _double_bytes_0_T_68 : _GEN_3140; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3142 = 8'h85 == _GEN_107 ? _double_bytes_0_T_69 : _GEN_3141; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3143 = 8'h86 == _GEN_107 ? _double_bytes_0_T_70 : _GEN_3142; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3144 = 8'h87 == _GEN_107 ? _double_bytes_0_T_71 : _GEN_3143; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3145 = 8'h88 == _GEN_107 ? _double_bytes_0_T_72 : _GEN_3144; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3146 = 8'h89 == _GEN_107 ? _double_bytes_0_T_73 : _GEN_3145; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3147 = 8'h8a == _GEN_107 ? _double_bytes_0_T_74 : _GEN_3146; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3148 = 8'h8b == _GEN_107 ? _double_bytes_0_T_75 : _GEN_3147; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3149 = 8'h8c == _GEN_107 ? _double_bytes_0_T_76 : _GEN_3148; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3150 = 8'h8d == _GEN_107 ? _double_bytes_0_T_77 : _GEN_3149; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3151 = 8'h8e == _GEN_107 ? _double_bytes_0_T_78 : _GEN_3150; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3152 = 8'h8f == _GEN_107 ? _double_bytes_0_T_79 : _GEN_3151; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3153 = 8'h90 == _GEN_107 ? _double_bytes_0_T_80 : _GEN_3152; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3154 = 8'h91 == _GEN_107 ? _double_bytes_0_T_81 : _GEN_3153; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3155 = 8'h92 == _GEN_107 ? _double_bytes_0_T_82 : _GEN_3154; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3156 = 8'h93 == _GEN_107 ? _double_bytes_0_T_83 : _GEN_3155; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3157 = 8'h94 == _GEN_107 ? _double_bytes_0_T_84 : _GEN_3156; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3158 = 8'h95 == _GEN_107 ? _double_bytes_0_T_85 : _GEN_3157; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3159 = 8'h96 == _GEN_107 ? _double_bytes_0_T_86 : _GEN_3158; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3160 = 8'h97 == _GEN_107 ? _double_bytes_0_T_87 : _GEN_3159; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3161 = 8'h98 == _GEN_107 ? _double_bytes_0_T_88 : _GEN_3160; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3162 = 8'h99 == _GEN_107 ? _double_bytes_0_T_89 : _GEN_3161; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3163 = 8'h9a == _GEN_107 ? _double_bytes_0_T_90 : _GEN_3162; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3164 = 8'h9b == _GEN_107 ? _double_bytes_0_T_91 : _GEN_3163; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3165 = 8'h9c == _GEN_107 ? _double_bytes_0_T_92 : _GEN_3164; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3166 = 8'h9d == _GEN_107 ? _double_bytes_0_T_93 : _GEN_3165; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3167 = 8'h9e == _GEN_107 ? _double_bytes_0_T_94 : _GEN_3166; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_3168 = 8'h9f == _GEN_107 ? _double_bytes_0_T_95 : _GEN_3167; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] double_bytes_5_1 = _GEN_83 ? _GEN_3168 : 16'h0; // @[matcher_pisa.scala 145:46 matcher_pisa.scala 144:41]
  wire [31:0] _groups_5_T_1 = {double_bytes_5_0,double_bytes_5_1}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_3170 = _GEN_61 == 2'h2 ? _groups_5_T_1 : _GEN_2975; // @[matcher_pisa.scala 139:50 matcher_pisa.scala 153:31]
  wire [31:0] _GEN_3171 = 8'ha0 == _GEN_106 ? _groups_0_T_2 : 32'h0; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39 matcher_pisa.scala 158:31]
  wire [31:0] _GEN_3172 = 8'ha1 == _GEN_106 ? _groups_0_T_3 : _GEN_3171; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_3173 = 8'ha2 == _GEN_106 ? _groups_0_T_4 : _GEN_3172; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_3174 = 8'ha3 == _GEN_106 ? _groups_0_T_5 : _GEN_3173; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_3175 = 8'ha4 == _GEN_106 ? _groups_0_T_6 : _GEN_3174; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_3176 = 8'ha5 == _GEN_106 ? _groups_0_T_7 : _GEN_3175; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_3177 = 8'ha6 == _GEN_106 ? _groups_0_T_8 : _GEN_3176; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_3178 = 8'ha7 == _GEN_106 ? _groups_0_T_9 : _GEN_3177; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_3179 = 8'ha8 == _GEN_106 ? _groups_0_T_10 : _GEN_3178; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_3180 = 8'ha9 == _GEN_106 ? _groups_0_T_11 : _GEN_3179; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_3181 = 8'haa == _GEN_106 ? _groups_0_T_12 : _GEN_3180; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_3182 = 8'hab == _GEN_106 ? _groups_0_T_13 : _GEN_3181; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_3183 = 8'hac == _GEN_106 ? _groups_0_T_14 : _GEN_3182; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_3184 = 8'had == _GEN_106 ? _groups_0_T_15 : _GEN_3183; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_3185 = 8'hae == _GEN_106 ? _groups_0_T_16 : _GEN_3184; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_3186 = 8'haf == _GEN_106 ? _groups_0_T_17 : _GEN_3185; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_3187 = 8'hb0 == _GEN_106 ? _groups_0_T_18 : _GEN_3186; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_3188 = 8'hb1 == _GEN_106 ? _groups_0_T_19 : _GEN_3187; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_3189 = 8'hb2 == _GEN_106 ? _groups_0_T_20 : _GEN_3188; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_3190 = 8'hb3 == _GEN_106 ? _groups_0_T_21 : _GEN_3189; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_3191 = 8'hb4 == _GEN_106 ? _groups_0_T_22 : _GEN_3190; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_3192 = 8'hb5 == _GEN_106 ? _groups_0_T_23 : _GEN_3191; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_3193 = 8'hb6 == _GEN_106 ? _groups_0_T_24 : _GEN_3192; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_3194 = 8'hb7 == _GEN_106 ? _groups_0_T_25 : _GEN_3193; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_3195 = 8'hb8 == _GEN_106 ? _groups_0_T_26 : _GEN_3194; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_3196 = 8'hb9 == _GEN_106 ? _groups_0_T_27 : _GEN_3195; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_3197 = 8'hba == _GEN_106 ? _groups_0_T_28 : _GEN_3196; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_3198 = 8'hbb == _GEN_106 ? _groups_0_T_29 : _GEN_3197; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_3199 = 8'hbc == _GEN_106 ? _groups_0_T_30 : _GEN_3198; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_3200 = 8'hbd == _GEN_106 ? _groups_0_T_31 : _GEN_3199; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_3201 = 8'hbe == _GEN_106 ? _groups_0_T_32 : _GEN_3200; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_3202 = 8'hbf == _GEN_106 ? _groups_0_T_33 : _GEN_3201; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_3203 = 8'hc0 == _GEN_106 ? _groups_0_T_34 : _GEN_3202; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_3204 = 8'hc1 == _GEN_106 ? _groups_0_T_35 : _GEN_3203; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_3205 = 8'hc2 == _GEN_106 ? _groups_0_T_36 : _GEN_3204; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_3206 = 8'hc3 == _GEN_106 ? _groups_0_T_37 : _GEN_3205; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_3207 = 8'hc4 == _GEN_106 ? _groups_0_T_38 : _GEN_3206; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_3208 = 8'hc5 == _GEN_106 ? _groups_0_T_39 : _GEN_3207; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_3209 = 8'hc6 == _GEN_106 ? _groups_0_T_40 : _GEN_3208; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_3210 = 8'hc7 == _GEN_106 ? _groups_0_T_41 : _GEN_3209; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_3211 = 8'hc8 == _GEN_106 ? _groups_0_T_42 : _GEN_3210; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_3212 = 8'hc9 == _GEN_106 ? _groups_0_T_43 : _GEN_3211; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_3213 = 8'hca == _GEN_106 ? _groups_0_T_44 : _GEN_3212; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_3214 = 8'hcb == _GEN_106 ? _groups_0_T_45 : _GEN_3213; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_3215 = 8'hcc == _GEN_106 ? _groups_0_T_46 : _GEN_3214; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_3216 = 8'hcd == _GEN_106 ? _groups_0_T_47 : _GEN_3215; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_3217 = 8'hce == _GEN_106 ? _groups_0_T_48 : _GEN_3216; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_3218 = 8'hcf == _GEN_106 ? _groups_0_T_49 : _GEN_3217; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_3219 = 8'hd0 == _GEN_106 ? _groups_0_T_50 : _GEN_3218; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_3220 = 8'hd1 == _GEN_106 ? _groups_0_T_51 : _GEN_3219; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_3221 = 8'hd2 == _GEN_106 ? _groups_0_T_52 : _GEN_3220; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_3222 = 8'hd3 == _GEN_106 ? _groups_0_T_53 : _GEN_3221; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_3223 = 8'hd4 == _GEN_106 ? _groups_0_T_54 : _GEN_3222; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_3224 = 8'hd5 == _GEN_106 ? _groups_0_T_55 : _GEN_3223; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_3225 = 8'hd6 == _GEN_106 ? _groups_0_T_56 : _GEN_3224; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_3226 = 8'hd7 == _GEN_106 ? _groups_0_T_57 : _GEN_3225; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_3227 = 8'hd8 == _GEN_106 ? _groups_0_T_58 : _GEN_3226; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_3228 = 8'hd9 == _GEN_106 ? _groups_0_T_59 : _GEN_3227; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_3229 = 8'hda == _GEN_106 ? _groups_0_T_60 : _GEN_3228; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_3230 = 8'hdb == _GEN_106 ? _groups_0_T_61 : _GEN_3229; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_3231 = 8'hdc == _GEN_106 ? _groups_0_T_62 : _GEN_3230; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_3232 = 8'hdd == _GEN_106 ? _groups_0_T_63 : _GEN_3231; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_3233 = 8'hde == _GEN_106 ? _groups_0_T_64 : _GEN_3232; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_3234 = 8'hdf == _GEN_106 ? _groups_0_T_65 : _GEN_3233; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] groups_5 = _GEN_61 == 2'h3 ? _GEN_3234 : _GEN_3170; // @[matcher_pisa.scala 155:50]
  wire [191:0] _io_match_key_T = {groups_0,groups_1,groups_2,groups_3,groups_4,groups_5}; // @[Cat.scala 30:58]
  assign io_pipe_phv_out_data_0 = phv_data_0; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_1 = phv_data_1; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_2 = phv_data_2; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_3 = phv_data_3; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_4 = phv_data_4; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_5 = phv_data_5; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_6 = phv_data_6; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_7 = phv_data_7; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_8 = phv_data_8; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_9 = phv_data_9; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_10 = phv_data_10; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_11 = phv_data_11; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_12 = phv_data_12; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_13 = phv_data_13; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_14 = phv_data_14; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_15 = phv_data_15; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_16 = phv_data_16; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_17 = phv_data_17; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_18 = phv_data_18; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_19 = phv_data_19; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_20 = phv_data_20; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_21 = phv_data_21; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_22 = phv_data_22; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_23 = phv_data_23; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_24 = phv_data_24; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_25 = phv_data_25; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_26 = phv_data_26; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_27 = phv_data_27; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_28 = phv_data_28; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_29 = phv_data_29; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_30 = phv_data_30; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_31 = phv_data_31; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_32 = phv_data_32; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_33 = phv_data_33; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_34 = phv_data_34; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_35 = phv_data_35; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_36 = phv_data_36; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_37 = phv_data_37; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_38 = phv_data_38; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_39 = phv_data_39; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_40 = phv_data_40; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_41 = phv_data_41; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_42 = phv_data_42; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_43 = phv_data_43; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_44 = phv_data_44; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_45 = phv_data_45; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_46 = phv_data_46; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_47 = phv_data_47; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_48 = phv_data_48; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_49 = phv_data_49; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_50 = phv_data_50; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_51 = phv_data_51; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_52 = phv_data_52; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_53 = phv_data_53; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_54 = phv_data_54; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_55 = phv_data_55; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_56 = phv_data_56; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_57 = phv_data_57; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_58 = phv_data_58; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_59 = phv_data_59; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_60 = phv_data_60; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_61 = phv_data_61; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_62 = phv_data_62; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_63 = phv_data_63; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_64 = phv_data_64; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_65 = phv_data_65; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_66 = phv_data_66; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_67 = phv_data_67; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_68 = phv_data_68; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_69 = phv_data_69; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_70 = phv_data_70; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_71 = phv_data_71; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_72 = phv_data_72; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_73 = phv_data_73; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_74 = phv_data_74; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_75 = phv_data_75; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_76 = phv_data_76; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_77 = phv_data_77; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_78 = phv_data_78; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_79 = phv_data_79; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_80 = phv_data_80; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_81 = phv_data_81; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_82 = phv_data_82; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_83 = phv_data_83; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_84 = phv_data_84; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_85 = phv_data_85; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_86 = phv_data_86; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_87 = phv_data_87; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_88 = phv_data_88; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_89 = phv_data_89; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_90 = phv_data_90; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_91 = phv_data_91; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_92 = phv_data_92; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_93 = phv_data_93; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_94 = phv_data_94; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_95 = phv_data_95; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_96 = phv_data_96; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_97 = phv_data_97; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_98 = phv_data_98; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_99 = phv_data_99; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_100 = phv_data_100; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_101 = phv_data_101; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_102 = phv_data_102; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_103 = phv_data_103; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_104 = phv_data_104; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_105 = phv_data_105; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_106 = phv_data_106; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_107 = phv_data_107; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_108 = phv_data_108; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_109 = phv_data_109; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_110 = phv_data_110; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_111 = phv_data_111; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_112 = phv_data_112; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_113 = phv_data_113; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_114 = phv_data_114; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_115 = phv_data_115; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_116 = phv_data_116; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_117 = phv_data_117; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_118 = phv_data_118; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_119 = phv_data_119; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_120 = phv_data_120; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_121 = phv_data_121; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_122 = phv_data_122; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_123 = phv_data_123; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_124 = phv_data_124; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_125 = phv_data_125; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_126 = phv_data_126; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_127 = phv_data_127; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_128 = phv_data_128; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_129 = phv_data_129; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_130 = phv_data_130; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_131 = phv_data_131; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_132 = phv_data_132; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_133 = phv_data_133; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_134 = phv_data_134; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_135 = phv_data_135; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_136 = phv_data_136; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_137 = phv_data_137; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_138 = phv_data_138; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_139 = phv_data_139; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_140 = phv_data_140; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_141 = phv_data_141; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_142 = phv_data_142; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_143 = phv_data_143; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_144 = phv_data_144; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_145 = phv_data_145; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_146 = phv_data_146; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_147 = phv_data_147; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_148 = phv_data_148; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_149 = phv_data_149; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_150 = phv_data_150; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_151 = phv_data_151; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_152 = phv_data_152; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_153 = phv_data_153; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_154 = phv_data_154; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_155 = phv_data_155; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_156 = phv_data_156; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_157 = phv_data_157; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_158 = phv_data_158; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_159 = phv_data_159; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_160 = phv_data_160; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_161 = phv_data_161; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_162 = phv_data_162; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_163 = phv_data_163; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_164 = phv_data_164; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_165 = phv_data_165; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_166 = phv_data_166; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_167 = phv_data_167; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_168 = phv_data_168; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_169 = phv_data_169; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_170 = phv_data_170; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_171 = phv_data_171; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_172 = phv_data_172; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_173 = phv_data_173; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_174 = phv_data_174; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_175 = phv_data_175; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_176 = phv_data_176; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_177 = phv_data_177; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_178 = phv_data_178; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_179 = phv_data_179; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_180 = phv_data_180; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_181 = phv_data_181; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_182 = phv_data_182; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_183 = phv_data_183; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_184 = phv_data_184; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_185 = phv_data_185; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_186 = phv_data_186; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_187 = phv_data_187; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_188 = phv_data_188; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_189 = phv_data_189; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_190 = phv_data_190; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_191 = phv_data_191; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_192 = phv_data_192; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_193 = phv_data_193; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_194 = phv_data_194; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_195 = phv_data_195; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_196 = phv_data_196; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_197 = phv_data_197; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_198 = phv_data_198; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_199 = phv_data_199; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_200 = phv_data_200; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_201 = phv_data_201; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_202 = phv_data_202; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_203 = phv_data_203; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_204 = phv_data_204; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_205 = phv_data_205; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_206 = phv_data_206; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_207 = phv_data_207; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_208 = phv_data_208; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_209 = phv_data_209; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_210 = phv_data_210; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_211 = phv_data_211; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_212 = phv_data_212; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_213 = phv_data_213; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_214 = phv_data_214; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_215 = phv_data_215; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_216 = phv_data_216; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_217 = phv_data_217; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_218 = phv_data_218; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_219 = phv_data_219; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_220 = phv_data_220; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_221 = phv_data_221; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_222 = phv_data_222; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_223 = phv_data_223; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_224 = phv_data_224; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_225 = phv_data_225; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_226 = phv_data_226; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_227 = phv_data_227; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_228 = phv_data_228; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_229 = phv_data_229; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_230 = phv_data_230; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_231 = phv_data_231; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_232 = phv_data_232; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_233 = phv_data_233; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_234 = phv_data_234; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_235 = phv_data_235; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_236 = phv_data_236; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_237 = phv_data_237; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_238 = phv_data_238; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_239 = phv_data_239; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_240 = phv_data_240; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_241 = phv_data_241; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_242 = phv_data_242; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_243 = phv_data_243; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_244 = phv_data_244; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_245 = phv_data_245; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_246 = phv_data_246; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_247 = phv_data_247; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_248 = phv_data_248; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_249 = phv_data_249; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_250 = phv_data_250; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_251 = phv_data_251; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_252 = phv_data_252; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_253 = phv_data_253; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_254 = phv_data_254; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_255 = phv_data_255; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_256 = phv_data_256; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_257 = phv_data_257; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_258 = phv_data_258; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_259 = phv_data_259; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_260 = phv_data_260; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_261 = phv_data_261; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_262 = phv_data_262; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_263 = phv_data_263; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_264 = phv_data_264; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_265 = phv_data_265; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_266 = phv_data_266; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_267 = phv_data_267; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_268 = phv_data_268; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_269 = phv_data_269; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_270 = phv_data_270; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_271 = phv_data_271; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_272 = phv_data_272; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_273 = phv_data_273; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_274 = phv_data_274; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_275 = phv_data_275; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_276 = phv_data_276; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_277 = phv_data_277; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_278 = phv_data_278; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_279 = phv_data_279; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_280 = phv_data_280; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_281 = phv_data_281; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_282 = phv_data_282; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_283 = phv_data_283; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_284 = phv_data_284; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_285 = phv_data_285; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_286 = phv_data_286; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_287 = phv_data_287; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_288 = phv_data_288; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_289 = phv_data_289; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_290 = phv_data_290; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_291 = phv_data_291; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_292 = phv_data_292; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_293 = phv_data_293; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_294 = phv_data_294; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_295 = phv_data_295; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_296 = phv_data_296; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_297 = phv_data_297; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_298 = phv_data_298; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_299 = phv_data_299; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_300 = phv_data_300; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_301 = phv_data_301; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_302 = phv_data_302; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_303 = phv_data_303; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_304 = phv_data_304; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_305 = phv_data_305; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_306 = phv_data_306; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_307 = phv_data_307; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_308 = phv_data_308; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_309 = phv_data_309; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_310 = phv_data_310; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_311 = phv_data_311; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_312 = phv_data_312; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_313 = phv_data_313; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_314 = phv_data_314; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_315 = phv_data_315; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_316 = phv_data_316; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_317 = phv_data_317; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_318 = phv_data_318; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_319 = phv_data_319; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_320 = phv_data_320; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_321 = phv_data_321; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_322 = phv_data_322; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_323 = phv_data_323; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_324 = phv_data_324; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_325 = phv_data_325; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_326 = phv_data_326; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_327 = phv_data_327; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_328 = phv_data_328; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_329 = phv_data_329; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_330 = phv_data_330; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_331 = phv_data_331; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_332 = phv_data_332; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_333 = phv_data_333; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_334 = phv_data_334; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_335 = phv_data_335; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_336 = phv_data_336; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_337 = phv_data_337; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_338 = phv_data_338; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_339 = phv_data_339; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_340 = phv_data_340; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_341 = phv_data_341; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_342 = phv_data_342; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_343 = phv_data_343; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_344 = phv_data_344; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_345 = phv_data_345; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_346 = phv_data_346; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_347 = phv_data_347; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_348 = phv_data_348; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_349 = phv_data_349; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_350 = phv_data_350; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_351 = phv_data_351; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_352 = phv_data_352; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_353 = phv_data_353; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_354 = phv_data_354; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_355 = phv_data_355; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_356 = phv_data_356; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_357 = phv_data_357; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_358 = phv_data_358; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_359 = phv_data_359; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_360 = phv_data_360; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_361 = phv_data_361; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_362 = phv_data_362; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_363 = phv_data_363; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_364 = phv_data_364; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_365 = phv_data_365; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_366 = phv_data_366; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_367 = phv_data_367; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_368 = phv_data_368; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_369 = phv_data_369; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_370 = phv_data_370; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_371 = phv_data_371; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_372 = phv_data_372; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_373 = phv_data_373; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_374 = phv_data_374; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_375 = phv_data_375; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_376 = phv_data_376; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_377 = phv_data_377; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_378 = phv_data_378; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_379 = phv_data_379; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_380 = phv_data_380; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_381 = phv_data_381; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_382 = phv_data_382; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_383 = phv_data_383; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_384 = phv_data_384; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_385 = phv_data_385; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_386 = phv_data_386; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_387 = phv_data_387; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_388 = phv_data_388; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_389 = phv_data_389; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_390 = phv_data_390; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_391 = phv_data_391; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_392 = phv_data_392; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_393 = phv_data_393; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_394 = phv_data_394; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_395 = phv_data_395; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_396 = phv_data_396; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_397 = phv_data_397; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_398 = phv_data_398; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_399 = phv_data_399; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_400 = phv_data_400; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_401 = phv_data_401; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_402 = phv_data_402; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_403 = phv_data_403; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_404 = phv_data_404; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_405 = phv_data_405; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_406 = phv_data_406; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_407 = phv_data_407; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_408 = phv_data_408; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_409 = phv_data_409; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_410 = phv_data_410; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_411 = phv_data_411; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_412 = phv_data_412; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_413 = phv_data_413; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_414 = phv_data_414; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_415 = phv_data_415; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_416 = phv_data_416; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_417 = phv_data_417; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_418 = phv_data_418; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_419 = phv_data_419; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_420 = phv_data_420; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_421 = phv_data_421; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_422 = phv_data_422; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_423 = phv_data_423; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_424 = phv_data_424; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_425 = phv_data_425; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_426 = phv_data_426; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_427 = phv_data_427; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_428 = phv_data_428; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_429 = phv_data_429; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_430 = phv_data_430; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_431 = phv_data_431; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_432 = phv_data_432; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_433 = phv_data_433; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_434 = phv_data_434; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_435 = phv_data_435; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_436 = phv_data_436; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_437 = phv_data_437; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_438 = phv_data_438; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_439 = phv_data_439; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_440 = phv_data_440; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_441 = phv_data_441; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_442 = phv_data_442; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_443 = phv_data_443; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_444 = phv_data_444; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_445 = phv_data_445; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_446 = phv_data_446; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_447 = phv_data_447; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_448 = phv_data_448; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_449 = phv_data_449; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_450 = phv_data_450; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_451 = phv_data_451; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_452 = phv_data_452; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_453 = phv_data_453; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_454 = phv_data_454; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_455 = phv_data_455; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_456 = phv_data_456; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_457 = phv_data_457; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_458 = phv_data_458; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_459 = phv_data_459; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_460 = phv_data_460; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_461 = phv_data_461; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_462 = phv_data_462; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_463 = phv_data_463; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_464 = phv_data_464; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_465 = phv_data_465; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_466 = phv_data_466; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_467 = phv_data_467; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_468 = phv_data_468; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_469 = phv_data_469; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_470 = phv_data_470; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_471 = phv_data_471; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_472 = phv_data_472; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_473 = phv_data_473; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_474 = phv_data_474; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_475 = phv_data_475; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_476 = phv_data_476; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_477 = phv_data_477; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_478 = phv_data_478; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_479 = phv_data_479; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_480 = phv_data_480; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_481 = phv_data_481; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_482 = phv_data_482; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_483 = phv_data_483; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_484 = phv_data_484; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_485 = phv_data_485; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_486 = phv_data_486; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_487 = phv_data_487; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_488 = phv_data_488; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_489 = phv_data_489; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_490 = phv_data_490; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_491 = phv_data_491; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_492 = phv_data_492; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_493 = phv_data_493; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_494 = phv_data_494; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_495 = phv_data_495; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_496 = phv_data_496; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_497 = phv_data_497; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_498 = phv_data_498; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_499 = phv_data_499; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_500 = phv_data_500; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_501 = phv_data_501; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_502 = phv_data_502; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_503 = phv_data_503; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_504 = phv_data_504; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_505 = phv_data_505; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_506 = phv_data_506; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_507 = phv_data_507; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_508 = phv_data_508; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_509 = phv_data_509; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_510 = phv_data_510; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_511 = phv_data_511; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_next_processor_id = phv_next_processor_id; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_next_config_id = phv_next_config_id; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_is_valid_processor = phv_is_valid_processor; // @[matcher_pisa.scala 112:25]
  assign io_match_key = phv_is_valid_processor ? _io_match_key_T : 192'h0; // @[matcher_pisa.scala 116:39 matcher_pisa.scala 166:26 matcher_pisa.scala 168:26]
  always @(posedge clock) begin
    phv_data_0 <= io_pipe_phv_in_data_0; // @[matcher_pisa.scala 111:13]
    phv_data_1 <= io_pipe_phv_in_data_1; // @[matcher_pisa.scala 111:13]
    phv_data_2 <= io_pipe_phv_in_data_2; // @[matcher_pisa.scala 111:13]
    phv_data_3 <= io_pipe_phv_in_data_3; // @[matcher_pisa.scala 111:13]
    phv_data_4 <= io_pipe_phv_in_data_4; // @[matcher_pisa.scala 111:13]
    phv_data_5 <= io_pipe_phv_in_data_5; // @[matcher_pisa.scala 111:13]
    phv_data_6 <= io_pipe_phv_in_data_6; // @[matcher_pisa.scala 111:13]
    phv_data_7 <= io_pipe_phv_in_data_7; // @[matcher_pisa.scala 111:13]
    phv_data_8 <= io_pipe_phv_in_data_8; // @[matcher_pisa.scala 111:13]
    phv_data_9 <= io_pipe_phv_in_data_9; // @[matcher_pisa.scala 111:13]
    phv_data_10 <= io_pipe_phv_in_data_10; // @[matcher_pisa.scala 111:13]
    phv_data_11 <= io_pipe_phv_in_data_11; // @[matcher_pisa.scala 111:13]
    phv_data_12 <= io_pipe_phv_in_data_12; // @[matcher_pisa.scala 111:13]
    phv_data_13 <= io_pipe_phv_in_data_13; // @[matcher_pisa.scala 111:13]
    phv_data_14 <= io_pipe_phv_in_data_14; // @[matcher_pisa.scala 111:13]
    phv_data_15 <= io_pipe_phv_in_data_15; // @[matcher_pisa.scala 111:13]
    phv_data_16 <= io_pipe_phv_in_data_16; // @[matcher_pisa.scala 111:13]
    phv_data_17 <= io_pipe_phv_in_data_17; // @[matcher_pisa.scala 111:13]
    phv_data_18 <= io_pipe_phv_in_data_18; // @[matcher_pisa.scala 111:13]
    phv_data_19 <= io_pipe_phv_in_data_19; // @[matcher_pisa.scala 111:13]
    phv_data_20 <= io_pipe_phv_in_data_20; // @[matcher_pisa.scala 111:13]
    phv_data_21 <= io_pipe_phv_in_data_21; // @[matcher_pisa.scala 111:13]
    phv_data_22 <= io_pipe_phv_in_data_22; // @[matcher_pisa.scala 111:13]
    phv_data_23 <= io_pipe_phv_in_data_23; // @[matcher_pisa.scala 111:13]
    phv_data_24 <= io_pipe_phv_in_data_24; // @[matcher_pisa.scala 111:13]
    phv_data_25 <= io_pipe_phv_in_data_25; // @[matcher_pisa.scala 111:13]
    phv_data_26 <= io_pipe_phv_in_data_26; // @[matcher_pisa.scala 111:13]
    phv_data_27 <= io_pipe_phv_in_data_27; // @[matcher_pisa.scala 111:13]
    phv_data_28 <= io_pipe_phv_in_data_28; // @[matcher_pisa.scala 111:13]
    phv_data_29 <= io_pipe_phv_in_data_29; // @[matcher_pisa.scala 111:13]
    phv_data_30 <= io_pipe_phv_in_data_30; // @[matcher_pisa.scala 111:13]
    phv_data_31 <= io_pipe_phv_in_data_31; // @[matcher_pisa.scala 111:13]
    phv_data_32 <= io_pipe_phv_in_data_32; // @[matcher_pisa.scala 111:13]
    phv_data_33 <= io_pipe_phv_in_data_33; // @[matcher_pisa.scala 111:13]
    phv_data_34 <= io_pipe_phv_in_data_34; // @[matcher_pisa.scala 111:13]
    phv_data_35 <= io_pipe_phv_in_data_35; // @[matcher_pisa.scala 111:13]
    phv_data_36 <= io_pipe_phv_in_data_36; // @[matcher_pisa.scala 111:13]
    phv_data_37 <= io_pipe_phv_in_data_37; // @[matcher_pisa.scala 111:13]
    phv_data_38 <= io_pipe_phv_in_data_38; // @[matcher_pisa.scala 111:13]
    phv_data_39 <= io_pipe_phv_in_data_39; // @[matcher_pisa.scala 111:13]
    phv_data_40 <= io_pipe_phv_in_data_40; // @[matcher_pisa.scala 111:13]
    phv_data_41 <= io_pipe_phv_in_data_41; // @[matcher_pisa.scala 111:13]
    phv_data_42 <= io_pipe_phv_in_data_42; // @[matcher_pisa.scala 111:13]
    phv_data_43 <= io_pipe_phv_in_data_43; // @[matcher_pisa.scala 111:13]
    phv_data_44 <= io_pipe_phv_in_data_44; // @[matcher_pisa.scala 111:13]
    phv_data_45 <= io_pipe_phv_in_data_45; // @[matcher_pisa.scala 111:13]
    phv_data_46 <= io_pipe_phv_in_data_46; // @[matcher_pisa.scala 111:13]
    phv_data_47 <= io_pipe_phv_in_data_47; // @[matcher_pisa.scala 111:13]
    phv_data_48 <= io_pipe_phv_in_data_48; // @[matcher_pisa.scala 111:13]
    phv_data_49 <= io_pipe_phv_in_data_49; // @[matcher_pisa.scala 111:13]
    phv_data_50 <= io_pipe_phv_in_data_50; // @[matcher_pisa.scala 111:13]
    phv_data_51 <= io_pipe_phv_in_data_51; // @[matcher_pisa.scala 111:13]
    phv_data_52 <= io_pipe_phv_in_data_52; // @[matcher_pisa.scala 111:13]
    phv_data_53 <= io_pipe_phv_in_data_53; // @[matcher_pisa.scala 111:13]
    phv_data_54 <= io_pipe_phv_in_data_54; // @[matcher_pisa.scala 111:13]
    phv_data_55 <= io_pipe_phv_in_data_55; // @[matcher_pisa.scala 111:13]
    phv_data_56 <= io_pipe_phv_in_data_56; // @[matcher_pisa.scala 111:13]
    phv_data_57 <= io_pipe_phv_in_data_57; // @[matcher_pisa.scala 111:13]
    phv_data_58 <= io_pipe_phv_in_data_58; // @[matcher_pisa.scala 111:13]
    phv_data_59 <= io_pipe_phv_in_data_59; // @[matcher_pisa.scala 111:13]
    phv_data_60 <= io_pipe_phv_in_data_60; // @[matcher_pisa.scala 111:13]
    phv_data_61 <= io_pipe_phv_in_data_61; // @[matcher_pisa.scala 111:13]
    phv_data_62 <= io_pipe_phv_in_data_62; // @[matcher_pisa.scala 111:13]
    phv_data_63 <= io_pipe_phv_in_data_63; // @[matcher_pisa.scala 111:13]
    phv_data_64 <= io_pipe_phv_in_data_64; // @[matcher_pisa.scala 111:13]
    phv_data_65 <= io_pipe_phv_in_data_65; // @[matcher_pisa.scala 111:13]
    phv_data_66 <= io_pipe_phv_in_data_66; // @[matcher_pisa.scala 111:13]
    phv_data_67 <= io_pipe_phv_in_data_67; // @[matcher_pisa.scala 111:13]
    phv_data_68 <= io_pipe_phv_in_data_68; // @[matcher_pisa.scala 111:13]
    phv_data_69 <= io_pipe_phv_in_data_69; // @[matcher_pisa.scala 111:13]
    phv_data_70 <= io_pipe_phv_in_data_70; // @[matcher_pisa.scala 111:13]
    phv_data_71 <= io_pipe_phv_in_data_71; // @[matcher_pisa.scala 111:13]
    phv_data_72 <= io_pipe_phv_in_data_72; // @[matcher_pisa.scala 111:13]
    phv_data_73 <= io_pipe_phv_in_data_73; // @[matcher_pisa.scala 111:13]
    phv_data_74 <= io_pipe_phv_in_data_74; // @[matcher_pisa.scala 111:13]
    phv_data_75 <= io_pipe_phv_in_data_75; // @[matcher_pisa.scala 111:13]
    phv_data_76 <= io_pipe_phv_in_data_76; // @[matcher_pisa.scala 111:13]
    phv_data_77 <= io_pipe_phv_in_data_77; // @[matcher_pisa.scala 111:13]
    phv_data_78 <= io_pipe_phv_in_data_78; // @[matcher_pisa.scala 111:13]
    phv_data_79 <= io_pipe_phv_in_data_79; // @[matcher_pisa.scala 111:13]
    phv_data_80 <= io_pipe_phv_in_data_80; // @[matcher_pisa.scala 111:13]
    phv_data_81 <= io_pipe_phv_in_data_81; // @[matcher_pisa.scala 111:13]
    phv_data_82 <= io_pipe_phv_in_data_82; // @[matcher_pisa.scala 111:13]
    phv_data_83 <= io_pipe_phv_in_data_83; // @[matcher_pisa.scala 111:13]
    phv_data_84 <= io_pipe_phv_in_data_84; // @[matcher_pisa.scala 111:13]
    phv_data_85 <= io_pipe_phv_in_data_85; // @[matcher_pisa.scala 111:13]
    phv_data_86 <= io_pipe_phv_in_data_86; // @[matcher_pisa.scala 111:13]
    phv_data_87 <= io_pipe_phv_in_data_87; // @[matcher_pisa.scala 111:13]
    phv_data_88 <= io_pipe_phv_in_data_88; // @[matcher_pisa.scala 111:13]
    phv_data_89 <= io_pipe_phv_in_data_89; // @[matcher_pisa.scala 111:13]
    phv_data_90 <= io_pipe_phv_in_data_90; // @[matcher_pisa.scala 111:13]
    phv_data_91 <= io_pipe_phv_in_data_91; // @[matcher_pisa.scala 111:13]
    phv_data_92 <= io_pipe_phv_in_data_92; // @[matcher_pisa.scala 111:13]
    phv_data_93 <= io_pipe_phv_in_data_93; // @[matcher_pisa.scala 111:13]
    phv_data_94 <= io_pipe_phv_in_data_94; // @[matcher_pisa.scala 111:13]
    phv_data_95 <= io_pipe_phv_in_data_95; // @[matcher_pisa.scala 111:13]
    phv_data_96 <= io_pipe_phv_in_data_96; // @[matcher_pisa.scala 111:13]
    phv_data_97 <= io_pipe_phv_in_data_97; // @[matcher_pisa.scala 111:13]
    phv_data_98 <= io_pipe_phv_in_data_98; // @[matcher_pisa.scala 111:13]
    phv_data_99 <= io_pipe_phv_in_data_99; // @[matcher_pisa.scala 111:13]
    phv_data_100 <= io_pipe_phv_in_data_100; // @[matcher_pisa.scala 111:13]
    phv_data_101 <= io_pipe_phv_in_data_101; // @[matcher_pisa.scala 111:13]
    phv_data_102 <= io_pipe_phv_in_data_102; // @[matcher_pisa.scala 111:13]
    phv_data_103 <= io_pipe_phv_in_data_103; // @[matcher_pisa.scala 111:13]
    phv_data_104 <= io_pipe_phv_in_data_104; // @[matcher_pisa.scala 111:13]
    phv_data_105 <= io_pipe_phv_in_data_105; // @[matcher_pisa.scala 111:13]
    phv_data_106 <= io_pipe_phv_in_data_106; // @[matcher_pisa.scala 111:13]
    phv_data_107 <= io_pipe_phv_in_data_107; // @[matcher_pisa.scala 111:13]
    phv_data_108 <= io_pipe_phv_in_data_108; // @[matcher_pisa.scala 111:13]
    phv_data_109 <= io_pipe_phv_in_data_109; // @[matcher_pisa.scala 111:13]
    phv_data_110 <= io_pipe_phv_in_data_110; // @[matcher_pisa.scala 111:13]
    phv_data_111 <= io_pipe_phv_in_data_111; // @[matcher_pisa.scala 111:13]
    phv_data_112 <= io_pipe_phv_in_data_112; // @[matcher_pisa.scala 111:13]
    phv_data_113 <= io_pipe_phv_in_data_113; // @[matcher_pisa.scala 111:13]
    phv_data_114 <= io_pipe_phv_in_data_114; // @[matcher_pisa.scala 111:13]
    phv_data_115 <= io_pipe_phv_in_data_115; // @[matcher_pisa.scala 111:13]
    phv_data_116 <= io_pipe_phv_in_data_116; // @[matcher_pisa.scala 111:13]
    phv_data_117 <= io_pipe_phv_in_data_117; // @[matcher_pisa.scala 111:13]
    phv_data_118 <= io_pipe_phv_in_data_118; // @[matcher_pisa.scala 111:13]
    phv_data_119 <= io_pipe_phv_in_data_119; // @[matcher_pisa.scala 111:13]
    phv_data_120 <= io_pipe_phv_in_data_120; // @[matcher_pisa.scala 111:13]
    phv_data_121 <= io_pipe_phv_in_data_121; // @[matcher_pisa.scala 111:13]
    phv_data_122 <= io_pipe_phv_in_data_122; // @[matcher_pisa.scala 111:13]
    phv_data_123 <= io_pipe_phv_in_data_123; // @[matcher_pisa.scala 111:13]
    phv_data_124 <= io_pipe_phv_in_data_124; // @[matcher_pisa.scala 111:13]
    phv_data_125 <= io_pipe_phv_in_data_125; // @[matcher_pisa.scala 111:13]
    phv_data_126 <= io_pipe_phv_in_data_126; // @[matcher_pisa.scala 111:13]
    phv_data_127 <= io_pipe_phv_in_data_127; // @[matcher_pisa.scala 111:13]
    phv_data_128 <= io_pipe_phv_in_data_128; // @[matcher_pisa.scala 111:13]
    phv_data_129 <= io_pipe_phv_in_data_129; // @[matcher_pisa.scala 111:13]
    phv_data_130 <= io_pipe_phv_in_data_130; // @[matcher_pisa.scala 111:13]
    phv_data_131 <= io_pipe_phv_in_data_131; // @[matcher_pisa.scala 111:13]
    phv_data_132 <= io_pipe_phv_in_data_132; // @[matcher_pisa.scala 111:13]
    phv_data_133 <= io_pipe_phv_in_data_133; // @[matcher_pisa.scala 111:13]
    phv_data_134 <= io_pipe_phv_in_data_134; // @[matcher_pisa.scala 111:13]
    phv_data_135 <= io_pipe_phv_in_data_135; // @[matcher_pisa.scala 111:13]
    phv_data_136 <= io_pipe_phv_in_data_136; // @[matcher_pisa.scala 111:13]
    phv_data_137 <= io_pipe_phv_in_data_137; // @[matcher_pisa.scala 111:13]
    phv_data_138 <= io_pipe_phv_in_data_138; // @[matcher_pisa.scala 111:13]
    phv_data_139 <= io_pipe_phv_in_data_139; // @[matcher_pisa.scala 111:13]
    phv_data_140 <= io_pipe_phv_in_data_140; // @[matcher_pisa.scala 111:13]
    phv_data_141 <= io_pipe_phv_in_data_141; // @[matcher_pisa.scala 111:13]
    phv_data_142 <= io_pipe_phv_in_data_142; // @[matcher_pisa.scala 111:13]
    phv_data_143 <= io_pipe_phv_in_data_143; // @[matcher_pisa.scala 111:13]
    phv_data_144 <= io_pipe_phv_in_data_144; // @[matcher_pisa.scala 111:13]
    phv_data_145 <= io_pipe_phv_in_data_145; // @[matcher_pisa.scala 111:13]
    phv_data_146 <= io_pipe_phv_in_data_146; // @[matcher_pisa.scala 111:13]
    phv_data_147 <= io_pipe_phv_in_data_147; // @[matcher_pisa.scala 111:13]
    phv_data_148 <= io_pipe_phv_in_data_148; // @[matcher_pisa.scala 111:13]
    phv_data_149 <= io_pipe_phv_in_data_149; // @[matcher_pisa.scala 111:13]
    phv_data_150 <= io_pipe_phv_in_data_150; // @[matcher_pisa.scala 111:13]
    phv_data_151 <= io_pipe_phv_in_data_151; // @[matcher_pisa.scala 111:13]
    phv_data_152 <= io_pipe_phv_in_data_152; // @[matcher_pisa.scala 111:13]
    phv_data_153 <= io_pipe_phv_in_data_153; // @[matcher_pisa.scala 111:13]
    phv_data_154 <= io_pipe_phv_in_data_154; // @[matcher_pisa.scala 111:13]
    phv_data_155 <= io_pipe_phv_in_data_155; // @[matcher_pisa.scala 111:13]
    phv_data_156 <= io_pipe_phv_in_data_156; // @[matcher_pisa.scala 111:13]
    phv_data_157 <= io_pipe_phv_in_data_157; // @[matcher_pisa.scala 111:13]
    phv_data_158 <= io_pipe_phv_in_data_158; // @[matcher_pisa.scala 111:13]
    phv_data_159 <= io_pipe_phv_in_data_159; // @[matcher_pisa.scala 111:13]
    phv_data_160 <= io_pipe_phv_in_data_160; // @[matcher_pisa.scala 111:13]
    phv_data_161 <= io_pipe_phv_in_data_161; // @[matcher_pisa.scala 111:13]
    phv_data_162 <= io_pipe_phv_in_data_162; // @[matcher_pisa.scala 111:13]
    phv_data_163 <= io_pipe_phv_in_data_163; // @[matcher_pisa.scala 111:13]
    phv_data_164 <= io_pipe_phv_in_data_164; // @[matcher_pisa.scala 111:13]
    phv_data_165 <= io_pipe_phv_in_data_165; // @[matcher_pisa.scala 111:13]
    phv_data_166 <= io_pipe_phv_in_data_166; // @[matcher_pisa.scala 111:13]
    phv_data_167 <= io_pipe_phv_in_data_167; // @[matcher_pisa.scala 111:13]
    phv_data_168 <= io_pipe_phv_in_data_168; // @[matcher_pisa.scala 111:13]
    phv_data_169 <= io_pipe_phv_in_data_169; // @[matcher_pisa.scala 111:13]
    phv_data_170 <= io_pipe_phv_in_data_170; // @[matcher_pisa.scala 111:13]
    phv_data_171 <= io_pipe_phv_in_data_171; // @[matcher_pisa.scala 111:13]
    phv_data_172 <= io_pipe_phv_in_data_172; // @[matcher_pisa.scala 111:13]
    phv_data_173 <= io_pipe_phv_in_data_173; // @[matcher_pisa.scala 111:13]
    phv_data_174 <= io_pipe_phv_in_data_174; // @[matcher_pisa.scala 111:13]
    phv_data_175 <= io_pipe_phv_in_data_175; // @[matcher_pisa.scala 111:13]
    phv_data_176 <= io_pipe_phv_in_data_176; // @[matcher_pisa.scala 111:13]
    phv_data_177 <= io_pipe_phv_in_data_177; // @[matcher_pisa.scala 111:13]
    phv_data_178 <= io_pipe_phv_in_data_178; // @[matcher_pisa.scala 111:13]
    phv_data_179 <= io_pipe_phv_in_data_179; // @[matcher_pisa.scala 111:13]
    phv_data_180 <= io_pipe_phv_in_data_180; // @[matcher_pisa.scala 111:13]
    phv_data_181 <= io_pipe_phv_in_data_181; // @[matcher_pisa.scala 111:13]
    phv_data_182 <= io_pipe_phv_in_data_182; // @[matcher_pisa.scala 111:13]
    phv_data_183 <= io_pipe_phv_in_data_183; // @[matcher_pisa.scala 111:13]
    phv_data_184 <= io_pipe_phv_in_data_184; // @[matcher_pisa.scala 111:13]
    phv_data_185 <= io_pipe_phv_in_data_185; // @[matcher_pisa.scala 111:13]
    phv_data_186 <= io_pipe_phv_in_data_186; // @[matcher_pisa.scala 111:13]
    phv_data_187 <= io_pipe_phv_in_data_187; // @[matcher_pisa.scala 111:13]
    phv_data_188 <= io_pipe_phv_in_data_188; // @[matcher_pisa.scala 111:13]
    phv_data_189 <= io_pipe_phv_in_data_189; // @[matcher_pisa.scala 111:13]
    phv_data_190 <= io_pipe_phv_in_data_190; // @[matcher_pisa.scala 111:13]
    phv_data_191 <= io_pipe_phv_in_data_191; // @[matcher_pisa.scala 111:13]
    phv_data_192 <= io_pipe_phv_in_data_192; // @[matcher_pisa.scala 111:13]
    phv_data_193 <= io_pipe_phv_in_data_193; // @[matcher_pisa.scala 111:13]
    phv_data_194 <= io_pipe_phv_in_data_194; // @[matcher_pisa.scala 111:13]
    phv_data_195 <= io_pipe_phv_in_data_195; // @[matcher_pisa.scala 111:13]
    phv_data_196 <= io_pipe_phv_in_data_196; // @[matcher_pisa.scala 111:13]
    phv_data_197 <= io_pipe_phv_in_data_197; // @[matcher_pisa.scala 111:13]
    phv_data_198 <= io_pipe_phv_in_data_198; // @[matcher_pisa.scala 111:13]
    phv_data_199 <= io_pipe_phv_in_data_199; // @[matcher_pisa.scala 111:13]
    phv_data_200 <= io_pipe_phv_in_data_200; // @[matcher_pisa.scala 111:13]
    phv_data_201 <= io_pipe_phv_in_data_201; // @[matcher_pisa.scala 111:13]
    phv_data_202 <= io_pipe_phv_in_data_202; // @[matcher_pisa.scala 111:13]
    phv_data_203 <= io_pipe_phv_in_data_203; // @[matcher_pisa.scala 111:13]
    phv_data_204 <= io_pipe_phv_in_data_204; // @[matcher_pisa.scala 111:13]
    phv_data_205 <= io_pipe_phv_in_data_205; // @[matcher_pisa.scala 111:13]
    phv_data_206 <= io_pipe_phv_in_data_206; // @[matcher_pisa.scala 111:13]
    phv_data_207 <= io_pipe_phv_in_data_207; // @[matcher_pisa.scala 111:13]
    phv_data_208 <= io_pipe_phv_in_data_208; // @[matcher_pisa.scala 111:13]
    phv_data_209 <= io_pipe_phv_in_data_209; // @[matcher_pisa.scala 111:13]
    phv_data_210 <= io_pipe_phv_in_data_210; // @[matcher_pisa.scala 111:13]
    phv_data_211 <= io_pipe_phv_in_data_211; // @[matcher_pisa.scala 111:13]
    phv_data_212 <= io_pipe_phv_in_data_212; // @[matcher_pisa.scala 111:13]
    phv_data_213 <= io_pipe_phv_in_data_213; // @[matcher_pisa.scala 111:13]
    phv_data_214 <= io_pipe_phv_in_data_214; // @[matcher_pisa.scala 111:13]
    phv_data_215 <= io_pipe_phv_in_data_215; // @[matcher_pisa.scala 111:13]
    phv_data_216 <= io_pipe_phv_in_data_216; // @[matcher_pisa.scala 111:13]
    phv_data_217 <= io_pipe_phv_in_data_217; // @[matcher_pisa.scala 111:13]
    phv_data_218 <= io_pipe_phv_in_data_218; // @[matcher_pisa.scala 111:13]
    phv_data_219 <= io_pipe_phv_in_data_219; // @[matcher_pisa.scala 111:13]
    phv_data_220 <= io_pipe_phv_in_data_220; // @[matcher_pisa.scala 111:13]
    phv_data_221 <= io_pipe_phv_in_data_221; // @[matcher_pisa.scala 111:13]
    phv_data_222 <= io_pipe_phv_in_data_222; // @[matcher_pisa.scala 111:13]
    phv_data_223 <= io_pipe_phv_in_data_223; // @[matcher_pisa.scala 111:13]
    phv_data_224 <= io_pipe_phv_in_data_224; // @[matcher_pisa.scala 111:13]
    phv_data_225 <= io_pipe_phv_in_data_225; // @[matcher_pisa.scala 111:13]
    phv_data_226 <= io_pipe_phv_in_data_226; // @[matcher_pisa.scala 111:13]
    phv_data_227 <= io_pipe_phv_in_data_227; // @[matcher_pisa.scala 111:13]
    phv_data_228 <= io_pipe_phv_in_data_228; // @[matcher_pisa.scala 111:13]
    phv_data_229 <= io_pipe_phv_in_data_229; // @[matcher_pisa.scala 111:13]
    phv_data_230 <= io_pipe_phv_in_data_230; // @[matcher_pisa.scala 111:13]
    phv_data_231 <= io_pipe_phv_in_data_231; // @[matcher_pisa.scala 111:13]
    phv_data_232 <= io_pipe_phv_in_data_232; // @[matcher_pisa.scala 111:13]
    phv_data_233 <= io_pipe_phv_in_data_233; // @[matcher_pisa.scala 111:13]
    phv_data_234 <= io_pipe_phv_in_data_234; // @[matcher_pisa.scala 111:13]
    phv_data_235 <= io_pipe_phv_in_data_235; // @[matcher_pisa.scala 111:13]
    phv_data_236 <= io_pipe_phv_in_data_236; // @[matcher_pisa.scala 111:13]
    phv_data_237 <= io_pipe_phv_in_data_237; // @[matcher_pisa.scala 111:13]
    phv_data_238 <= io_pipe_phv_in_data_238; // @[matcher_pisa.scala 111:13]
    phv_data_239 <= io_pipe_phv_in_data_239; // @[matcher_pisa.scala 111:13]
    phv_data_240 <= io_pipe_phv_in_data_240; // @[matcher_pisa.scala 111:13]
    phv_data_241 <= io_pipe_phv_in_data_241; // @[matcher_pisa.scala 111:13]
    phv_data_242 <= io_pipe_phv_in_data_242; // @[matcher_pisa.scala 111:13]
    phv_data_243 <= io_pipe_phv_in_data_243; // @[matcher_pisa.scala 111:13]
    phv_data_244 <= io_pipe_phv_in_data_244; // @[matcher_pisa.scala 111:13]
    phv_data_245 <= io_pipe_phv_in_data_245; // @[matcher_pisa.scala 111:13]
    phv_data_246 <= io_pipe_phv_in_data_246; // @[matcher_pisa.scala 111:13]
    phv_data_247 <= io_pipe_phv_in_data_247; // @[matcher_pisa.scala 111:13]
    phv_data_248 <= io_pipe_phv_in_data_248; // @[matcher_pisa.scala 111:13]
    phv_data_249 <= io_pipe_phv_in_data_249; // @[matcher_pisa.scala 111:13]
    phv_data_250 <= io_pipe_phv_in_data_250; // @[matcher_pisa.scala 111:13]
    phv_data_251 <= io_pipe_phv_in_data_251; // @[matcher_pisa.scala 111:13]
    phv_data_252 <= io_pipe_phv_in_data_252; // @[matcher_pisa.scala 111:13]
    phv_data_253 <= io_pipe_phv_in_data_253; // @[matcher_pisa.scala 111:13]
    phv_data_254 <= io_pipe_phv_in_data_254; // @[matcher_pisa.scala 111:13]
    phv_data_255 <= io_pipe_phv_in_data_255; // @[matcher_pisa.scala 111:13]
    phv_data_256 <= io_pipe_phv_in_data_256; // @[matcher_pisa.scala 111:13]
    phv_data_257 <= io_pipe_phv_in_data_257; // @[matcher_pisa.scala 111:13]
    phv_data_258 <= io_pipe_phv_in_data_258; // @[matcher_pisa.scala 111:13]
    phv_data_259 <= io_pipe_phv_in_data_259; // @[matcher_pisa.scala 111:13]
    phv_data_260 <= io_pipe_phv_in_data_260; // @[matcher_pisa.scala 111:13]
    phv_data_261 <= io_pipe_phv_in_data_261; // @[matcher_pisa.scala 111:13]
    phv_data_262 <= io_pipe_phv_in_data_262; // @[matcher_pisa.scala 111:13]
    phv_data_263 <= io_pipe_phv_in_data_263; // @[matcher_pisa.scala 111:13]
    phv_data_264 <= io_pipe_phv_in_data_264; // @[matcher_pisa.scala 111:13]
    phv_data_265 <= io_pipe_phv_in_data_265; // @[matcher_pisa.scala 111:13]
    phv_data_266 <= io_pipe_phv_in_data_266; // @[matcher_pisa.scala 111:13]
    phv_data_267 <= io_pipe_phv_in_data_267; // @[matcher_pisa.scala 111:13]
    phv_data_268 <= io_pipe_phv_in_data_268; // @[matcher_pisa.scala 111:13]
    phv_data_269 <= io_pipe_phv_in_data_269; // @[matcher_pisa.scala 111:13]
    phv_data_270 <= io_pipe_phv_in_data_270; // @[matcher_pisa.scala 111:13]
    phv_data_271 <= io_pipe_phv_in_data_271; // @[matcher_pisa.scala 111:13]
    phv_data_272 <= io_pipe_phv_in_data_272; // @[matcher_pisa.scala 111:13]
    phv_data_273 <= io_pipe_phv_in_data_273; // @[matcher_pisa.scala 111:13]
    phv_data_274 <= io_pipe_phv_in_data_274; // @[matcher_pisa.scala 111:13]
    phv_data_275 <= io_pipe_phv_in_data_275; // @[matcher_pisa.scala 111:13]
    phv_data_276 <= io_pipe_phv_in_data_276; // @[matcher_pisa.scala 111:13]
    phv_data_277 <= io_pipe_phv_in_data_277; // @[matcher_pisa.scala 111:13]
    phv_data_278 <= io_pipe_phv_in_data_278; // @[matcher_pisa.scala 111:13]
    phv_data_279 <= io_pipe_phv_in_data_279; // @[matcher_pisa.scala 111:13]
    phv_data_280 <= io_pipe_phv_in_data_280; // @[matcher_pisa.scala 111:13]
    phv_data_281 <= io_pipe_phv_in_data_281; // @[matcher_pisa.scala 111:13]
    phv_data_282 <= io_pipe_phv_in_data_282; // @[matcher_pisa.scala 111:13]
    phv_data_283 <= io_pipe_phv_in_data_283; // @[matcher_pisa.scala 111:13]
    phv_data_284 <= io_pipe_phv_in_data_284; // @[matcher_pisa.scala 111:13]
    phv_data_285 <= io_pipe_phv_in_data_285; // @[matcher_pisa.scala 111:13]
    phv_data_286 <= io_pipe_phv_in_data_286; // @[matcher_pisa.scala 111:13]
    phv_data_287 <= io_pipe_phv_in_data_287; // @[matcher_pisa.scala 111:13]
    phv_data_288 <= io_pipe_phv_in_data_288; // @[matcher_pisa.scala 111:13]
    phv_data_289 <= io_pipe_phv_in_data_289; // @[matcher_pisa.scala 111:13]
    phv_data_290 <= io_pipe_phv_in_data_290; // @[matcher_pisa.scala 111:13]
    phv_data_291 <= io_pipe_phv_in_data_291; // @[matcher_pisa.scala 111:13]
    phv_data_292 <= io_pipe_phv_in_data_292; // @[matcher_pisa.scala 111:13]
    phv_data_293 <= io_pipe_phv_in_data_293; // @[matcher_pisa.scala 111:13]
    phv_data_294 <= io_pipe_phv_in_data_294; // @[matcher_pisa.scala 111:13]
    phv_data_295 <= io_pipe_phv_in_data_295; // @[matcher_pisa.scala 111:13]
    phv_data_296 <= io_pipe_phv_in_data_296; // @[matcher_pisa.scala 111:13]
    phv_data_297 <= io_pipe_phv_in_data_297; // @[matcher_pisa.scala 111:13]
    phv_data_298 <= io_pipe_phv_in_data_298; // @[matcher_pisa.scala 111:13]
    phv_data_299 <= io_pipe_phv_in_data_299; // @[matcher_pisa.scala 111:13]
    phv_data_300 <= io_pipe_phv_in_data_300; // @[matcher_pisa.scala 111:13]
    phv_data_301 <= io_pipe_phv_in_data_301; // @[matcher_pisa.scala 111:13]
    phv_data_302 <= io_pipe_phv_in_data_302; // @[matcher_pisa.scala 111:13]
    phv_data_303 <= io_pipe_phv_in_data_303; // @[matcher_pisa.scala 111:13]
    phv_data_304 <= io_pipe_phv_in_data_304; // @[matcher_pisa.scala 111:13]
    phv_data_305 <= io_pipe_phv_in_data_305; // @[matcher_pisa.scala 111:13]
    phv_data_306 <= io_pipe_phv_in_data_306; // @[matcher_pisa.scala 111:13]
    phv_data_307 <= io_pipe_phv_in_data_307; // @[matcher_pisa.scala 111:13]
    phv_data_308 <= io_pipe_phv_in_data_308; // @[matcher_pisa.scala 111:13]
    phv_data_309 <= io_pipe_phv_in_data_309; // @[matcher_pisa.scala 111:13]
    phv_data_310 <= io_pipe_phv_in_data_310; // @[matcher_pisa.scala 111:13]
    phv_data_311 <= io_pipe_phv_in_data_311; // @[matcher_pisa.scala 111:13]
    phv_data_312 <= io_pipe_phv_in_data_312; // @[matcher_pisa.scala 111:13]
    phv_data_313 <= io_pipe_phv_in_data_313; // @[matcher_pisa.scala 111:13]
    phv_data_314 <= io_pipe_phv_in_data_314; // @[matcher_pisa.scala 111:13]
    phv_data_315 <= io_pipe_phv_in_data_315; // @[matcher_pisa.scala 111:13]
    phv_data_316 <= io_pipe_phv_in_data_316; // @[matcher_pisa.scala 111:13]
    phv_data_317 <= io_pipe_phv_in_data_317; // @[matcher_pisa.scala 111:13]
    phv_data_318 <= io_pipe_phv_in_data_318; // @[matcher_pisa.scala 111:13]
    phv_data_319 <= io_pipe_phv_in_data_319; // @[matcher_pisa.scala 111:13]
    phv_data_320 <= io_pipe_phv_in_data_320; // @[matcher_pisa.scala 111:13]
    phv_data_321 <= io_pipe_phv_in_data_321; // @[matcher_pisa.scala 111:13]
    phv_data_322 <= io_pipe_phv_in_data_322; // @[matcher_pisa.scala 111:13]
    phv_data_323 <= io_pipe_phv_in_data_323; // @[matcher_pisa.scala 111:13]
    phv_data_324 <= io_pipe_phv_in_data_324; // @[matcher_pisa.scala 111:13]
    phv_data_325 <= io_pipe_phv_in_data_325; // @[matcher_pisa.scala 111:13]
    phv_data_326 <= io_pipe_phv_in_data_326; // @[matcher_pisa.scala 111:13]
    phv_data_327 <= io_pipe_phv_in_data_327; // @[matcher_pisa.scala 111:13]
    phv_data_328 <= io_pipe_phv_in_data_328; // @[matcher_pisa.scala 111:13]
    phv_data_329 <= io_pipe_phv_in_data_329; // @[matcher_pisa.scala 111:13]
    phv_data_330 <= io_pipe_phv_in_data_330; // @[matcher_pisa.scala 111:13]
    phv_data_331 <= io_pipe_phv_in_data_331; // @[matcher_pisa.scala 111:13]
    phv_data_332 <= io_pipe_phv_in_data_332; // @[matcher_pisa.scala 111:13]
    phv_data_333 <= io_pipe_phv_in_data_333; // @[matcher_pisa.scala 111:13]
    phv_data_334 <= io_pipe_phv_in_data_334; // @[matcher_pisa.scala 111:13]
    phv_data_335 <= io_pipe_phv_in_data_335; // @[matcher_pisa.scala 111:13]
    phv_data_336 <= io_pipe_phv_in_data_336; // @[matcher_pisa.scala 111:13]
    phv_data_337 <= io_pipe_phv_in_data_337; // @[matcher_pisa.scala 111:13]
    phv_data_338 <= io_pipe_phv_in_data_338; // @[matcher_pisa.scala 111:13]
    phv_data_339 <= io_pipe_phv_in_data_339; // @[matcher_pisa.scala 111:13]
    phv_data_340 <= io_pipe_phv_in_data_340; // @[matcher_pisa.scala 111:13]
    phv_data_341 <= io_pipe_phv_in_data_341; // @[matcher_pisa.scala 111:13]
    phv_data_342 <= io_pipe_phv_in_data_342; // @[matcher_pisa.scala 111:13]
    phv_data_343 <= io_pipe_phv_in_data_343; // @[matcher_pisa.scala 111:13]
    phv_data_344 <= io_pipe_phv_in_data_344; // @[matcher_pisa.scala 111:13]
    phv_data_345 <= io_pipe_phv_in_data_345; // @[matcher_pisa.scala 111:13]
    phv_data_346 <= io_pipe_phv_in_data_346; // @[matcher_pisa.scala 111:13]
    phv_data_347 <= io_pipe_phv_in_data_347; // @[matcher_pisa.scala 111:13]
    phv_data_348 <= io_pipe_phv_in_data_348; // @[matcher_pisa.scala 111:13]
    phv_data_349 <= io_pipe_phv_in_data_349; // @[matcher_pisa.scala 111:13]
    phv_data_350 <= io_pipe_phv_in_data_350; // @[matcher_pisa.scala 111:13]
    phv_data_351 <= io_pipe_phv_in_data_351; // @[matcher_pisa.scala 111:13]
    phv_data_352 <= io_pipe_phv_in_data_352; // @[matcher_pisa.scala 111:13]
    phv_data_353 <= io_pipe_phv_in_data_353; // @[matcher_pisa.scala 111:13]
    phv_data_354 <= io_pipe_phv_in_data_354; // @[matcher_pisa.scala 111:13]
    phv_data_355 <= io_pipe_phv_in_data_355; // @[matcher_pisa.scala 111:13]
    phv_data_356 <= io_pipe_phv_in_data_356; // @[matcher_pisa.scala 111:13]
    phv_data_357 <= io_pipe_phv_in_data_357; // @[matcher_pisa.scala 111:13]
    phv_data_358 <= io_pipe_phv_in_data_358; // @[matcher_pisa.scala 111:13]
    phv_data_359 <= io_pipe_phv_in_data_359; // @[matcher_pisa.scala 111:13]
    phv_data_360 <= io_pipe_phv_in_data_360; // @[matcher_pisa.scala 111:13]
    phv_data_361 <= io_pipe_phv_in_data_361; // @[matcher_pisa.scala 111:13]
    phv_data_362 <= io_pipe_phv_in_data_362; // @[matcher_pisa.scala 111:13]
    phv_data_363 <= io_pipe_phv_in_data_363; // @[matcher_pisa.scala 111:13]
    phv_data_364 <= io_pipe_phv_in_data_364; // @[matcher_pisa.scala 111:13]
    phv_data_365 <= io_pipe_phv_in_data_365; // @[matcher_pisa.scala 111:13]
    phv_data_366 <= io_pipe_phv_in_data_366; // @[matcher_pisa.scala 111:13]
    phv_data_367 <= io_pipe_phv_in_data_367; // @[matcher_pisa.scala 111:13]
    phv_data_368 <= io_pipe_phv_in_data_368; // @[matcher_pisa.scala 111:13]
    phv_data_369 <= io_pipe_phv_in_data_369; // @[matcher_pisa.scala 111:13]
    phv_data_370 <= io_pipe_phv_in_data_370; // @[matcher_pisa.scala 111:13]
    phv_data_371 <= io_pipe_phv_in_data_371; // @[matcher_pisa.scala 111:13]
    phv_data_372 <= io_pipe_phv_in_data_372; // @[matcher_pisa.scala 111:13]
    phv_data_373 <= io_pipe_phv_in_data_373; // @[matcher_pisa.scala 111:13]
    phv_data_374 <= io_pipe_phv_in_data_374; // @[matcher_pisa.scala 111:13]
    phv_data_375 <= io_pipe_phv_in_data_375; // @[matcher_pisa.scala 111:13]
    phv_data_376 <= io_pipe_phv_in_data_376; // @[matcher_pisa.scala 111:13]
    phv_data_377 <= io_pipe_phv_in_data_377; // @[matcher_pisa.scala 111:13]
    phv_data_378 <= io_pipe_phv_in_data_378; // @[matcher_pisa.scala 111:13]
    phv_data_379 <= io_pipe_phv_in_data_379; // @[matcher_pisa.scala 111:13]
    phv_data_380 <= io_pipe_phv_in_data_380; // @[matcher_pisa.scala 111:13]
    phv_data_381 <= io_pipe_phv_in_data_381; // @[matcher_pisa.scala 111:13]
    phv_data_382 <= io_pipe_phv_in_data_382; // @[matcher_pisa.scala 111:13]
    phv_data_383 <= io_pipe_phv_in_data_383; // @[matcher_pisa.scala 111:13]
    phv_data_384 <= io_pipe_phv_in_data_384; // @[matcher_pisa.scala 111:13]
    phv_data_385 <= io_pipe_phv_in_data_385; // @[matcher_pisa.scala 111:13]
    phv_data_386 <= io_pipe_phv_in_data_386; // @[matcher_pisa.scala 111:13]
    phv_data_387 <= io_pipe_phv_in_data_387; // @[matcher_pisa.scala 111:13]
    phv_data_388 <= io_pipe_phv_in_data_388; // @[matcher_pisa.scala 111:13]
    phv_data_389 <= io_pipe_phv_in_data_389; // @[matcher_pisa.scala 111:13]
    phv_data_390 <= io_pipe_phv_in_data_390; // @[matcher_pisa.scala 111:13]
    phv_data_391 <= io_pipe_phv_in_data_391; // @[matcher_pisa.scala 111:13]
    phv_data_392 <= io_pipe_phv_in_data_392; // @[matcher_pisa.scala 111:13]
    phv_data_393 <= io_pipe_phv_in_data_393; // @[matcher_pisa.scala 111:13]
    phv_data_394 <= io_pipe_phv_in_data_394; // @[matcher_pisa.scala 111:13]
    phv_data_395 <= io_pipe_phv_in_data_395; // @[matcher_pisa.scala 111:13]
    phv_data_396 <= io_pipe_phv_in_data_396; // @[matcher_pisa.scala 111:13]
    phv_data_397 <= io_pipe_phv_in_data_397; // @[matcher_pisa.scala 111:13]
    phv_data_398 <= io_pipe_phv_in_data_398; // @[matcher_pisa.scala 111:13]
    phv_data_399 <= io_pipe_phv_in_data_399; // @[matcher_pisa.scala 111:13]
    phv_data_400 <= io_pipe_phv_in_data_400; // @[matcher_pisa.scala 111:13]
    phv_data_401 <= io_pipe_phv_in_data_401; // @[matcher_pisa.scala 111:13]
    phv_data_402 <= io_pipe_phv_in_data_402; // @[matcher_pisa.scala 111:13]
    phv_data_403 <= io_pipe_phv_in_data_403; // @[matcher_pisa.scala 111:13]
    phv_data_404 <= io_pipe_phv_in_data_404; // @[matcher_pisa.scala 111:13]
    phv_data_405 <= io_pipe_phv_in_data_405; // @[matcher_pisa.scala 111:13]
    phv_data_406 <= io_pipe_phv_in_data_406; // @[matcher_pisa.scala 111:13]
    phv_data_407 <= io_pipe_phv_in_data_407; // @[matcher_pisa.scala 111:13]
    phv_data_408 <= io_pipe_phv_in_data_408; // @[matcher_pisa.scala 111:13]
    phv_data_409 <= io_pipe_phv_in_data_409; // @[matcher_pisa.scala 111:13]
    phv_data_410 <= io_pipe_phv_in_data_410; // @[matcher_pisa.scala 111:13]
    phv_data_411 <= io_pipe_phv_in_data_411; // @[matcher_pisa.scala 111:13]
    phv_data_412 <= io_pipe_phv_in_data_412; // @[matcher_pisa.scala 111:13]
    phv_data_413 <= io_pipe_phv_in_data_413; // @[matcher_pisa.scala 111:13]
    phv_data_414 <= io_pipe_phv_in_data_414; // @[matcher_pisa.scala 111:13]
    phv_data_415 <= io_pipe_phv_in_data_415; // @[matcher_pisa.scala 111:13]
    phv_data_416 <= io_pipe_phv_in_data_416; // @[matcher_pisa.scala 111:13]
    phv_data_417 <= io_pipe_phv_in_data_417; // @[matcher_pisa.scala 111:13]
    phv_data_418 <= io_pipe_phv_in_data_418; // @[matcher_pisa.scala 111:13]
    phv_data_419 <= io_pipe_phv_in_data_419; // @[matcher_pisa.scala 111:13]
    phv_data_420 <= io_pipe_phv_in_data_420; // @[matcher_pisa.scala 111:13]
    phv_data_421 <= io_pipe_phv_in_data_421; // @[matcher_pisa.scala 111:13]
    phv_data_422 <= io_pipe_phv_in_data_422; // @[matcher_pisa.scala 111:13]
    phv_data_423 <= io_pipe_phv_in_data_423; // @[matcher_pisa.scala 111:13]
    phv_data_424 <= io_pipe_phv_in_data_424; // @[matcher_pisa.scala 111:13]
    phv_data_425 <= io_pipe_phv_in_data_425; // @[matcher_pisa.scala 111:13]
    phv_data_426 <= io_pipe_phv_in_data_426; // @[matcher_pisa.scala 111:13]
    phv_data_427 <= io_pipe_phv_in_data_427; // @[matcher_pisa.scala 111:13]
    phv_data_428 <= io_pipe_phv_in_data_428; // @[matcher_pisa.scala 111:13]
    phv_data_429 <= io_pipe_phv_in_data_429; // @[matcher_pisa.scala 111:13]
    phv_data_430 <= io_pipe_phv_in_data_430; // @[matcher_pisa.scala 111:13]
    phv_data_431 <= io_pipe_phv_in_data_431; // @[matcher_pisa.scala 111:13]
    phv_data_432 <= io_pipe_phv_in_data_432; // @[matcher_pisa.scala 111:13]
    phv_data_433 <= io_pipe_phv_in_data_433; // @[matcher_pisa.scala 111:13]
    phv_data_434 <= io_pipe_phv_in_data_434; // @[matcher_pisa.scala 111:13]
    phv_data_435 <= io_pipe_phv_in_data_435; // @[matcher_pisa.scala 111:13]
    phv_data_436 <= io_pipe_phv_in_data_436; // @[matcher_pisa.scala 111:13]
    phv_data_437 <= io_pipe_phv_in_data_437; // @[matcher_pisa.scala 111:13]
    phv_data_438 <= io_pipe_phv_in_data_438; // @[matcher_pisa.scala 111:13]
    phv_data_439 <= io_pipe_phv_in_data_439; // @[matcher_pisa.scala 111:13]
    phv_data_440 <= io_pipe_phv_in_data_440; // @[matcher_pisa.scala 111:13]
    phv_data_441 <= io_pipe_phv_in_data_441; // @[matcher_pisa.scala 111:13]
    phv_data_442 <= io_pipe_phv_in_data_442; // @[matcher_pisa.scala 111:13]
    phv_data_443 <= io_pipe_phv_in_data_443; // @[matcher_pisa.scala 111:13]
    phv_data_444 <= io_pipe_phv_in_data_444; // @[matcher_pisa.scala 111:13]
    phv_data_445 <= io_pipe_phv_in_data_445; // @[matcher_pisa.scala 111:13]
    phv_data_446 <= io_pipe_phv_in_data_446; // @[matcher_pisa.scala 111:13]
    phv_data_447 <= io_pipe_phv_in_data_447; // @[matcher_pisa.scala 111:13]
    phv_data_448 <= io_pipe_phv_in_data_448; // @[matcher_pisa.scala 111:13]
    phv_data_449 <= io_pipe_phv_in_data_449; // @[matcher_pisa.scala 111:13]
    phv_data_450 <= io_pipe_phv_in_data_450; // @[matcher_pisa.scala 111:13]
    phv_data_451 <= io_pipe_phv_in_data_451; // @[matcher_pisa.scala 111:13]
    phv_data_452 <= io_pipe_phv_in_data_452; // @[matcher_pisa.scala 111:13]
    phv_data_453 <= io_pipe_phv_in_data_453; // @[matcher_pisa.scala 111:13]
    phv_data_454 <= io_pipe_phv_in_data_454; // @[matcher_pisa.scala 111:13]
    phv_data_455 <= io_pipe_phv_in_data_455; // @[matcher_pisa.scala 111:13]
    phv_data_456 <= io_pipe_phv_in_data_456; // @[matcher_pisa.scala 111:13]
    phv_data_457 <= io_pipe_phv_in_data_457; // @[matcher_pisa.scala 111:13]
    phv_data_458 <= io_pipe_phv_in_data_458; // @[matcher_pisa.scala 111:13]
    phv_data_459 <= io_pipe_phv_in_data_459; // @[matcher_pisa.scala 111:13]
    phv_data_460 <= io_pipe_phv_in_data_460; // @[matcher_pisa.scala 111:13]
    phv_data_461 <= io_pipe_phv_in_data_461; // @[matcher_pisa.scala 111:13]
    phv_data_462 <= io_pipe_phv_in_data_462; // @[matcher_pisa.scala 111:13]
    phv_data_463 <= io_pipe_phv_in_data_463; // @[matcher_pisa.scala 111:13]
    phv_data_464 <= io_pipe_phv_in_data_464; // @[matcher_pisa.scala 111:13]
    phv_data_465 <= io_pipe_phv_in_data_465; // @[matcher_pisa.scala 111:13]
    phv_data_466 <= io_pipe_phv_in_data_466; // @[matcher_pisa.scala 111:13]
    phv_data_467 <= io_pipe_phv_in_data_467; // @[matcher_pisa.scala 111:13]
    phv_data_468 <= io_pipe_phv_in_data_468; // @[matcher_pisa.scala 111:13]
    phv_data_469 <= io_pipe_phv_in_data_469; // @[matcher_pisa.scala 111:13]
    phv_data_470 <= io_pipe_phv_in_data_470; // @[matcher_pisa.scala 111:13]
    phv_data_471 <= io_pipe_phv_in_data_471; // @[matcher_pisa.scala 111:13]
    phv_data_472 <= io_pipe_phv_in_data_472; // @[matcher_pisa.scala 111:13]
    phv_data_473 <= io_pipe_phv_in_data_473; // @[matcher_pisa.scala 111:13]
    phv_data_474 <= io_pipe_phv_in_data_474; // @[matcher_pisa.scala 111:13]
    phv_data_475 <= io_pipe_phv_in_data_475; // @[matcher_pisa.scala 111:13]
    phv_data_476 <= io_pipe_phv_in_data_476; // @[matcher_pisa.scala 111:13]
    phv_data_477 <= io_pipe_phv_in_data_477; // @[matcher_pisa.scala 111:13]
    phv_data_478 <= io_pipe_phv_in_data_478; // @[matcher_pisa.scala 111:13]
    phv_data_479 <= io_pipe_phv_in_data_479; // @[matcher_pisa.scala 111:13]
    phv_data_480 <= io_pipe_phv_in_data_480; // @[matcher_pisa.scala 111:13]
    phv_data_481 <= io_pipe_phv_in_data_481; // @[matcher_pisa.scala 111:13]
    phv_data_482 <= io_pipe_phv_in_data_482; // @[matcher_pisa.scala 111:13]
    phv_data_483 <= io_pipe_phv_in_data_483; // @[matcher_pisa.scala 111:13]
    phv_data_484 <= io_pipe_phv_in_data_484; // @[matcher_pisa.scala 111:13]
    phv_data_485 <= io_pipe_phv_in_data_485; // @[matcher_pisa.scala 111:13]
    phv_data_486 <= io_pipe_phv_in_data_486; // @[matcher_pisa.scala 111:13]
    phv_data_487 <= io_pipe_phv_in_data_487; // @[matcher_pisa.scala 111:13]
    phv_data_488 <= io_pipe_phv_in_data_488; // @[matcher_pisa.scala 111:13]
    phv_data_489 <= io_pipe_phv_in_data_489; // @[matcher_pisa.scala 111:13]
    phv_data_490 <= io_pipe_phv_in_data_490; // @[matcher_pisa.scala 111:13]
    phv_data_491 <= io_pipe_phv_in_data_491; // @[matcher_pisa.scala 111:13]
    phv_data_492 <= io_pipe_phv_in_data_492; // @[matcher_pisa.scala 111:13]
    phv_data_493 <= io_pipe_phv_in_data_493; // @[matcher_pisa.scala 111:13]
    phv_data_494 <= io_pipe_phv_in_data_494; // @[matcher_pisa.scala 111:13]
    phv_data_495 <= io_pipe_phv_in_data_495; // @[matcher_pisa.scala 111:13]
    phv_data_496 <= io_pipe_phv_in_data_496; // @[matcher_pisa.scala 111:13]
    phv_data_497 <= io_pipe_phv_in_data_497; // @[matcher_pisa.scala 111:13]
    phv_data_498 <= io_pipe_phv_in_data_498; // @[matcher_pisa.scala 111:13]
    phv_data_499 <= io_pipe_phv_in_data_499; // @[matcher_pisa.scala 111:13]
    phv_data_500 <= io_pipe_phv_in_data_500; // @[matcher_pisa.scala 111:13]
    phv_data_501 <= io_pipe_phv_in_data_501; // @[matcher_pisa.scala 111:13]
    phv_data_502 <= io_pipe_phv_in_data_502; // @[matcher_pisa.scala 111:13]
    phv_data_503 <= io_pipe_phv_in_data_503; // @[matcher_pisa.scala 111:13]
    phv_data_504 <= io_pipe_phv_in_data_504; // @[matcher_pisa.scala 111:13]
    phv_data_505 <= io_pipe_phv_in_data_505; // @[matcher_pisa.scala 111:13]
    phv_data_506 <= io_pipe_phv_in_data_506; // @[matcher_pisa.scala 111:13]
    phv_data_507 <= io_pipe_phv_in_data_507; // @[matcher_pisa.scala 111:13]
    phv_data_508 <= io_pipe_phv_in_data_508; // @[matcher_pisa.scala 111:13]
    phv_data_509 <= io_pipe_phv_in_data_509; // @[matcher_pisa.scala 111:13]
    phv_data_510 <= io_pipe_phv_in_data_510; // @[matcher_pisa.scala 111:13]
    phv_data_511 <= io_pipe_phv_in_data_511; // @[matcher_pisa.scala 111:13]
    phv_next_processor_id <= io_pipe_phv_in_next_processor_id; // @[matcher_pisa.scala 111:13]
    phv_next_config_id <= io_pipe_phv_in_next_config_id; // @[matcher_pisa.scala 111:13]
    phv_is_valid_processor <= io_pipe_phv_in_is_valid_processor; // @[matcher_pisa.scala 111:13]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  phv_data_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  phv_data_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  phv_data_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  phv_data_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  phv_data_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  phv_data_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  phv_data_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  phv_data_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  phv_data_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  phv_data_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  phv_data_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  phv_data_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  phv_data_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  phv_data_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  phv_data_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  phv_data_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  phv_data_16 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  phv_data_17 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  phv_data_18 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  phv_data_19 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  phv_data_20 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  phv_data_21 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  phv_data_22 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  phv_data_23 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  phv_data_24 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  phv_data_25 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  phv_data_26 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  phv_data_27 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  phv_data_28 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  phv_data_29 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  phv_data_30 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  phv_data_31 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  phv_data_32 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  phv_data_33 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  phv_data_34 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  phv_data_35 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  phv_data_36 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  phv_data_37 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  phv_data_38 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  phv_data_39 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  phv_data_40 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  phv_data_41 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  phv_data_42 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  phv_data_43 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  phv_data_44 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  phv_data_45 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  phv_data_46 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  phv_data_47 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  phv_data_48 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  phv_data_49 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  phv_data_50 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  phv_data_51 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  phv_data_52 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  phv_data_53 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  phv_data_54 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  phv_data_55 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  phv_data_56 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  phv_data_57 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  phv_data_58 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  phv_data_59 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  phv_data_60 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  phv_data_61 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  phv_data_62 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  phv_data_63 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  phv_data_64 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  phv_data_65 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  phv_data_66 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  phv_data_67 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  phv_data_68 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  phv_data_69 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  phv_data_70 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  phv_data_71 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  phv_data_72 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  phv_data_73 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  phv_data_74 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  phv_data_75 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  phv_data_76 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  phv_data_77 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  phv_data_78 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  phv_data_79 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  phv_data_80 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  phv_data_81 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  phv_data_82 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  phv_data_83 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  phv_data_84 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  phv_data_85 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  phv_data_86 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  phv_data_87 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  phv_data_88 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  phv_data_89 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  phv_data_90 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  phv_data_91 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  phv_data_92 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  phv_data_93 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  phv_data_94 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  phv_data_95 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  phv_data_96 = _RAND_96[7:0];
  _RAND_97 = {1{`RANDOM}};
  phv_data_97 = _RAND_97[7:0];
  _RAND_98 = {1{`RANDOM}};
  phv_data_98 = _RAND_98[7:0];
  _RAND_99 = {1{`RANDOM}};
  phv_data_99 = _RAND_99[7:0];
  _RAND_100 = {1{`RANDOM}};
  phv_data_100 = _RAND_100[7:0];
  _RAND_101 = {1{`RANDOM}};
  phv_data_101 = _RAND_101[7:0];
  _RAND_102 = {1{`RANDOM}};
  phv_data_102 = _RAND_102[7:0];
  _RAND_103 = {1{`RANDOM}};
  phv_data_103 = _RAND_103[7:0];
  _RAND_104 = {1{`RANDOM}};
  phv_data_104 = _RAND_104[7:0];
  _RAND_105 = {1{`RANDOM}};
  phv_data_105 = _RAND_105[7:0];
  _RAND_106 = {1{`RANDOM}};
  phv_data_106 = _RAND_106[7:0];
  _RAND_107 = {1{`RANDOM}};
  phv_data_107 = _RAND_107[7:0];
  _RAND_108 = {1{`RANDOM}};
  phv_data_108 = _RAND_108[7:0];
  _RAND_109 = {1{`RANDOM}};
  phv_data_109 = _RAND_109[7:0];
  _RAND_110 = {1{`RANDOM}};
  phv_data_110 = _RAND_110[7:0];
  _RAND_111 = {1{`RANDOM}};
  phv_data_111 = _RAND_111[7:0];
  _RAND_112 = {1{`RANDOM}};
  phv_data_112 = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  phv_data_113 = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  phv_data_114 = _RAND_114[7:0];
  _RAND_115 = {1{`RANDOM}};
  phv_data_115 = _RAND_115[7:0];
  _RAND_116 = {1{`RANDOM}};
  phv_data_116 = _RAND_116[7:0];
  _RAND_117 = {1{`RANDOM}};
  phv_data_117 = _RAND_117[7:0];
  _RAND_118 = {1{`RANDOM}};
  phv_data_118 = _RAND_118[7:0];
  _RAND_119 = {1{`RANDOM}};
  phv_data_119 = _RAND_119[7:0];
  _RAND_120 = {1{`RANDOM}};
  phv_data_120 = _RAND_120[7:0];
  _RAND_121 = {1{`RANDOM}};
  phv_data_121 = _RAND_121[7:0];
  _RAND_122 = {1{`RANDOM}};
  phv_data_122 = _RAND_122[7:0];
  _RAND_123 = {1{`RANDOM}};
  phv_data_123 = _RAND_123[7:0];
  _RAND_124 = {1{`RANDOM}};
  phv_data_124 = _RAND_124[7:0];
  _RAND_125 = {1{`RANDOM}};
  phv_data_125 = _RAND_125[7:0];
  _RAND_126 = {1{`RANDOM}};
  phv_data_126 = _RAND_126[7:0];
  _RAND_127 = {1{`RANDOM}};
  phv_data_127 = _RAND_127[7:0];
  _RAND_128 = {1{`RANDOM}};
  phv_data_128 = _RAND_128[7:0];
  _RAND_129 = {1{`RANDOM}};
  phv_data_129 = _RAND_129[7:0];
  _RAND_130 = {1{`RANDOM}};
  phv_data_130 = _RAND_130[7:0];
  _RAND_131 = {1{`RANDOM}};
  phv_data_131 = _RAND_131[7:0];
  _RAND_132 = {1{`RANDOM}};
  phv_data_132 = _RAND_132[7:0];
  _RAND_133 = {1{`RANDOM}};
  phv_data_133 = _RAND_133[7:0];
  _RAND_134 = {1{`RANDOM}};
  phv_data_134 = _RAND_134[7:0];
  _RAND_135 = {1{`RANDOM}};
  phv_data_135 = _RAND_135[7:0];
  _RAND_136 = {1{`RANDOM}};
  phv_data_136 = _RAND_136[7:0];
  _RAND_137 = {1{`RANDOM}};
  phv_data_137 = _RAND_137[7:0];
  _RAND_138 = {1{`RANDOM}};
  phv_data_138 = _RAND_138[7:0];
  _RAND_139 = {1{`RANDOM}};
  phv_data_139 = _RAND_139[7:0];
  _RAND_140 = {1{`RANDOM}};
  phv_data_140 = _RAND_140[7:0];
  _RAND_141 = {1{`RANDOM}};
  phv_data_141 = _RAND_141[7:0];
  _RAND_142 = {1{`RANDOM}};
  phv_data_142 = _RAND_142[7:0];
  _RAND_143 = {1{`RANDOM}};
  phv_data_143 = _RAND_143[7:0];
  _RAND_144 = {1{`RANDOM}};
  phv_data_144 = _RAND_144[7:0];
  _RAND_145 = {1{`RANDOM}};
  phv_data_145 = _RAND_145[7:0];
  _RAND_146 = {1{`RANDOM}};
  phv_data_146 = _RAND_146[7:0];
  _RAND_147 = {1{`RANDOM}};
  phv_data_147 = _RAND_147[7:0];
  _RAND_148 = {1{`RANDOM}};
  phv_data_148 = _RAND_148[7:0];
  _RAND_149 = {1{`RANDOM}};
  phv_data_149 = _RAND_149[7:0];
  _RAND_150 = {1{`RANDOM}};
  phv_data_150 = _RAND_150[7:0];
  _RAND_151 = {1{`RANDOM}};
  phv_data_151 = _RAND_151[7:0];
  _RAND_152 = {1{`RANDOM}};
  phv_data_152 = _RAND_152[7:0];
  _RAND_153 = {1{`RANDOM}};
  phv_data_153 = _RAND_153[7:0];
  _RAND_154 = {1{`RANDOM}};
  phv_data_154 = _RAND_154[7:0];
  _RAND_155 = {1{`RANDOM}};
  phv_data_155 = _RAND_155[7:0];
  _RAND_156 = {1{`RANDOM}};
  phv_data_156 = _RAND_156[7:0];
  _RAND_157 = {1{`RANDOM}};
  phv_data_157 = _RAND_157[7:0];
  _RAND_158 = {1{`RANDOM}};
  phv_data_158 = _RAND_158[7:0];
  _RAND_159 = {1{`RANDOM}};
  phv_data_159 = _RAND_159[7:0];
  _RAND_160 = {1{`RANDOM}};
  phv_data_160 = _RAND_160[7:0];
  _RAND_161 = {1{`RANDOM}};
  phv_data_161 = _RAND_161[7:0];
  _RAND_162 = {1{`RANDOM}};
  phv_data_162 = _RAND_162[7:0];
  _RAND_163 = {1{`RANDOM}};
  phv_data_163 = _RAND_163[7:0];
  _RAND_164 = {1{`RANDOM}};
  phv_data_164 = _RAND_164[7:0];
  _RAND_165 = {1{`RANDOM}};
  phv_data_165 = _RAND_165[7:0];
  _RAND_166 = {1{`RANDOM}};
  phv_data_166 = _RAND_166[7:0];
  _RAND_167 = {1{`RANDOM}};
  phv_data_167 = _RAND_167[7:0];
  _RAND_168 = {1{`RANDOM}};
  phv_data_168 = _RAND_168[7:0];
  _RAND_169 = {1{`RANDOM}};
  phv_data_169 = _RAND_169[7:0];
  _RAND_170 = {1{`RANDOM}};
  phv_data_170 = _RAND_170[7:0];
  _RAND_171 = {1{`RANDOM}};
  phv_data_171 = _RAND_171[7:0];
  _RAND_172 = {1{`RANDOM}};
  phv_data_172 = _RAND_172[7:0];
  _RAND_173 = {1{`RANDOM}};
  phv_data_173 = _RAND_173[7:0];
  _RAND_174 = {1{`RANDOM}};
  phv_data_174 = _RAND_174[7:0];
  _RAND_175 = {1{`RANDOM}};
  phv_data_175 = _RAND_175[7:0];
  _RAND_176 = {1{`RANDOM}};
  phv_data_176 = _RAND_176[7:0];
  _RAND_177 = {1{`RANDOM}};
  phv_data_177 = _RAND_177[7:0];
  _RAND_178 = {1{`RANDOM}};
  phv_data_178 = _RAND_178[7:0];
  _RAND_179 = {1{`RANDOM}};
  phv_data_179 = _RAND_179[7:0];
  _RAND_180 = {1{`RANDOM}};
  phv_data_180 = _RAND_180[7:0];
  _RAND_181 = {1{`RANDOM}};
  phv_data_181 = _RAND_181[7:0];
  _RAND_182 = {1{`RANDOM}};
  phv_data_182 = _RAND_182[7:0];
  _RAND_183 = {1{`RANDOM}};
  phv_data_183 = _RAND_183[7:0];
  _RAND_184 = {1{`RANDOM}};
  phv_data_184 = _RAND_184[7:0];
  _RAND_185 = {1{`RANDOM}};
  phv_data_185 = _RAND_185[7:0];
  _RAND_186 = {1{`RANDOM}};
  phv_data_186 = _RAND_186[7:0];
  _RAND_187 = {1{`RANDOM}};
  phv_data_187 = _RAND_187[7:0];
  _RAND_188 = {1{`RANDOM}};
  phv_data_188 = _RAND_188[7:0];
  _RAND_189 = {1{`RANDOM}};
  phv_data_189 = _RAND_189[7:0];
  _RAND_190 = {1{`RANDOM}};
  phv_data_190 = _RAND_190[7:0];
  _RAND_191 = {1{`RANDOM}};
  phv_data_191 = _RAND_191[7:0];
  _RAND_192 = {1{`RANDOM}};
  phv_data_192 = _RAND_192[7:0];
  _RAND_193 = {1{`RANDOM}};
  phv_data_193 = _RAND_193[7:0];
  _RAND_194 = {1{`RANDOM}};
  phv_data_194 = _RAND_194[7:0];
  _RAND_195 = {1{`RANDOM}};
  phv_data_195 = _RAND_195[7:0];
  _RAND_196 = {1{`RANDOM}};
  phv_data_196 = _RAND_196[7:0];
  _RAND_197 = {1{`RANDOM}};
  phv_data_197 = _RAND_197[7:0];
  _RAND_198 = {1{`RANDOM}};
  phv_data_198 = _RAND_198[7:0];
  _RAND_199 = {1{`RANDOM}};
  phv_data_199 = _RAND_199[7:0];
  _RAND_200 = {1{`RANDOM}};
  phv_data_200 = _RAND_200[7:0];
  _RAND_201 = {1{`RANDOM}};
  phv_data_201 = _RAND_201[7:0];
  _RAND_202 = {1{`RANDOM}};
  phv_data_202 = _RAND_202[7:0];
  _RAND_203 = {1{`RANDOM}};
  phv_data_203 = _RAND_203[7:0];
  _RAND_204 = {1{`RANDOM}};
  phv_data_204 = _RAND_204[7:0];
  _RAND_205 = {1{`RANDOM}};
  phv_data_205 = _RAND_205[7:0];
  _RAND_206 = {1{`RANDOM}};
  phv_data_206 = _RAND_206[7:0];
  _RAND_207 = {1{`RANDOM}};
  phv_data_207 = _RAND_207[7:0];
  _RAND_208 = {1{`RANDOM}};
  phv_data_208 = _RAND_208[7:0];
  _RAND_209 = {1{`RANDOM}};
  phv_data_209 = _RAND_209[7:0];
  _RAND_210 = {1{`RANDOM}};
  phv_data_210 = _RAND_210[7:0];
  _RAND_211 = {1{`RANDOM}};
  phv_data_211 = _RAND_211[7:0];
  _RAND_212 = {1{`RANDOM}};
  phv_data_212 = _RAND_212[7:0];
  _RAND_213 = {1{`RANDOM}};
  phv_data_213 = _RAND_213[7:0];
  _RAND_214 = {1{`RANDOM}};
  phv_data_214 = _RAND_214[7:0];
  _RAND_215 = {1{`RANDOM}};
  phv_data_215 = _RAND_215[7:0];
  _RAND_216 = {1{`RANDOM}};
  phv_data_216 = _RAND_216[7:0];
  _RAND_217 = {1{`RANDOM}};
  phv_data_217 = _RAND_217[7:0];
  _RAND_218 = {1{`RANDOM}};
  phv_data_218 = _RAND_218[7:0];
  _RAND_219 = {1{`RANDOM}};
  phv_data_219 = _RAND_219[7:0];
  _RAND_220 = {1{`RANDOM}};
  phv_data_220 = _RAND_220[7:0];
  _RAND_221 = {1{`RANDOM}};
  phv_data_221 = _RAND_221[7:0];
  _RAND_222 = {1{`RANDOM}};
  phv_data_222 = _RAND_222[7:0];
  _RAND_223 = {1{`RANDOM}};
  phv_data_223 = _RAND_223[7:0];
  _RAND_224 = {1{`RANDOM}};
  phv_data_224 = _RAND_224[7:0];
  _RAND_225 = {1{`RANDOM}};
  phv_data_225 = _RAND_225[7:0];
  _RAND_226 = {1{`RANDOM}};
  phv_data_226 = _RAND_226[7:0];
  _RAND_227 = {1{`RANDOM}};
  phv_data_227 = _RAND_227[7:0];
  _RAND_228 = {1{`RANDOM}};
  phv_data_228 = _RAND_228[7:0];
  _RAND_229 = {1{`RANDOM}};
  phv_data_229 = _RAND_229[7:0];
  _RAND_230 = {1{`RANDOM}};
  phv_data_230 = _RAND_230[7:0];
  _RAND_231 = {1{`RANDOM}};
  phv_data_231 = _RAND_231[7:0];
  _RAND_232 = {1{`RANDOM}};
  phv_data_232 = _RAND_232[7:0];
  _RAND_233 = {1{`RANDOM}};
  phv_data_233 = _RAND_233[7:0];
  _RAND_234 = {1{`RANDOM}};
  phv_data_234 = _RAND_234[7:0];
  _RAND_235 = {1{`RANDOM}};
  phv_data_235 = _RAND_235[7:0];
  _RAND_236 = {1{`RANDOM}};
  phv_data_236 = _RAND_236[7:0];
  _RAND_237 = {1{`RANDOM}};
  phv_data_237 = _RAND_237[7:0];
  _RAND_238 = {1{`RANDOM}};
  phv_data_238 = _RAND_238[7:0];
  _RAND_239 = {1{`RANDOM}};
  phv_data_239 = _RAND_239[7:0];
  _RAND_240 = {1{`RANDOM}};
  phv_data_240 = _RAND_240[7:0];
  _RAND_241 = {1{`RANDOM}};
  phv_data_241 = _RAND_241[7:0];
  _RAND_242 = {1{`RANDOM}};
  phv_data_242 = _RAND_242[7:0];
  _RAND_243 = {1{`RANDOM}};
  phv_data_243 = _RAND_243[7:0];
  _RAND_244 = {1{`RANDOM}};
  phv_data_244 = _RAND_244[7:0];
  _RAND_245 = {1{`RANDOM}};
  phv_data_245 = _RAND_245[7:0];
  _RAND_246 = {1{`RANDOM}};
  phv_data_246 = _RAND_246[7:0];
  _RAND_247 = {1{`RANDOM}};
  phv_data_247 = _RAND_247[7:0];
  _RAND_248 = {1{`RANDOM}};
  phv_data_248 = _RAND_248[7:0];
  _RAND_249 = {1{`RANDOM}};
  phv_data_249 = _RAND_249[7:0];
  _RAND_250 = {1{`RANDOM}};
  phv_data_250 = _RAND_250[7:0];
  _RAND_251 = {1{`RANDOM}};
  phv_data_251 = _RAND_251[7:0];
  _RAND_252 = {1{`RANDOM}};
  phv_data_252 = _RAND_252[7:0];
  _RAND_253 = {1{`RANDOM}};
  phv_data_253 = _RAND_253[7:0];
  _RAND_254 = {1{`RANDOM}};
  phv_data_254 = _RAND_254[7:0];
  _RAND_255 = {1{`RANDOM}};
  phv_data_255 = _RAND_255[7:0];
  _RAND_256 = {1{`RANDOM}};
  phv_data_256 = _RAND_256[7:0];
  _RAND_257 = {1{`RANDOM}};
  phv_data_257 = _RAND_257[7:0];
  _RAND_258 = {1{`RANDOM}};
  phv_data_258 = _RAND_258[7:0];
  _RAND_259 = {1{`RANDOM}};
  phv_data_259 = _RAND_259[7:0];
  _RAND_260 = {1{`RANDOM}};
  phv_data_260 = _RAND_260[7:0];
  _RAND_261 = {1{`RANDOM}};
  phv_data_261 = _RAND_261[7:0];
  _RAND_262 = {1{`RANDOM}};
  phv_data_262 = _RAND_262[7:0];
  _RAND_263 = {1{`RANDOM}};
  phv_data_263 = _RAND_263[7:0];
  _RAND_264 = {1{`RANDOM}};
  phv_data_264 = _RAND_264[7:0];
  _RAND_265 = {1{`RANDOM}};
  phv_data_265 = _RAND_265[7:0];
  _RAND_266 = {1{`RANDOM}};
  phv_data_266 = _RAND_266[7:0];
  _RAND_267 = {1{`RANDOM}};
  phv_data_267 = _RAND_267[7:0];
  _RAND_268 = {1{`RANDOM}};
  phv_data_268 = _RAND_268[7:0];
  _RAND_269 = {1{`RANDOM}};
  phv_data_269 = _RAND_269[7:0];
  _RAND_270 = {1{`RANDOM}};
  phv_data_270 = _RAND_270[7:0];
  _RAND_271 = {1{`RANDOM}};
  phv_data_271 = _RAND_271[7:0];
  _RAND_272 = {1{`RANDOM}};
  phv_data_272 = _RAND_272[7:0];
  _RAND_273 = {1{`RANDOM}};
  phv_data_273 = _RAND_273[7:0];
  _RAND_274 = {1{`RANDOM}};
  phv_data_274 = _RAND_274[7:0];
  _RAND_275 = {1{`RANDOM}};
  phv_data_275 = _RAND_275[7:0];
  _RAND_276 = {1{`RANDOM}};
  phv_data_276 = _RAND_276[7:0];
  _RAND_277 = {1{`RANDOM}};
  phv_data_277 = _RAND_277[7:0];
  _RAND_278 = {1{`RANDOM}};
  phv_data_278 = _RAND_278[7:0];
  _RAND_279 = {1{`RANDOM}};
  phv_data_279 = _RAND_279[7:0];
  _RAND_280 = {1{`RANDOM}};
  phv_data_280 = _RAND_280[7:0];
  _RAND_281 = {1{`RANDOM}};
  phv_data_281 = _RAND_281[7:0];
  _RAND_282 = {1{`RANDOM}};
  phv_data_282 = _RAND_282[7:0];
  _RAND_283 = {1{`RANDOM}};
  phv_data_283 = _RAND_283[7:0];
  _RAND_284 = {1{`RANDOM}};
  phv_data_284 = _RAND_284[7:0];
  _RAND_285 = {1{`RANDOM}};
  phv_data_285 = _RAND_285[7:0];
  _RAND_286 = {1{`RANDOM}};
  phv_data_286 = _RAND_286[7:0];
  _RAND_287 = {1{`RANDOM}};
  phv_data_287 = _RAND_287[7:0];
  _RAND_288 = {1{`RANDOM}};
  phv_data_288 = _RAND_288[7:0];
  _RAND_289 = {1{`RANDOM}};
  phv_data_289 = _RAND_289[7:0];
  _RAND_290 = {1{`RANDOM}};
  phv_data_290 = _RAND_290[7:0];
  _RAND_291 = {1{`RANDOM}};
  phv_data_291 = _RAND_291[7:0];
  _RAND_292 = {1{`RANDOM}};
  phv_data_292 = _RAND_292[7:0];
  _RAND_293 = {1{`RANDOM}};
  phv_data_293 = _RAND_293[7:0];
  _RAND_294 = {1{`RANDOM}};
  phv_data_294 = _RAND_294[7:0];
  _RAND_295 = {1{`RANDOM}};
  phv_data_295 = _RAND_295[7:0];
  _RAND_296 = {1{`RANDOM}};
  phv_data_296 = _RAND_296[7:0];
  _RAND_297 = {1{`RANDOM}};
  phv_data_297 = _RAND_297[7:0];
  _RAND_298 = {1{`RANDOM}};
  phv_data_298 = _RAND_298[7:0];
  _RAND_299 = {1{`RANDOM}};
  phv_data_299 = _RAND_299[7:0];
  _RAND_300 = {1{`RANDOM}};
  phv_data_300 = _RAND_300[7:0];
  _RAND_301 = {1{`RANDOM}};
  phv_data_301 = _RAND_301[7:0];
  _RAND_302 = {1{`RANDOM}};
  phv_data_302 = _RAND_302[7:0];
  _RAND_303 = {1{`RANDOM}};
  phv_data_303 = _RAND_303[7:0];
  _RAND_304 = {1{`RANDOM}};
  phv_data_304 = _RAND_304[7:0];
  _RAND_305 = {1{`RANDOM}};
  phv_data_305 = _RAND_305[7:0];
  _RAND_306 = {1{`RANDOM}};
  phv_data_306 = _RAND_306[7:0];
  _RAND_307 = {1{`RANDOM}};
  phv_data_307 = _RAND_307[7:0];
  _RAND_308 = {1{`RANDOM}};
  phv_data_308 = _RAND_308[7:0];
  _RAND_309 = {1{`RANDOM}};
  phv_data_309 = _RAND_309[7:0];
  _RAND_310 = {1{`RANDOM}};
  phv_data_310 = _RAND_310[7:0];
  _RAND_311 = {1{`RANDOM}};
  phv_data_311 = _RAND_311[7:0];
  _RAND_312 = {1{`RANDOM}};
  phv_data_312 = _RAND_312[7:0];
  _RAND_313 = {1{`RANDOM}};
  phv_data_313 = _RAND_313[7:0];
  _RAND_314 = {1{`RANDOM}};
  phv_data_314 = _RAND_314[7:0];
  _RAND_315 = {1{`RANDOM}};
  phv_data_315 = _RAND_315[7:0];
  _RAND_316 = {1{`RANDOM}};
  phv_data_316 = _RAND_316[7:0];
  _RAND_317 = {1{`RANDOM}};
  phv_data_317 = _RAND_317[7:0];
  _RAND_318 = {1{`RANDOM}};
  phv_data_318 = _RAND_318[7:0];
  _RAND_319 = {1{`RANDOM}};
  phv_data_319 = _RAND_319[7:0];
  _RAND_320 = {1{`RANDOM}};
  phv_data_320 = _RAND_320[7:0];
  _RAND_321 = {1{`RANDOM}};
  phv_data_321 = _RAND_321[7:0];
  _RAND_322 = {1{`RANDOM}};
  phv_data_322 = _RAND_322[7:0];
  _RAND_323 = {1{`RANDOM}};
  phv_data_323 = _RAND_323[7:0];
  _RAND_324 = {1{`RANDOM}};
  phv_data_324 = _RAND_324[7:0];
  _RAND_325 = {1{`RANDOM}};
  phv_data_325 = _RAND_325[7:0];
  _RAND_326 = {1{`RANDOM}};
  phv_data_326 = _RAND_326[7:0];
  _RAND_327 = {1{`RANDOM}};
  phv_data_327 = _RAND_327[7:0];
  _RAND_328 = {1{`RANDOM}};
  phv_data_328 = _RAND_328[7:0];
  _RAND_329 = {1{`RANDOM}};
  phv_data_329 = _RAND_329[7:0];
  _RAND_330 = {1{`RANDOM}};
  phv_data_330 = _RAND_330[7:0];
  _RAND_331 = {1{`RANDOM}};
  phv_data_331 = _RAND_331[7:0];
  _RAND_332 = {1{`RANDOM}};
  phv_data_332 = _RAND_332[7:0];
  _RAND_333 = {1{`RANDOM}};
  phv_data_333 = _RAND_333[7:0];
  _RAND_334 = {1{`RANDOM}};
  phv_data_334 = _RAND_334[7:0];
  _RAND_335 = {1{`RANDOM}};
  phv_data_335 = _RAND_335[7:0];
  _RAND_336 = {1{`RANDOM}};
  phv_data_336 = _RAND_336[7:0];
  _RAND_337 = {1{`RANDOM}};
  phv_data_337 = _RAND_337[7:0];
  _RAND_338 = {1{`RANDOM}};
  phv_data_338 = _RAND_338[7:0];
  _RAND_339 = {1{`RANDOM}};
  phv_data_339 = _RAND_339[7:0];
  _RAND_340 = {1{`RANDOM}};
  phv_data_340 = _RAND_340[7:0];
  _RAND_341 = {1{`RANDOM}};
  phv_data_341 = _RAND_341[7:0];
  _RAND_342 = {1{`RANDOM}};
  phv_data_342 = _RAND_342[7:0];
  _RAND_343 = {1{`RANDOM}};
  phv_data_343 = _RAND_343[7:0];
  _RAND_344 = {1{`RANDOM}};
  phv_data_344 = _RAND_344[7:0];
  _RAND_345 = {1{`RANDOM}};
  phv_data_345 = _RAND_345[7:0];
  _RAND_346 = {1{`RANDOM}};
  phv_data_346 = _RAND_346[7:0];
  _RAND_347 = {1{`RANDOM}};
  phv_data_347 = _RAND_347[7:0];
  _RAND_348 = {1{`RANDOM}};
  phv_data_348 = _RAND_348[7:0];
  _RAND_349 = {1{`RANDOM}};
  phv_data_349 = _RAND_349[7:0];
  _RAND_350 = {1{`RANDOM}};
  phv_data_350 = _RAND_350[7:0];
  _RAND_351 = {1{`RANDOM}};
  phv_data_351 = _RAND_351[7:0];
  _RAND_352 = {1{`RANDOM}};
  phv_data_352 = _RAND_352[7:0];
  _RAND_353 = {1{`RANDOM}};
  phv_data_353 = _RAND_353[7:0];
  _RAND_354 = {1{`RANDOM}};
  phv_data_354 = _RAND_354[7:0];
  _RAND_355 = {1{`RANDOM}};
  phv_data_355 = _RAND_355[7:0];
  _RAND_356 = {1{`RANDOM}};
  phv_data_356 = _RAND_356[7:0];
  _RAND_357 = {1{`RANDOM}};
  phv_data_357 = _RAND_357[7:0];
  _RAND_358 = {1{`RANDOM}};
  phv_data_358 = _RAND_358[7:0];
  _RAND_359 = {1{`RANDOM}};
  phv_data_359 = _RAND_359[7:0];
  _RAND_360 = {1{`RANDOM}};
  phv_data_360 = _RAND_360[7:0];
  _RAND_361 = {1{`RANDOM}};
  phv_data_361 = _RAND_361[7:0];
  _RAND_362 = {1{`RANDOM}};
  phv_data_362 = _RAND_362[7:0];
  _RAND_363 = {1{`RANDOM}};
  phv_data_363 = _RAND_363[7:0];
  _RAND_364 = {1{`RANDOM}};
  phv_data_364 = _RAND_364[7:0];
  _RAND_365 = {1{`RANDOM}};
  phv_data_365 = _RAND_365[7:0];
  _RAND_366 = {1{`RANDOM}};
  phv_data_366 = _RAND_366[7:0];
  _RAND_367 = {1{`RANDOM}};
  phv_data_367 = _RAND_367[7:0];
  _RAND_368 = {1{`RANDOM}};
  phv_data_368 = _RAND_368[7:0];
  _RAND_369 = {1{`RANDOM}};
  phv_data_369 = _RAND_369[7:0];
  _RAND_370 = {1{`RANDOM}};
  phv_data_370 = _RAND_370[7:0];
  _RAND_371 = {1{`RANDOM}};
  phv_data_371 = _RAND_371[7:0];
  _RAND_372 = {1{`RANDOM}};
  phv_data_372 = _RAND_372[7:0];
  _RAND_373 = {1{`RANDOM}};
  phv_data_373 = _RAND_373[7:0];
  _RAND_374 = {1{`RANDOM}};
  phv_data_374 = _RAND_374[7:0];
  _RAND_375 = {1{`RANDOM}};
  phv_data_375 = _RAND_375[7:0];
  _RAND_376 = {1{`RANDOM}};
  phv_data_376 = _RAND_376[7:0];
  _RAND_377 = {1{`RANDOM}};
  phv_data_377 = _RAND_377[7:0];
  _RAND_378 = {1{`RANDOM}};
  phv_data_378 = _RAND_378[7:0];
  _RAND_379 = {1{`RANDOM}};
  phv_data_379 = _RAND_379[7:0];
  _RAND_380 = {1{`RANDOM}};
  phv_data_380 = _RAND_380[7:0];
  _RAND_381 = {1{`RANDOM}};
  phv_data_381 = _RAND_381[7:0];
  _RAND_382 = {1{`RANDOM}};
  phv_data_382 = _RAND_382[7:0];
  _RAND_383 = {1{`RANDOM}};
  phv_data_383 = _RAND_383[7:0];
  _RAND_384 = {1{`RANDOM}};
  phv_data_384 = _RAND_384[7:0];
  _RAND_385 = {1{`RANDOM}};
  phv_data_385 = _RAND_385[7:0];
  _RAND_386 = {1{`RANDOM}};
  phv_data_386 = _RAND_386[7:0];
  _RAND_387 = {1{`RANDOM}};
  phv_data_387 = _RAND_387[7:0];
  _RAND_388 = {1{`RANDOM}};
  phv_data_388 = _RAND_388[7:0];
  _RAND_389 = {1{`RANDOM}};
  phv_data_389 = _RAND_389[7:0];
  _RAND_390 = {1{`RANDOM}};
  phv_data_390 = _RAND_390[7:0];
  _RAND_391 = {1{`RANDOM}};
  phv_data_391 = _RAND_391[7:0];
  _RAND_392 = {1{`RANDOM}};
  phv_data_392 = _RAND_392[7:0];
  _RAND_393 = {1{`RANDOM}};
  phv_data_393 = _RAND_393[7:0];
  _RAND_394 = {1{`RANDOM}};
  phv_data_394 = _RAND_394[7:0];
  _RAND_395 = {1{`RANDOM}};
  phv_data_395 = _RAND_395[7:0];
  _RAND_396 = {1{`RANDOM}};
  phv_data_396 = _RAND_396[7:0];
  _RAND_397 = {1{`RANDOM}};
  phv_data_397 = _RAND_397[7:0];
  _RAND_398 = {1{`RANDOM}};
  phv_data_398 = _RAND_398[7:0];
  _RAND_399 = {1{`RANDOM}};
  phv_data_399 = _RAND_399[7:0];
  _RAND_400 = {1{`RANDOM}};
  phv_data_400 = _RAND_400[7:0];
  _RAND_401 = {1{`RANDOM}};
  phv_data_401 = _RAND_401[7:0];
  _RAND_402 = {1{`RANDOM}};
  phv_data_402 = _RAND_402[7:0];
  _RAND_403 = {1{`RANDOM}};
  phv_data_403 = _RAND_403[7:0];
  _RAND_404 = {1{`RANDOM}};
  phv_data_404 = _RAND_404[7:0];
  _RAND_405 = {1{`RANDOM}};
  phv_data_405 = _RAND_405[7:0];
  _RAND_406 = {1{`RANDOM}};
  phv_data_406 = _RAND_406[7:0];
  _RAND_407 = {1{`RANDOM}};
  phv_data_407 = _RAND_407[7:0];
  _RAND_408 = {1{`RANDOM}};
  phv_data_408 = _RAND_408[7:0];
  _RAND_409 = {1{`RANDOM}};
  phv_data_409 = _RAND_409[7:0];
  _RAND_410 = {1{`RANDOM}};
  phv_data_410 = _RAND_410[7:0];
  _RAND_411 = {1{`RANDOM}};
  phv_data_411 = _RAND_411[7:0];
  _RAND_412 = {1{`RANDOM}};
  phv_data_412 = _RAND_412[7:0];
  _RAND_413 = {1{`RANDOM}};
  phv_data_413 = _RAND_413[7:0];
  _RAND_414 = {1{`RANDOM}};
  phv_data_414 = _RAND_414[7:0];
  _RAND_415 = {1{`RANDOM}};
  phv_data_415 = _RAND_415[7:0];
  _RAND_416 = {1{`RANDOM}};
  phv_data_416 = _RAND_416[7:0];
  _RAND_417 = {1{`RANDOM}};
  phv_data_417 = _RAND_417[7:0];
  _RAND_418 = {1{`RANDOM}};
  phv_data_418 = _RAND_418[7:0];
  _RAND_419 = {1{`RANDOM}};
  phv_data_419 = _RAND_419[7:0];
  _RAND_420 = {1{`RANDOM}};
  phv_data_420 = _RAND_420[7:0];
  _RAND_421 = {1{`RANDOM}};
  phv_data_421 = _RAND_421[7:0];
  _RAND_422 = {1{`RANDOM}};
  phv_data_422 = _RAND_422[7:0];
  _RAND_423 = {1{`RANDOM}};
  phv_data_423 = _RAND_423[7:0];
  _RAND_424 = {1{`RANDOM}};
  phv_data_424 = _RAND_424[7:0];
  _RAND_425 = {1{`RANDOM}};
  phv_data_425 = _RAND_425[7:0];
  _RAND_426 = {1{`RANDOM}};
  phv_data_426 = _RAND_426[7:0];
  _RAND_427 = {1{`RANDOM}};
  phv_data_427 = _RAND_427[7:0];
  _RAND_428 = {1{`RANDOM}};
  phv_data_428 = _RAND_428[7:0];
  _RAND_429 = {1{`RANDOM}};
  phv_data_429 = _RAND_429[7:0];
  _RAND_430 = {1{`RANDOM}};
  phv_data_430 = _RAND_430[7:0];
  _RAND_431 = {1{`RANDOM}};
  phv_data_431 = _RAND_431[7:0];
  _RAND_432 = {1{`RANDOM}};
  phv_data_432 = _RAND_432[7:0];
  _RAND_433 = {1{`RANDOM}};
  phv_data_433 = _RAND_433[7:0];
  _RAND_434 = {1{`RANDOM}};
  phv_data_434 = _RAND_434[7:0];
  _RAND_435 = {1{`RANDOM}};
  phv_data_435 = _RAND_435[7:0];
  _RAND_436 = {1{`RANDOM}};
  phv_data_436 = _RAND_436[7:0];
  _RAND_437 = {1{`RANDOM}};
  phv_data_437 = _RAND_437[7:0];
  _RAND_438 = {1{`RANDOM}};
  phv_data_438 = _RAND_438[7:0];
  _RAND_439 = {1{`RANDOM}};
  phv_data_439 = _RAND_439[7:0];
  _RAND_440 = {1{`RANDOM}};
  phv_data_440 = _RAND_440[7:0];
  _RAND_441 = {1{`RANDOM}};
  phv_data_441 = _RAND_441[7:0];
  _RAND_442 = {1{`RANDOM}};
  phv_data_442 = _RAND_442[7:0];
  _RAND_443 = {1{`RANDOM}};
  phv_data_443 = _RAND_443[7:0];
  _RAND_444 = {1{`RANDOM}};
  phv_data_444 = _RAND_444[7:0];
  _RAND_445 = {1{`RANDOM}};
  phv_data_445 = _RAND_445[7:0];
  _RAND_446 = {1{`RANDOM}};
  phv_data_446 = _RAND_446[7:0];
  _RAND_447 = {1{`RANDOM}};
  phv_data_447 = _RAND_447[7:0];
  _RAND_448 = {1{`RANDOM}};
  phv_data_448 = _RAND_448[7:0];
  _RAND_449 = {1{`RANDOM}};
  phv_data_449 = _RAND_449[7:0];
  _RAND_450 = {1{`RANDOM}};
  phv_data_450 = _RAND_450[7:0];
  _RAND_451 = {1{`RANDOM}};
  phv_data_451 = _RAND_451[7:0];
  _RAND_452 = {1{`RANDOM}};
  phv_data_452 = _RAND_452[7:0];
  _RAND_453 = {1{`RANDOM}};
  phv_data_453 = _RAND_453[7:0];
  _RAND_454 = {1{`RANDOM}};
  phv_data_454 = _RAND_454[7:0];
  _RAND_455 = {1{`RANDOM}};
  phv_data_455 = _RAND_455[7:0];
  _RAND_456 = {1{`RANDOM}};
  phv_data_456 = _RAND_456[7:0];
  _RAND_457 = {1{`RANDOM}};
  phv_data_457 = _RAND_457[7:0];
  _RAND_458 = {1{`RANDOM}};
  phv_data_458 = _RAND_458[7:0];
  _RAND_459 = {1{`RANDOM}};
  phv_data_459 = _RAND_459[7:0];
  _RAND_460 = {1{`RANDOM}};
  phv_data_460 = _RAND_460[7:0];
  _RAND_461 = {1{`RANDOM}};
  phv_data_461 = _RAND_461[7:0];
  _RAND_462 = {1{`RANDOM}};
  phv_data_462 = _RAND_462[7:0];
  _RAND_463 = {1{`RANDOM}};
  phv_data_463 = _RAND_463[7:0];
  _RAND_464 = {1{`RANDOM}};
  phv_data_464 = _RAND_464[7:0];
  _RAND_465 = {1{`RANDOM}};
  phv_data_465 = _RAND_465[7:0];
  _RAND_466 = {1{`RANDOM}};
  phv_data_466 = _RAND_466[7:0];
  _RAND_467 = {1{`RANDOM}};
  phv_data_467 = _RAND_467[7:0];
  _RAND_468 = {1{`RANDOM}};
  phv_data_468 = _RAND_468[7:0];
  _RAND_469 = {1{`RANDOM}};
  phv_data_469 = _RAND_469[7:0];
  _RAND_470 = {1{`RANDOM}};
  phv_data_470 = _RAND_470[7:0];
  _RAND_471 = {1{`RANDOM}};
  phv_data_471 = _RAND_471[7:0];
  _RAND_472 = {1{`RANDOM}};
  phv_data_472 = _RAND_472[7:0];
  _RAND_473 = {1{`RANDOM}};
  phv_data_473 = _RAND_473[7:0];
  _RAND_474 = {1{`RANDOM}};
  phv_data_474 = _RAND_474[7:0];
  _RAND_475 = {1{`RANDOM}};
  phv_data_475 = _RAND_475[7:0];
  _RAND_476 = {1{`RANDOM}};
  phv_data_476 = _RAND_476[7:0];
  _RAND_477 = {1{`RANDOM}};
  phv_data_477 = _RAND_477[7:0];
  _RAND_478 = {1{`RANDOM}};
  phv_data_478 = _RAND_478[7:0];
  _RAND_479 = {1{`RANDOM}};
  phv_data_479 = _RAND_479[7:0];
  _RAND_480 = {1{`RANDOM}};
  phv_data_480 = _RAND_480[7:0];
  _RAND_481 = {1{`RANDOM}};
  phv_data_481 = _RAND_481[7:0];
  _RAND_482 = {1{`RANDOM}};
  phv_data_482 = _RAND_482[7:0];
  _RAND_483 = {1{`RANDOM}};
  phv_data_483 = _RAND_483[7:0];
  _RAND_484 = {1{`RANDOM}};
  phv_data_484 = _RAND_484[7:0];
  _RAND_485 = {1{`RANDOM}};
  phv_data_485 = _RAND_485[7:0];
  _RAND_486 = {1{`RANDOM}};
  phv_data_486 = _RAND_486[7:0];
  _RAND_487 = {1{`RANDOM}};
  phv_data_487 = _RAND_487[7:0];
  _RAND_488 = {1{`RANDOM}};
  phv_data_488 = _RAND_488[7:0];
  _RAND_489 = {1{`RANDOM}};
  phv_data_489 = _RAND_489[7:0];
  _RAND_490 = {1{`RANDOM}};
  phv_data_490 = _RAND_490[7:0];
  _RAND_491 = {1{`RANDOM}};
  phv_data_491 = _RAND_491[7:0];
  _RAND_492 = {1{`RANDOM}};
  phv_data_492 = _RAND_492[7:0];
  _RAND_493 = {1{`RANDOM}};
  phv_data_493 = _RAND_493[7:0];
  _RAND_494 = {1{`RANDOM}};
  phv_data_494 = _RAND_494[7:0];
  _RAND_495 = {1{`RANDOM}};
  phv_data_495 = _RAND_495[7:0];
  _RAND_496 = {1{`RANDOM}};
  phv_data_496 = _RAND_496[7:0];
  _RAND_497 = {1{`RANDOM}};
  phv_data_497 = _RAND_497[7:0];
  _RAND_498 = {1{`RANDOM}};
  phv_data_498 = _RAND_498[7:0];
  _RAND_499 = {1{`RANDOM}};
  phv_data_499 = _RAND_499[7:0];
  _RAND_500 = {1{`RANDOM}};
  phv_data_500 = _RAND_500[7:0];
  _RAND_501 = {1{`RANDOM}};
  phv_data_501 = _RAND_501[7:0];
  _RAND_502 = {1{`RANDOM}};
  phv_data_502 = _RAND_502[7:0];
  _RAND_503 = {1{`RANDOM}};
  phv_data_503 = _RAND_503[7:0];
  _RAND_504 = {1{`RANDOM}};
  phv_data_504 = _RAND_504[7:0];
  _RAND_505 = {1{`RANDOM}};
  phv_data_505 = _RAND_505[7:0];
  _RAND_506 = {1{`RANDOM}};
  phv_data_506 = _RAND_506[7:0];
  _RAND_507 = {1{`RANDOM}};
  phv_data_507 = _RAND_507[7:0];
  _RAND_508 = {1{`RANDOM}};
  phv_data_508 = _RAND_508[7:0];
  _RAND_509 = {1{`RANDOM}};
  phv_data_509 = _RAND_509[7:0];
  _RAND_510 = {1{`RANDOM}};
  phv_data_510 = _RAND_510[7:0];
  _RAND_511 = {1{`RANDOM}};
  phv_data_511 = _RAND_511[7:0];
  _RAND_512 = {1{`RANDOM}};
  phv_next_processor_id = _RAND_512[3:0];
  _RAND_513 = {1{`RANDOM}};
  phv_next_config_id = _RAND_513[0:0];
  _RAND_514 = {1{`RANDOM}};
  phv_is_valid_processor = _RAND_514[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
