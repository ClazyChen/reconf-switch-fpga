module Controller(
  input         clock,
  input         reset,
  input         io_start,
  input  [7:0]  io_packet_header_0,
  input  [7:0]  io_packet_header_1,
  input  [7:0]  io_packet_header_2,
  input  [7:0]  io_packet_header_3,
  input  [7:0]  io_packet_header_4,
  input  [7:0]  io_packet_header_5,
  input  [7:0]  io_packet_header_6,
  input  [7:0]  io_packet_header_7,
  input  [7:0]  io_packet_header_8,
  input  [7:0]  io_packet_header_9,
  input  [7:0]  io_packet_header_10,
  input  [7:0]  io_packet_header_11,
  input  [7:0]  io_packet_header_12,
  input  [7:0]  io_packet_header_13,
  input  [7:0]  io_packet_header_14,
  input  [7:0]  io_packet_header_15,
  input  [7:0]  io_packet_header_16,
  input  [7:0]  io_packet_header_17,
  input  [7:0]  io_packet_header_18,
  input  [7:0]  io_packet_header_19,
  input  [7:0]  io_packet_header_20,
  input  [7:0]  io_packet_header_21,
  input  [7:0]  io_packet_header_22,
  input  [7:0]  io_packet_header_23,
  input  [7:0]  io_packet_header_24,
  input  [7:0]  io_packet_header_25,
  input  [7:0]  io_packet_header_26,
  input  [7:0]  io_packet_header_27,
  input  [7:0]  io_packet_header_28,
  input  [7:0]  io_packet_header_29,
  input  [7:0]  io_packet_header_30,
  input  [7:0]  io_packet_header_31,
  input  [7:0]  io_packet_header_32,
  input  [7:0]  io_packet_header_33,
  input  [7:0]  io_packet_header_34,
  input  [7:0]  io_packet_header_35,
  input  [7:0]  io_packet_header_36,
  input  [7:0]  io_packet_header_37,
  input  [7:0]  io_packet_header_38,
  input  [7:0]  io_packet_header_39,
  input  [7:0]  io_packet_header_40,
  input  [7:0]  io_packet_header_41,
  input  [7:0]  io_packet_header_42,
  input  [7:0]  io_packet_header_43,
  input  [7:0]  io_packet_header_44,
  input  [7:0]  io_packet_header_45,
  input  [7:0]  io_packet_header_46,
  input  [7:0]  io_packet_header_47,
  input  [7:0]  io_packet_header_48,
  input  [7:0]  io_packet_header_49,
  input  [7:0]  io_packet_header_50,
  input  [7:0]  io_packet_header_51,
  input  [7:0]  io_packet_header_52,
  input  [7:0]  io_packet_header_53,
  input  [7:0]  io_packet_header_54,
  input  [7:0]  io_packet_header_55,
  input  [7:0]  io_packet_header_56,
  input  [7:0]  io_packet_header_57,
  input  [7:0]  io_packet_header_58,
  input  [7:0]  io_packet_header_59,
  input  [7:0]  io_packet_header_60,
  input  [7:0]  io_packet_header_61,
  input  [7:0]  io_packet_header_62,
  input  [7:0]  io_packet_header_63,
  input  [2:0]  io_mod_proc,
  input         io_mod_start,
  input  [31:0] io_mod_hit_action_addr,
  input  [31:0] io_mod_miss_action_addr,
  input         io_mod_ps_mod_start,
  input         io_mod_ps_mod_header_id,
  input  [31:0] io_mod_ps_mod_header_length,
  input  [31:0] io_mod_ps_mod_next_tag_start,
  input  [31:0] io_mod_ps_mod_next_tag_length,
  input  [31:0] io_mod_ps_mod_next_table_0,
  input  [31:0] io_mod_ps_mod_next_table_1,
  input         io_mod_mt_mod_start,
  input  [3:0]  io_mod_mt_mod_header_id,
  input  [5:0]  io_mod_mt_mod_key_off,
  input  [5:0]  io_mod_mt_mod_key_len,
  input  [5:0]  io_mod_mt_mod_val_len,
  input         io_mod_ex_mod_start,
  input  [63:0] io_mod_ex_mod_ops_0,
  input  [63:0] io_mod_ex_mod_ops_1,
  input  [63:0] io_mod_ex_mod_ops_2,
  input  [63:0] io_mod_ex_mod_ops_3,
  input  [63:0] io_mod_ex_mod_ops_4,
  input  [63:0] io_mod_ex_mod_ops_5,
  input  [63:0] io_mod_ex_mod_ops_6,
  input  [63:0] io_mod_ex_mod_ops_7,
  input  [63:0] io_mod_ex_mod_ops_8,
  input  [63:0] io_mod_ex_mod_ops_9,
  input  [63:0] io_mod_ex_mod_ops_10,
  input  [63:0] io_mod_ex_mod_ops_11,
  input  [63:0] io_mod_ex_mod_ops_12,
  input  [63:0] io_mod_ex_mod_ops_13,
  input  [63:0] io_mod_ex_mod_ops_14,
  input  [63:0] io_mod_ex_mod_ops_15,
  output        io_ready_0,
  output        io_ready_1,
  output        io_ready_2,
  output        io_ready_3,
  output        io_ready_4,
  output        io_ready_5,
  output        io_ready_6,
  output        io_ready_7
);
  wire  mem_0_clock; // @[controller.scala 18:25]
  wire [31:0] mem_0_io_mem_a_addr; // @[controller.scala 18:25]
  wire [31:0] mem_0_io_mem_a_rdata; // @[controller.scala 18:25]
  wire [31:0] mem_0_io_mem_b_addr; // @[controller.scala 18:25]
  wire [31:0] mem_0_io_mem_b_rdata; // @[controller.scala 18:25]
  wire  mem_1_clock; // @[controller.scala 18:25]
  wire [31:0] mem_1_io_mem_a_addr; // @[controller.scala 18:25]
  wire [31:0] mem_1_io_mem_a_rdata; // @[controller.scala 18:25]
  wire [31:0] mem_1_io_mem_b_addr; // @[controller.scala 18:25]
  wire [31:0] mem_1_io_mem_b_rdata; // @[controller.scala 18:25]
  wire  mem_2_clock; // @[controller.scala 18:25]
  wire [31:0] mem_2_io_mem_a_addr; // @[controller.scala 18:25]
  wire [31:0] mem_2_io_mem_a_rdata; // @[controller.scala 18:25]
  wire [31:0] mem_2_io_mem_b_addr; // @[controller.scala 18:25]
  wire [31:0] mem_2_io_mem_b_rdata; // @[controller.scala 18:25]
  wire  mem_3_clock; // @[controller.scala 18:25]
  wire [31:0] mem_3_io_mem_a_addr; // @[controller.scala 18:25]
  wire [31:0] mem_3_io_mem_a_rdata; // @[controller.scala 18:25]
  wire [31:0] mem_3_io_mem_b_addr; // @[controller.scala 18:25]
  wire [31:0] mem_3_io_mem_b_rdata; // @[controller.scala 18:25]
  wire [7:0] encoders_0_io_input; // @[controller.scala 23:25]
  wire [2:0] encoders_0_io_output; // @[controller.scala 23:25]
  wire  encoders_0_io_valid; // @[controller.scala 23:25]
  wire [7:0] encoders_1_io_input; // @[controller.scala 23:25]
  wire [2:0] encoders_1_io_output; // @[controller.scala 23:25]
  wire  encoders_1_io_valid; // @[controller.scala 23:25]
  wire [7:0] encoders_2_io_input; // @[controller.scala 23:25]
  wire [2:0] encoders_2_io_output; // @[controller.scala 23:25]
  wire  encoders_2_io_valid; // @[controller.scala 23:25]
  wire [7:0] encoders_3_io_input; // @[controller.scala 23:25]
  wire [2:0] encoders_3_io_output; // @[controller.scala 23:25]
  wire  encoders_3_io_valid; // @[controller.scala 23:25]
  wire [7:0] encoders_4_io_input; // @[controller.scala 23:25]
  wire [2:0] encoders_4_io_output; // @[controller.scala 23:25]
  wire  encoders_4_io_valid; // @[controller.scala 23:25]
  wire [7:0] encoders_5_io_input; // @[controller.scala 23:25]
  wire [2:0] encoders_5_io_output; // @[controller.scala 23:25]
  wire  encoders_5_io_valid; // @[controller.scala 23:25]
  wire [7:0] encoders_6_io_input; // @[controller.scala 23:25]
  wire [2:0] encoders_6_io_output; // @[controller.scala 23:25]
  wire  encoders_6_io_valid; // @[controller.scala 23:25]
  wire [7:0] encoders_7_io_input; // @[controller.scala 23:25]
  wire [2:0] encoders_7_io_output; // @[controller.scala 23:25]
  wire  encoders_7_io_valid; // @[controller.scala 23:25]
  wire  proc_0_clock; // @[controller.scala 29:25]
  wire  proc_0_reset; // @[controller.scala 29:25]
  wire  proc_0_io_update; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_packet_header_0; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_packet_header_1; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_packet_header_2; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_packet_header_3; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_packet_header_4; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_packet_header_5; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_packet_header_6; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_packet_header_7; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_packet_header_8; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_packet_header_9; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_packet_header_10; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_packet_header_11; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_packet_header_12; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_packet_header_13; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_packet_header_14; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_packet_header_15; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_packet_header_16; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_packet_header_17; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_packet_header_18; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_packet_header_19; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_packet_header_20; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_packet_header_21; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_packet_header_22; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_packet_header_23; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_packet_header_24; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_packet_header_25; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_packet_header_26; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_packet_header_27; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_packet_header_28; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_packet_header_29; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_packet_header_30; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_packet_header_31; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_packet_header_32; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_packet_header_33; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_packet_header_34; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_packet_header_35; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_packet_header_36; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_packet_header_37; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_packet_header_38; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_packet_header_39; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_packet_header_40; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_packet_header_41; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_packet_header_42; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_packet_header_43; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_packet_header_44; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_packet_header_45; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_packet_header_46; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_packet_header_47; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_packet_header_48; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_packet_header_49; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_packet_header_50; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_packet_header_51; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_packet_header_52; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_packet_header_53; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_packet_header_54; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_packet_header_55; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_packet_header_56; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_packet_header_57; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_packet_header_58; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_packet_header_59; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_packet_header_60; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_packet_header_61; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_packet_header_62; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_packet_header_63; // @[controller.scala 29:25]
  wire  proc_0_io_end; // @[controller.scala 29:25]
  wire [31:0] proc_0_io_mem_addr; // @[controller.scala 29:25]
  wire [31:0] proc_0_io_mem_rdata; // @[controller.scala 29:25]
  wire  proc_0_io_ready; // @[controller.scala 29:25]
  wire  proc_0_io_mod_start; // @[controller.scala 29:25]
  wire [31:0] proc_0_io_mod_hit_action_addr; // @[controller.scala 29:25]
  wire [31:0] proc_0_io_mod_miss_action_addr; // @[controller.scala 29:25]
  wire  proc_0_io_mod_ps_mod_start; // @[controller.scala 29:25]
  wire  proc_0_io_mod_ps_mod_header_id; // @[controller.scala 29:25]
  wire [31:0] proc_0_io_mod_ps_mod_header_length; // @[controller.scala 29:25]
  wire [31:0] proc_0_io_mod_ps_mod_next_tag_start; // @[controller.scala 29:25]
  wire [31:0] proc_0_io_mod_ps_mod_next_table_0; // @[controller.scala 29:25]
  wire [31:0] proc_0_io_mod_ps_mod_next_table_1; // @[controller.scala 29:25]
  wire  proc_0_io_mod_mt_mod_start; // @[controller.scala 29:25]
  wire [3:0] proc_0_io_mod_mt_mod_header_id; // @[controller.scala 29:25]
  wire [5:0] proc_0_io_mod_mt_mod_key_off; // @[controller.scala 29:25]
  wire [5:0] proc_0_io_mod_mt_mod_key_len; // @[controller.scala 29:25]
  wire [5:0] proc_0_io_mod_mt_mod_val_len; // @[controller.scala 29:25]
  wire  proc_0_io_mod_ex_mod_start; // @[controller.scala 29:25]
  wire [63:0] proc_0_io_mod_ex_mod_ops_0; // @[controller.scala 29:25]
  wire [63:0] proc_0_io_mod_ex_mod_ops_1; // @[controller.scala 29:25]
  wire [63:0] proc_0_io_mod_ex_mod_ops_2; // @[controller.scala 29:25]
  wire [63:0] proc_0_io_mod_ex_mod_ops_3; // @[controller.scala 29:25]
  wire [63:0] proc_0_io_mod_ex_mod_ops_4; // @[controller.scala 29:25]
  wire [63:0] proc_0_io_mod_ex_mod_ops_5; // @[controller.scala 29:25]
  wire [63:0] proc_0_io_mod_ex_mod_ops_6; // @[controller.scala 29:25]
  wire [63:0] proc_0_io_mod_ex_mod_ops_7; // @[controller.scala 29:25]
  wire [63:0] proc_0_io_mod_ex_mod_ops_8; // @[controller.scala 29:25]
  wire [63:0] proc_0_io_mod_ex_mod_ops_9; // @[controller.scala 29:25]
  wire [63:0] proc_0_io_mod_ex_mod_ops_10; // @[controller.scala 29:25]
  wire [63:0] proc_0_io_mod_ex_mod_ops_11; // @[controller.scala 29:25]
  wire [63:0] proc_0_io_mod_ex_mod_ops_12; // @[controller.scala 29:25]
  wire [63:0] proc_0_io_mod_ex_mod_ops_13; // @[controller.scala 29:25]
  wire [63:0] proc_0_io_mod_ex_mod_ops_14; // @[controller.scala 29:25]
  wire [63:0] proc_0_io_mod_ex_mod_ops_15; // @[controller.scala 29:25]
  wire  proc_0_io_next_en; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_next_header_0; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_next_header_1; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_next_header_2; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_next_header_3; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_next_header_4; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_next_header_5; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_next_header_6; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_next_header_7; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_next_header_8; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_next_header_9; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_next_header_10; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_next_header_11; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_next_header_12; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_next_header_13; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_next_header_14; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_next_header_15; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_next_header_16; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_next_header_17; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_next_header_18; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_next_header_19; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_next_header_20; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_next_header_21; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_next_header_22; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_next_header_23; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_next_header_24; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_next_header_25; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_next_header_26; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_next_header_27; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_next_header_28; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_next_header_29; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_next_header_30; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_next_header_31; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_next_header_32; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_next_header_33; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_next_header_34; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_next_header_35; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_next_header_36; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_next_header_37; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_next_header_38; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_next_header_39; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_next_header_40; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_next_header_41; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_next_header_42; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_next_header_43; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_next_header_44; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_next_header_45; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_next_header_46; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_next_header_47; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_next_header_48; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_next_header_49; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_next_header_50; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_next_header_51; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_next_header_52; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_next_header_53; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_next_header_54; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_next_header_55; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_next_header_56; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_next_header_57; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_next_header_58; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_next_header_59; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_next_header_60; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_next_header_61; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_next_header_62; // @[controller.scala 29:25]
  wire [7:0] proc_0_io_next_header_63; // @[controller.scala 29:25]
  wire [2:0] proc_0_io_next_proc; // @[controller.scala 29:25]
  wire  proc_1_clock; // @[controller.scala 29:25]
  wire  proc_1_reset; // @[controller.scala 29:25]
  wire  proc_1_io_update; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_packet_header_0; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_packet_header_1; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_packet_header_2; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_packet_header_3; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_packet_header_4; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_packet_header_5; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_packet_header_6; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_packet_header_7; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_packet_header_8; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_packet_header_9; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_packet_header_10; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_packet_header_11; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_packet_header_12; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_packet_header_13; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_packet_header_14; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_packet_header_15; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_packet_header_16; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_packet_header_17; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_packet_header_18; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_packet_header_19; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_packet_header_20; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_packet_header_21; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_packet_header_22; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_packet_header_23; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_packet_header_24; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_packet_header_25; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_packet_header_26; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_packet_header_27; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_packet_header_28; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_packet_header_29; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_packet_header_30; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_packet_header_31; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_packet_header_32; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_packet_header_33; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_packet_header_34; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_packet_header_35; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_packet_header_36; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_packet_header_37; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_packet_header_38; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_packet_header_39; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_packet_header_40; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_packet_header_41; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_packet_header_42; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_packet_header_43; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_packet_header_44; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_packet_header_45; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_packet_header_46; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_packet_header_47; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_packet_header_48; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_packet_header_49; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_packet_header_50; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_packet_header_51; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_packet_header_52; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_packet_header_53; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_packet_header_54; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_packet_header_55; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_packet_header_56; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_packet_header_57; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_packet_header_58; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_packet_header_59; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_packet_header_60; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_packet_header_61; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_packet_header_62; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_packet_header_63; // @[controller.scala 29:25]
  wire  proc_1_io_end; // @[controller.scala 29:25]
  wire [31:0] proc_1_io_mem_addr; // @[controller.scala 29:25]
  wire [31:0] proc_1_io_mem_rdata; // @[controller.scala 29:25]
  wire  proc_1_io_ready; // @[controller.scala 29:25]
  wire  proc_1_io_mod_start; // @[controller.scala 29:25]
  wire [31:0] proc_1_io_mod_hit_action_addr; // @[controller.scala 29:25]
  wire [31:0] proc_1_io_mod_miss_action_addr; // @[controller.scala 29:25]
  wire  proc_1_io_mod_ps_mod_start; // @[controller.scala 29:25]
  wire  proc_1_io_mod_ps_mod_header_id; // @[controller.scala 29:25]
  wire [31:0] proc_1_io_mod_ps_mod_header_length; // @[controller.scala 29:25]
  wire [31:0] proc_1_io_mod_ps_mod_next_tag_start; // @[controller.scala 29:25]
  wire [31:0] proc_1_io_mod_ps_mod_next_table_0; // @[controller.scala 29:25]
  wire [31:0] proc_1_io_mod_ps_mod_next_table_1; // @[controller.scala 29:25]
  wire  proc_1_io_mod_mt_mod_start; // @[controller.scala 29:25]
  wire [3:0] proc_1_io_mod_mt_mod_header_id; // @[controller.scala 29:25]
  wire [5:0] proc_1_io_mod_mt_mod_key_off; // @[controller.scala 29:25]
  wire [5:0] proc_1_io_mod_mt_mod_key_len; // @[controller.scala 29:25]
  wire [5:0] proc_1_io_mod_mt_mod_val_len; // @[controller.scala 29:25]
  wire  proc_1_io_mod_ex_mod_start; // @[controller.scala 29:25]
  wire [63:0] proc_1_io_mod_ex_mod_ops_0; // @[controller.scala 29:25]
  wire [63:0] proc_1_io_mod_ex_mod_ops_1; // @[controller.scala 29:25]
  wire [63:0] proc_1_io_mod_ex_mod_ops_2; // @[controller.scala 29:25]
  wire [63:0] proc_1_io_mod_ex_mod_ops_3; // @[controller.scala 29:25]
  wire [63:0] proc_1_io_mod_ex_mod_ops_4; // @[controller.scala 29:25]
  wire [63:0] proc_1_io_mod_ex_mod_ops_5; // @[controller.scala 29:25]
  wire [63:0] proc_1_io_mod_ex_mod_ops_6; // @[controller.scala 29:25]
  wire [63:0] proc_1_io_mod_ex_mod_ops_7; // @[controller.scala 29:25]
  wire [63:0] proc_1_io_mod_ex_mod_ops_8; // @[controller.scala 29:25]
  wire [63:0] proc_1_io_mod_ex_mod_ops_9; // @[controller.scala 29:25]
  wire [63:0] proc_1_io_mod_ex_mod_ops_10; // @[controller.scala 29:25]
  wire [63:0] proc_1_io_mod_ex_mod_ops_11; // @[controller.scala 29:25]
  wire [63:0] proc_1_io_mod_ex_mod_ops_12; // @[controller.scala 29:25]
  wire [63:0] proc_1_io_mod_ex_mod_ops_13; // @[controller.scala 29:25]
  wire [63:0] proc_1_io_mod_ex_mod_ops_14; // @[controller.scala 29:25]
  wire [63:0] proc_1_io_mod_ex_mod_ops_15; // @[controller.scala 29:25]
  wire  proc_1_io_next_en; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_next_header_0; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_next_header_1; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_next_header_2; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_next_header_3; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_next_header_4; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_next_header_5; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_next_header_6; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_next_header_7; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_next_header_8; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_next_header_9; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_next_header_10; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_next_header_11; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_next_header_12; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_next_header_13; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_next_header_14; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_next_header_15; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_next_header_16; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_next_header_17; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_next_header_18; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_next_header_19; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_next_header_20; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_next_header_21; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_next_header_22; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_next_header_23; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_next_header_24; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_next_header_25; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_next_header_26; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_next_header_27; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_next_header_28; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_next_header_29; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_next_header_30; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_next_header_31; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_next_header_32; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_next_header_33; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_next_header_34; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_next_header_35; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_next_header_36; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_next_header_37; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_next_header_38; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_next_header_39; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_next_header_40; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_next_header_41; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_next_header_42; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_next_header_43; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_next_header_44; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_next_header_45; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_next_header_46; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_next_header_47; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_next_header_48; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_next_header_49; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_next_header_50; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_next_header_51; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_next_header_52; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_next_header_53; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_next_header_54; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_next_header_55; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_next_header_56; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_next_header_57; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_next_header_58; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_next_header_59; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_next_header_60; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_next_header_61; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_next_header_62; // @[controller.scala 29:25]
  wire [7:0] proc_1_io_next_header_63; // @[controller.scala 29:25]
  wire [2:0] proc_1_io_next_proc; // @[controller.scala 29:25]
  wire  proc_2_clock; // @[controller.scala 29:25]
  wire  proc_2_reset; // @[controller.scala 29:25]
  wire  proc_2_io_update; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_packet_header_0; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_packet_header_1; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_packet_header_2; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_packet_header_3; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_packet_header_4; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_packet_header_5; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_packet_header_6; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_packet_header_7; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_packet_header_8; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_packet_header_9; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_packet_header_10; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_packet_header_11; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_packet_header_12; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_packet_header_13; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_packet_header_14; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_packet_header_15; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_packet_header_16; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_packet_header_17; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_packet_header_18; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_packet_header_19; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_packet_header_20; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_packet_header_21; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_packet_header_22; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_packet_header_23; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_packet_header_24; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_packet_header_25; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_packet_header_26; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_packet_header_27; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_packet_header_28; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_packet_header_29; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_packet_header_30; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_packet_header_31; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_packet_header_32; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_packet_header_33; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_packet_header_34; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_packet_header_35; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_packet_header_36; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_packet_header_37; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_packet_header_38; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_packet_header_39; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_packet_header_40; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_packet_header_41; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_packet_header_42; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_packet_header_43; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_packet_header_44; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_packet_header_45; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_packet_header_46; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_packet_header_47; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_packet_header_48; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_packet_header_49; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_packet_header_50; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_packet_header_51; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_packet_header_52; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_packet_header_53; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_packet_header_54; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_packet_header_55; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_packet_header_56; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_packet_header_57; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_packet_header_58; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_packet_header_59; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_packet_header_60; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_packet_header_61; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_packet_header_62; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_packet_header_63; // @[controller.scala 29:25]
  wire  proc_2_io_end; // @[controller.scala 29:25]
  wire [31:0] proc_2_io_mem_addr; // @[controller.scala 29:25]
  wire [31:0] proc_2_io_mem_rdata; // @[controller.scala 29:25]
  wire  proc_2_io_ready; // @[controller.scala 29:25]
  wire  proc_2_io_mod_start; // @[controller.scala 29:25]
  wire [31:0] proc_2_io_mod_hit_action_addr; // @[controller.scala 29:25]
  wire [31:0] proc_2_io_mod_miss_action_addr; // @[controller.scala 29:25]
  wire  proc_2_io_mod_ps_mod_start; // @[controller.scala 29:25]
  wire  proc_2_io_mod_ps_mod_header_id; // @[controller.scala 29:25]
  wire [31:0] proc_2_io_mod_ps_mod_header_length; // @[controller.scala 29:25]
  wire [31:0] proc_2_io_mod_ps_mod_next_tag_start; // @[controller.scala 29:25]
  wire [31:0] proc_2_io_mod_ps_mod_next_table_0; // @[controller.scala 29:25]
  wire [31:0] proc_2_io_mod_ps_mod_next_table_1; // @[controller.scala 29:25]
  wire  proc_2_io_mod_mt_mod_start; // @[controller.scala 29:25]
  wire [3:0] proc_2_io_mod_mt_mod_header_id; // @[controller.scala 29:25]
  wire [5:0] proc_2_io_mod_mt_mod_key_off; // @[controller.scala 29:25]
  wire [5:0] proc_2_io_mod_mt_mod_key_len; // @[controller.scala 29:25]
  wire [5:0] proc_2_io_mod_mt_mod_val_len; // @[controller.scala 29:25]
  wire  proc_2_io_mod_ex_mod_start; // @[controller.scala 29:25]
  wire [63:0] proc_2_io_mod_ex_mod_ops_0; // @[controller.scala 29:25]
  wire [63:0] proc_2_io_mod_ex_mod_ops_1; // @[controller.scala 29:25]
  wire [63:0] proc_2_io_mod_ex_mod_ops_2; // @[controller.scala 29:25]
  wire [63:0] proc_2_io_mod_ex_mod_ops_3; // @[controller.scala 29:25]
  wire [63:0] proc_2_io_mod_ex_mod_ops_4; // @[controller.scala 29:25]
  wire [63:0] proc_2_io_mod_ex_mod_ops_5; // @[controller.scala 29:25]
  wire [63:0] proc_2_io_mod_ex_mod_ops_6; // @[controller.scala 29:25]
  wire [63:0] proc_2_io_mod_ex_mod_ops_7; // @[controller.scala 29:25]
  wire [63:0] proc_2_io_mod_ex_mod_ops_8; // @[controller.scala 29:25]
  wire [63:0] proc_2_io_mod_ex_mod_ops_9; // @[controller.scala 29:25]
  wire [63:0] proc_2_io_mod_ex_mod_ops_10; // @[controller.scala 29:25]
  wire [63:0] proc_2_io_mod_ex_mod_ops_11; // @[controller.scala 29:25]
  wire [63:0] proc_2_io_mod_ex_mod_ops_12; // @[controller.scala 29:25]
  wire [63:0] proc_2_io_mod_ex_mod_ops_13; // @[controller.scala 29:25]
  wire [63:0] proc_2_io_mod_ex_mod_ops_14; // @[controller.scala 29:25]
  wire [63:0] proc_2_io_mod_ex_mod_ops_15; // @[controller.scala 29:25]
  wire  proc_2_io_next_en; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_next_header_0; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_next_header_1; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_next_header_2; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_next_header_3; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_next_header_4; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_next_header_5; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_next_header_6; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_next_header_7; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_next_header_8; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_next_header_9; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_next_header_10; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_next_header_11; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_next_header_12; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_next_header_13; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_next_header_14; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_next_header_15; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_next_header_16; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_next_header_17; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_next_header_18; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_next_header_19; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_next_header_20; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_next_header_21; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_next_header_22; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_next_header_23; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_next_header_24; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_next_header_25; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_next_header_26; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_next_header_27; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_next_header_28; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_next_header_29; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_next_header_30; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_next_header_31; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_next_header_32; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_next_header_33; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_next_header_34; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_next_header_35; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_next_header_36; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_next_header_37; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_next_header_38; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_next_header_39; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_next_header_40; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_next_header_41; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_next_header_42; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_next_header_43; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_next_header_44; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_next_header_45; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_next_header_46; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_next_header_47; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_next_header_48; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_next_header_49; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_next_header_50; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_next_header_51; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_next_header_52; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_next_header_53; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_next_header_54; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_next_header_55; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_next_header_56; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_next_header_57; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_next_header_58; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_next_header_59; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_next_header_60; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_next_header_61; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_next_header_62; // @[controller.scala 29:25]
  wire [7:0] proc_2_io_next_header_63; // @[controller.scala 29:25]
  wire [2:0] proc_2_io_next_proc; // @[controller.scala 29:25]
  wire  proc_3_clock; // @[controller.scala 29:25]
  wire  proc_3_reset; // @[controller.scala 29:25]
  wire  proc_3_io_update; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_packet_header_0; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_packet_header_1; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_packet_header_2; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_packet_header_3; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_packet_header_4; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_packet_header_5; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_packet_header_6; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_packet_header_7; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_packet_header_8; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_packet_header_9; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_packet_header_10; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_packet_header_11; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_packet_header_12; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_packet_header_13; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_packet_header_14; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_packet_header_15; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_packet_header_16; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_packet_header_17; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_packet_header_18; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_packet_header_19; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_packet_header_20; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_packet_header_21; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_packet_header_22; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_packet_header_23; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_packet_header_24; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_packet_header_25; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_packet_header_26; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_packet_header_27; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_packet_header_28; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_packet_header_29; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_packet_header_30; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_packet_header_31; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_packet_header_32; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_packet_header_33; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_packet_header_34; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_packet_header_35; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_packet_header_36; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_packet_header_37; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_packet_header_38; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_packet_header_39; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_packet_header_40; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_packet_header_41; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_packet_header_42; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_packet_header_43; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_packet_header_44; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_packet_header_45; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_packet_header_46; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_packet_header_47; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_packet_header_48; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_packet_header_49; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_packet_header_50; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_packet_header_51; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_packet_header_52; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_packet_header_53; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_packet_header_54; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_packet_header_55; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_packet_header_56; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_packet_header_57; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_packet_header_58; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_packet_header_59; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_packet_header_60; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_packet_header_61; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_packet_header_62; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_packet_header_63; // @[controller.scala 29:25]
  wire  proc_3_io_end; // @[controller.scala 29:25]
  wire [31:0] proc_3_io_mem_addr; // @[controller.scala 29:25]
  wire [31:0] proc_3_io_mem_rdata; // @[controller.scala 29:25]
  wire  proc_3_io_ready; // @[controller.scala 29:25]
  wire  proc_3_io_mod_start; // @[controller.scala 29:25]
  wire [31:0] proc_3_io_mod_hit_action_addr; // @[controller.scala 29:25]
  wire [31:0] proc_3_io_mod_miss_action_addr; // @[controller.scala 29:25]
  wire  proc_3_io_mod_ps_mod_start; // @[controller.scala 29:25]
  wire  proc_3_io_mod_ps_mod_header_id; // @[controller.scala 29:25]
  wire [31:0] proc_3_io_mod_ps_mod_header_length; // @[controller.scala 29:25]
  wire [31:0] proc_3_io_mod_ps_mod_next_tag_start; // @[controller.scala 29:25]
  wire [31:0] proc_3_io_mod_ps_mod_next_table_0; // @[controller.scala 29:25]
  wire [31:0] proc_3_io_mod_ps_mod_next_table_1; // @[controller.scala 29:25]
  wire  proc_3_io_mod_mt_mod_start; // @[controller.scala 29:25]
  wire [3:0] proc_3_io_mod_mt_mod_header_id; // @[controller.scala 29:25]
  wire [5:0] proc_3_io_mod_mt_mod_key_off; // @[controller.scala 29:25]
  wire [5:0] proc_3_io_mod_mt_mod_key_len; // @[controller.scala 29:25]
  wire [5:0] proc_3_io_mod_mt_mod_val_len; // @[controller.scala 29:25]
  wire  proc_3_io_mod_ex_mod_start; // @[controller.scala 29:25]
  wire [63:0] proc_3_io_mod_ex_mod_ops_0; // @[controller.scala 29:25]
  wire [63:0] proc_3_io_mod_ex_mod_ops_1; // @[controller.scala 29:25]
  wire [63:0] proc_3_io_mod_ex_mod_ops_2; // @[controller.scala 29:25]
  wire [63:0] proc_3_io_mod_ex_mod_ops_3; // @[controller.scala 29:25]
  wire [63:0] proc_3_io_mod_ex_mod_ops_4; // @[controller.scala 29:25]
  wire [63:0] proc_3_io_mod_ex_mod_ops_5; // @[controller.scala 29:25]
  wire [63:0] proc_3_io_mod_ex_mod_ops_6; // @[controller.scala 29:25]
  wire [63:0] proc_3_io_mod_ex_mod_ops_7; // @[controller.scala 29:25]
  wire [63:0] proc_3_io_mod_ex_mod_ops_8; // @[controller.scala 29:25]
  wire [63:0] proc_3_io_mod_ex_mod_ops_9; // @[controller.scala 29:25]
  wire [63:0] proc_3_io_mod_ex_mod_ops_10; // @[controller.scala 29:25]
  wire [63:0] proc_3_io_mod_ex_mod_ops_11; // @[controller.scala 29:25]
  wire [63:0] proc_3_io_mod_ex_mod_ops_12; // @[controller.scala 29:25]
  wire [63:0] proc_3_io_mod_ex_mod_ops_13; // @[controller.scala 29:25]
  wire [63:0] proc_3_io_mod_ex_mod_ops_14; // @[controller.scala 29:25]
  wire [63:0] proc_3_io_mod_ex_mod_ops_15; // @[controller.scala 29:25]
  wire  proc_3_io_next_en; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_next_header_0; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_next_header_1; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_next_header_2; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_next_header_3; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_next_header_4; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_next_header_5; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_next_header_6; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_next_header_7; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_next_header_8; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_next_header_9; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_next_header_10; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_next_header_11; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_next_header_12; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_next_header_13; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_next_header_14; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_next_header_15; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_next_header_16; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_next_header_17; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_next_header_18; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_next_header_19; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_next_header_20; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_next_header_21; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_next_header_22; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_next_header_23; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_next_header_24; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_next_header_25; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_next_header_26; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_next_header_27; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_next_header_28; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_next_header_29; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_next_header_30; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_next_header_31; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_next_header_32; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_next_header_33; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_next_header_34; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_next_header_35; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_next_header_36; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_next_header_37; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_next_header_38; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_next_header_39; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_next_header_40; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_next_header_41; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_next_header_42; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_next_header_43; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_next_header_44; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_next_header_45; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_next_header_46; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_next_header_47; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_next_header_48; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_next_header_49; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_next_header_50; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_next_header_51; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_next_header_52; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_next_header_53; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_next_header_54; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_next_header_55; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_next_header_56; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_next_header_57; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_next_header_58; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_next_header_59; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_next_header_60; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_next_header_61; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_next_header_62; // @[controller.scala 29:25]
  wire [7:0] proc_3_io_next_header_63; // @[controller.scala 29:25]
  wire [2:0] proc_3_io_next_proc; // @[controller.scala 29:25]
  wire  proc_4_clock; // @[controller.scala 29:25]
  wire  proc_4_reset; // @[controller.scala 29:25]
  wire  proc_4_io_update; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_packet_header_0; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_packet_header_1; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_packet_header_2; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_packet_header_3; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_packet_header_4; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_packet_header_5; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_packet_header_6; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_packet_header_7; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_packet_header_8; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_packet_header_9; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_packet_header_10; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_packet_header_11; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_packet_header_12; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_packet_header_13; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_packet_header_14; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_packet_header_15; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_packet_header_16; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_packet_header_17; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_packet_header_18; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_packet_header_19; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_packet_header_20; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_packet_header_21; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_packet_header_22; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_packet_header_23; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_packet_header_24; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_packet_header_25; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_packet_header_26; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_packet_header_27; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_packet_header_28; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_packet_header_29; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_packet_header_30; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_packet_header_31; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_packet_header_32; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_packet_header_33; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_packet_header_34; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_packet_header_35; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_packet_header_36; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_packet_header_37; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_packet_header_38; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_packet_header_39; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_packet_header_40; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_packet_header_41; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_packet_header_42; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_packet_header_43; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_packet_header_44; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_packet_header_45; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_packet_header_46; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_packet_header_47; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_packet_header_48; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_packet_header_49; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_packet_header_50; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_packet_header_51; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_packet_header_52; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_packet_header_53; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_packet_header_54; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_packet_header_55; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_packet_header_56; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_packet_header_57; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_packet_header_58; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_packet_header_59; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_packet_header_60; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_packet_header_61; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_packet_header_62; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_packet_header_63; // @[controller.scala 29:25]
  wire  proc_4_io_end; // @[controller.scala 29:25]
  wire [31:0] proc_4_io_mem_addr; // @[controller.scala 29:25]
  wire [31:0] proc_4_io_mem_rdata; // @[controller.scala 29:25]
  wire  proc_4_io_ready; // @[controller.scala 29:25]
  wire  proc_4_io_mod_start; // @[controller.scala 29:25]
  wire [31:0] proc_4_io_mod_hit_action_addr; // @[controller.scala 29:25]
  wire [31:0] proc_4_io_mod_miss_action_addr; // @[controller.scala 29:25]
  wire  proc_4_io_mod_ps_mod_start; // @[controller.scala 29:25]
  wire  proc_4_io_mod_ps_mod_header_id; // @[controller.scala 29:25]
  wire [31:0] proc_4_io_mod_ps_mod_header_length; // @[controller.scala 29:25]
  wire [31:0] proc_4_io_mod_ps_mod_next_tag_start; // @[controller.scala 29:25]
  wire [31:0] proc_4_io_mod_ps_mod_next_table_0; // @[controller.scala 29:25]
  wire [31:0] proc_4_io_mod_ps_mod_next_table_1; // @[controller.scala 29:25]
  wire  proc_4_io_mod_mt_mod_start; // @[controller.scala 29:25]
  wire [3:0] proc_4_io_mod_mt_mod_header_id; // @[controller.scala 29:25]
  wire [5:0] proc_4_io_mod_mt_mod_key_off; // @[controller.scala 29:25]
  wire [5:0] proc_4_io_mod_mt_mod_key_len; // @[controller.scala 29:25]
  wire [5:0] proc_4_io_mod_mt_mod_val_len; // @[controller.scala 29:25]
  wire  proc_4_io_mod_ex_mod_start; // @[controller.scala 29:25]
  wire [63:0] proc_4_io_mod_ex_mod_ops_0; // @[controller.scala 29:25]
  wire [63:0] proc_4_io_mod_ex_mod_ops_1; // @[controller.scala 29:25]
  wire [63:0] proc_4_io_mod_ex_mod_ops_2; // @[controller.scala 29:25]
  wire [63:0] proc_4_io_mod_ex_mod_ops_3; // @[controller.scala 29:25]
  wire [63:0] proc_4_io_mod_ex_mod_ops_4; // @[controller.scala 29:25]
  wire [63:0] proc_4_io_mod_ex_mod_ops_5; // @[controller.scala 29:25]
  wire [63:0] proc_4_io_mod_ex_mod_ops_6; // @[controller.scala 29:25]
  wire [63:0] proc_4_io_mod_ex_mod_ops_7; // @[controller.scala 29:25]
  wire [63:0] proc_4_io_mod_ex_mod_ops_8; // @[controller.scala 29:25]
  wire [63:0] proc_4_io_mod_ex_mod_ops_9; // @[controller.scala 29:25]
  wire [63:0] proc_4_io_mod_ex_mod_ops_10; // @[controller.scala 29:25]
  wire [63:0] proc_4_io_mod_ex_mod_ops_11; // @[controller.scala 29:25]
  wire [63:0] proc_4_io_mod_ex_mod_ops_12; // @[controller.scala 29:25]
  wire [63:0] proc_4_io_mod_ex_mod_ops_13; // @[controller.scala 29:25]
  wire [63:0] proc_4_io_mod_ex_mod_ops_14; // @[controller.scala 29:25]
  wire [63:0] proc_4_io_mod_ex_mod_ops_15; // @[controller.scala 29:25]
  wire  proc_4_io_next_en; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_next_header_0; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_next_header_1; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_next_header_2; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_next_header_3; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_next_header_4; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_next_header_5; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_next_header_6; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_next_header_7; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_next_header_8; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_next_header_9; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_next_header_10; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_next_header_11; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_next_header_12; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_next_header_13; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_next_header_14; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_next_header_15; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_next_header_16; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_next_header_17; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_next_header_18; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_next_header_19; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_next_header_20; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_next_header_21; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_next_header_22; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_next_header_23; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_next_header_24; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_next_header_25; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_next_header_26; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_next_header_27; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_next_header_28; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_next_header_29; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_next_header_30; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_next_header_31; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_next_header_32; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_next_header_33; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_next_header_34; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_next_header_35; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_next_header_36; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_next_header_37; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_next_header_38; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_next_header_39; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_next_header_40; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_next_header_41; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_next_header_42; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_next_header_43; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_next_header_44; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_next_header_45; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_next_header_46; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_next_header_47; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_next_header_48; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_next_header_49; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_next_header_50; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_next_header_51; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_next_header_52; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_next_header_53; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_next_header_54; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_next_header_55; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_next_header_56; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_next_header_57; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_next_header_58; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_next_header_59; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_next_header_60; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_next_header_61; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_next_header_62; // @[controller.scala 29:25]
  wire [7:0] proc_4_io_next_header_63; // @[controller.scala 29:25]
  wire [2:0] proc_4_io_next_proc; // @[controller.scala 29:25]
  wire  proc_5_clock; // @[controller.scala 29:25]
  wire  proc_5_reset; // @[controller.scala 29:25]
  wire  proc_5_io_update; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_packet_header_0; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_packet_header_1; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_packet_header_2; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_packet_header_3; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_packet_header_4; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_packet_header_5; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_packet_header_6; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_packet_header_7; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_packet_header_8; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_packet_header_9; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_packet_header_10; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_packet_header_11; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_packet_header_12; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_packet_header_13; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_packet_header_14; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_packet_header_15; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_packet_header_16; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_packet_header_17; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_packet_header_18; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_packet_header_19; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_packet_header_20; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_packet_header_21; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_packet_header_22; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_packet_header_23; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_packet_header_24; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_packet_header_25; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_packet_header_26; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_packet_header_27; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_packet_header_28; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_packet_header_29; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_packet_header_30; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_packet_header_31; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_packet_header_32; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_packet_header_33; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_packet_header_34; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_packet_header_35; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_packet_header_36; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_packet_header_37; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_packet_header_38; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_packet_header_39; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_packet_header_40; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_packet_header_41; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_packet_header_42; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_packet_header_43; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_packet_header_44; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_packet_header_45; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_packet_header_46; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_packet_header_47; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_packet_header_48; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_packet_header_49; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_packet_header_50; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_packet_header_51; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_packet_header_52; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_packet_header_53; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_packet_header_54; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_packet_header_55; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_packet_header_56; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_packet_header_57; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_packet_header_58; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_packet_header_59; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_packet_header_60; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_packet_header_61; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_packet_header_62; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_packet_header_63; // @[controller.scala 29:25]
  wire  proc_5_io_end; // @[controller.scala 29:25]
  wire [31:0] proc_5_io_mem_addr; // @[controller.scala 29:25]
  wire [31:0] proc_5_io_mem_rdata; // @[controller.scala 29:25]
  wire  proc_5_io_ready; // @[controller.scala 29:25]
  wire  proc_5_io_mod_start; // @[controller.scala 29:25]
  wire [31:0] proc_5_io_mod_hit_action_addr; // @[controller.scala 29:25]
  wire [31:0] proc_5_io_mod_miss_action_addr; // @[controller.scala 29:25]
  wire  proc_5_io_mod_ps_mod_start; // @[controller.scala 29:25]
  wire  proc_5_io_mod_ps_mod_header_id; // @[controller.scala 29:25]
  wire [31:0] proc_5_io_mod_ps_mod_header_length; // @[controller.scala 29:25]
  wire [31:0] proc_5_io_mod_ps_mod_next_tag_start; // @[controller.scala 29:25]
  wire [31:0] proc_5_io_mod_ps_mod_next_table_0; // @[controller.scala 29:25]
  wire [31:0] proc_5_io_mod_ps_mod_next_table_1; // @[controller.scala 29:25]
  wire  proc_5_io_mod_mt_mod_start; // @[controller.scala 29:25]
  wire [3:0] proc_5_io_mod_mt_mod_header_id; // @[controller.scala 29:25]
  wire [5:0] proc_5_io_mod_mt_mod_key_off; // @[controller.scala 29:25]
  wire [5:0] proc_5_io_mod_mt_mod_key_len; // @[controller.scala 29:25]
  wire [5:0] proc_5_io_mod_mt_mod_val_len; // @[controller.scala 29:25]
  wire  proc_5_io_mod_ex_mod_start; // @[controller.scala 29:25]
  wire [63:0] proc_5_io_mod_ex_mod_ops_0; // @[controller.scala 29:25]
  wire [63:0] proc_5_io_mod_ex_mod_ops_1; // @[controller.scala 29:25]
  wire [63:0] proc_5_io_mod_ex_mod_ops_2; // @[controller.scala 29:25]
  wire [63:0] proc_5_io_mod_ex_mod_ops_3; // @[controller.scala 29:25]
  wire [63:0] proc_5_io_mod_ex_mod_ops_4; // @[controller.scala 29:25]
  wire [63:0] proc_5_io_mod_ex_mod_ops_5; // @[controller.scala 29:25]
  wire [63:0] proc_5_io_mod_ex_mod_ops_6; // @[controller.scala 29:25]
  wire [63:0] proc_5_io_mod_ex_mod_ops_7; // @[controller.scala 29:25]
  wire [63:0] proc_5_io_mod_ex_mod_ops_8; // @[controller.scala 29:25]
  wire [63:0] proc_5_io_mod_ex_mod_ops_9; // @[controller.scala 29:25]
  wire [63:0] proc_5_io_mod_ex_mod_ops_10; // @[controller.scala 29:25]
  wire [63:0] proc_5_io_mod_ex_mod_ops_11; // @[controller.scala 29:25]
  wire [63:0] proc_5_io_mod_ex_mod_ops_12; // @[controller.scala 29:25]
  wire [63:0] proc_5_io_mod_ex_mod_ops_13; // @[controller.scala 29:25]
  wire [63:0] proc_5_io_mod_ex_mod_ops_14; // @[controller.scala 29:25]
  wire [63:0] proc_5_io_mod_ex_mod_ops_15; // @[controller.scala 29:25]
  wire  proc_5_io_next_en; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_next_header_0; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_next_header_1; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_next_header_2; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_next_header_3; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_next_header_4; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_next_header_5; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_next_header_6; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_next_header_7; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_next_header_8; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_next_header_9; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_next_header_10; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_next_header_11; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_next_header_12; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_next_header_13; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_next_header_14; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_next_header_15; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_next_header_16; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_next_header_17; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_next_header_18; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_next_header_19; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_next_header_20; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_next_header_21; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_next_header_22; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_next_header_23; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_next_header_24; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_next_header_25; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_next_header_26; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_next_header_27; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_next_header_28; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_next_header_29; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_next_header_30; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_next_header_31; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_next_header_32; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_next_header_33; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_next_header_34; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_next_header_35; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_next_header_36; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_next_header_37; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_next_header_38; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_next_header_39; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_next_header_40; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_next_header_41; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_next_header_42; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_next_header_43; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_next_header_44; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_next_header_45; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_next_header_46; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_next_header_47; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_next_header_48; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_next_header_49; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_next_header_50; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_next_header_51; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_next_header_52; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_next_header_53; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_next_header_54; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_next_header_55; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_next_header_56; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_next_header_57; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_next_header_58; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_next_header_59; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_next_header_60; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_next_header_61; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_next_header_62; // @[controller.scala 29:25]
  wire [7:0] proc_5_io_next_header_63; // @[controller.scala 29:25]
  wire [2:0] proc_5_io_next_proc; // @[controller.scala 29:25]
  wire  proc_6_clock; // @[controller.scala 29:25]
  wire  proc_6_reset; // @[controller.scala 29:25]
  wire  proc_6_io_update; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_packet_header_0; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_packet_header_1; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_packet_header_2; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_packet_header_3; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_packet_header_4; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_packet_header_5; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_packet_header_6; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_packet_header_7; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_packet_header_8; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_packet_header_9; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_packet_header_10; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_packet_header_11; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_packet_header_12; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_packet_header_13; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_packet_header_14; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_packet_header_15; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_packet_header_16; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_packet_header_17; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_packet_header_18; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_packet_header_19; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_packet_header_20; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_packet_header_21; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_packet_header_22; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_packet_header_23; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_packet_header_24; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_packet_header_25; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_packet_header_26; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_packet_header_27; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_packet_header_28; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_packet_header_29; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_packet_header_30; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_packet_header_31; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_packet_header_32; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_packet_header_33; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_packet_header_34; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_packet_header_35; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_packet_header_36; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_packet_header_37; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_packet_header_38; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_packet_header_39; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_packet_header_40; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_packet_header_41; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_packet_header_42; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_packet_header_43; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_packet_header_44; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_packet_header_45; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_packet_header_46; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_packet_header_47; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_packet_header_48; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_packet_header_49; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_packet_header_50; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_packet_header_51; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_packet_header_52; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_packet_header_53; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_packet_header_54; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_packet_header_55; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_packet_header_56; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_packet_header_57; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_packet_header_58; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_packet_header_59; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_packet_header_60; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_packet_header_61; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_packet_header_62; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_packet_header_63; // @[controller.scala 29:25]
  wire  proc_6_io_end; // @[controller.scala 29:25]
  wire [31:0] proc_6_io_mem_addr; // @[controller.scala 29:25]
  wire [31:0] proc_6_io_mem_rdata; // @[controller.scala 29:25]
  wire  proc_6_io_ready; // @[controller.scala 29:25]
  wire  proc_6_io_mod_start; // @[controller.scala 29:25]
  wire [31:0] proc_6_io_mod_hit_action_addr; // @[controller.scala 29:25]
  wire [31:0] proc_6_io_mod_miss_action_addr; // @[controller.scala 29:25]
  wire  proc_6_io_mod_ps_mod_start; // @[controller.scala 29:25]
  wire  proc_6_io_mod_ps_mod_header_id; // @[controller.scala 29:25]
  wire [31:0] proc_6_io_mod_ps_mod_header_length; // @[controller.scala 29:25]
  wire [31:0] proc_6_io_mod_ps_mod_next_tag_start; // @[controller.scala 29:25]
  wire [31:0] proc_6_io_mod_ps_mod_next_table_0; // @[controller.scala 29:25]
  wire [31:0] proc_6_io_mod_ps_mod_next_table_1; // @[controller.scala 29:25]
  wire  proc_6_io_mod_mt_mod_start; // @[controller.scala 29:25]
  wire [3:0] proc_6_io_mod_mt_mod_header_id; // @[controller.scala 29:25]
  wire [5:0] proc_6_io_mod_mt_mod_key_off; // @[controller.scala 29:25]
  wire [5:0] proc_6_io_mod_mt_mod_key_len; // @[controller.scala 29:25]
  wire [5:0] proc_6_io_mod_mt_mod_val_len; // @[controller.scala 29:25]
  wire  proc_6_io_mod_ex_mod_start; // @[controller.scala 29:25]
  wire [63:0] proc_6_io_mod_ex_mod_ops_0; // @[controller.scala 29:25]
  wire [63:0] proc_6_io_mod_ex_mod_ops_1; // @[controller.scala 29:25]
  wire [63:0] proc_6_io_mod_ex_mod_ops_2; // @[controller.scala 29:25]
  wire [63:0] proc_6_io_mod_ex_mod_ops_3; // @[controller.scala 29:25]
  wire [63:0] proc_6_io_mod_ex_mod_ops_4; // @[controller.scala 29:25]
  wire [63:0] proc_6_io_mod_ex_mod_ops_5; // @[controller.scala 29:25]
  wire [63:0] proc_6_io_mod_ex_mod_ops_6; // @[controller.scala 29:25]
  wire [63:0] proc_6_io_mod_ex_mod_ops_7; // @[controller.scala 29:25]
  wire [63:0] proc_6_io_mod_ex_mod_ops_8; // @[controller.scala 29:25]
  wire [63:0] proc_6_io_mod_ex_mod_ops_9; // @[controller.scala 29:25]
  wire [63:0] proc_6_io_mod_ex_mod_ops_10; // @[controller.scala 29:25]
  wire [63:0] proc_6_io_mod_ex_mod_ops_11; // @[controller.scala 29:25]
  wire [63:0] proc_6_io_mod_ex_mod_ops_12; // @[controller.scala 29:25]
  wire [63:0] proc_6_io_mod_ex_mod_ops_13; // @[controller.scala 29:25]
  wire [63:0] proc_6_io_mod_ex_mod_ops_14; // @[controller.scala 29:25]
  wire [63:0] proc_6_io_mod_ex_mod_ops_15; // @[controller.scala 29:25]
  wire  proc_6_io_next_en; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_next_header_0; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_next_header_1; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_next_header_2; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_next_header_3; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_next_header_4; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_next_header_5; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_next_header_6; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_next_header_7; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_next_header_8; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_next_header_9; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_next_header_10; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_next_header_11; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_next_header_12; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_next_header_13; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_next_header_14; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_next_header_15; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_next_header_16; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_next_header_17; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_next_header_18; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_next_header_19; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_next_header_20; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_next_header_21; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_next_header_22; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_next_header_23; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_next_header_24; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_next_header_25; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_next_header_26; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_next_header_27; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_next_header_28; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_next_header_29; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_next_header_30; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_next_header_31; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_next_header_32; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_next_header_33; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_next_header_34; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_next_header_35; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_next_header_36; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_next_header_37; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_next_header_38; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_next_header_39; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_next_header_40; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_next_header_41; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_next_header_42; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_next_header_43; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_next_header_44; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_next_header_45; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_next_header_46; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_next_header_47; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_next_header_48; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_next_header_49; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_next_header_50; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_next_header_51; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_next_header_52; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_next_header_53; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_next_header_54; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_next_header_55; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_next_header_56; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_next_header_57; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_next_header_58; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_next_header_59; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_next_header_60; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_next_header_61; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_next_header_62; // @[controller.scala 29:25]
  wire [7:0] proc_6_io_next_header_63; // @[controller.scala 29:25]
  wire [2:0] proc_6_io_next_proc; // @[controller.scala 29:25]
  wire  proc_7_clock; // @[controller.scala 29:25]
  wire  proc_7_reset; // @[controller.scala 29:25]
  wire  proc_7_io_update; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_packet_header_0; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_packet_header_1; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_packet_header_2; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_packet_header_3; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_packet_header_4; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_packet_header_5; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_packet_header_6; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_packet_header_7; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_packet_header_8; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_packet_header_9; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_packet_header_10; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_packet_header_11; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_packet_header_12; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_packet_header_13; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_packet_header_14; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_packet_header_15; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_packet_header_16; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_packet_header_17; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_packet_header_18; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_packet_header_19; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_packet_header_20; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_packet_header_21; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_packet_header_22; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_packet_header_23; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_packet_header_24; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_packet_header_25; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_packet_header_26; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_packet_header_27; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_packet_header_28; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_packet_header_29; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_packet_header_30; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_packet_header_31; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_packet_header_32; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_packet_header_33; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_packet_header_34; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_packet_header_35; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_packet_header_36; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_packet_header_37; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_packet_header_38; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_packet_header_39; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_packet_header_40; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_packet_header_41; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_packet_header_42; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_packet_header_43; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_packet_header_44; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_packet_header_45; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_packet_header_46; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_packet_header_47; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_packet_header_48; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_packet_header_49; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_packet_header_50; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_packet_header_51; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_packet_header_52; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_packet_header_53; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_packet_header_54; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_packet_header_55; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_packet_header_56; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_packet_header_57; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_packet_header_58; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_packet_header_59; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_packet_header_60; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_packet_header_61; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_packet_header_62; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_packet_header_63; // @[controller.scala 29:25]
  wire  proc_7_io_end; // @[controller.scala 29:25]
  wire [31:0] proc_7_io_mem_addr; // @[controller.scala 29:25]
  wire [31:0] proc_7_io_mem_rdata; // @[controller.scala 29:25]
  wire  proc_7_io_ready; // @[controller.scala 29:25]
  wire  proc_7_io_mod_start; // @[controller.scala 29:25]
  wire [31:0] proc_7_io_mod_hit_action_addr; // @[controller.scala 29:25]
  wire [31:0] proc_7_io_mod_miss_action_addr; // @[controller.scala 29:25]
  wire  proc_7_io_mod_ps_mod_start; // @[controller.scala 29:25]
  wire  proc_7_io_mod_ps_mod_header_id; // @[controller.scala 29:25]
  wire [31:0] proc_7_io_mod_ps_mod_header_length; // @[controller.scala 29:25]
  wire [31:0] proc_7_io_mod_ps_mod_next_tag_start; // @[controller.scala 29:25]
  wire [31:0] proc_7_io_mod_ps_mod_next_table_0; // @[controller.scala 29:25]
  wire [31:0] proc_7_io_mod_ps_mod_next_table_1; // @[controller.scala 29:25]
  wire  proc_7_io_mod_mt_mod_start; // @[controller.scala 29:25]
  wire [3:0] proc_7_io_mod_mt_mod_header_id; // @[controller.scala 29:25]
  wire [5:0] proc_7_io_mod_mt_mod_key_off; // @[controller.scala 29:25]
  wire [5:0] proc_7_io_mod_mt_mod_key_len; // @[controller.scala 29:25]
  wire [5:0] proc_7_io_mod_mt_mod_val_len; // @[controller.scala 29:25]
  wire  proc_7_io_mod_ex_mod_start; // @[controller.scala 29:25]
  wire [63:0] proc_7_io_mod_ex_mod_ops_0; // @[controller.scala 29:25]
  wire [63:0] proc_7_io_mod_ex_mod_ops_1; // @[controller.scala 29:25]
  wire [63:0] proc_7_io_mod_ex_mod_ops_2; // @[controller.scala 29:25]
  wire [63:0] proc_7_io_mod_ex_mod_ops_3; // @[controller.scala 29:25]
  wire [63:0] proc_7_io_mod_ex_mod_ops_4; // @[controller.scala 29:25]
  wire [63:0] proc_7_io_mod_ex_mod_ops_5; // @[controller.scala 29:25]
  wire [63:0] proc_7_io_mod_ex_mod_ops_6; // @[controller.scala 29:25]
  wire [63:0] proc_7_io_mod_ex_mod_ops_7; // @[controller.scala 29:25]
  wire [63:0] proc_7_io_mod_ex_mod_ops_8; // @[controller.scala 29:25]
  wire [63:0] proc_7_io_mod_ex_mod_ops_9; // @[controller.scala 29:25]
  wire [63:0] proc_7_io_mod_ex_mod_ops_10; // @[controller.scala 29:25]
  wire [63:0] proc_7_io_mod_ex_mod_ops_11; // @[controller.scala 29:25]
  wire [63:0] proc_7_io_mod_ex_mod_ops_12; // @[controller.scala 29:25]
  wire [63:0] proc_7_io_mod_ex_mod_ops_13; // @[controller.scala 29:25]
  wire [63:0] proc_7_io_mod_ex_mod_ops_14; // @[controller.scala 29:25]
  wire [63:0] proc_7_io_mod_ex_mod_ops_15; // @[controller.scala 29:25]
  wire  proc_7_io_next_en; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_next_header_0; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_next_header_1; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_next_header_2; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_next_header_3; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_next_header_4; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_next_header_5; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_next_header_6; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_next_header_7; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_next_header_8; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_next_header_9; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_next_header_10; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_next_header_11; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_next_header_12; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_next_header_13; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_next_header_14; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_next_header_15; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_next_header_16; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_next_header_17; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_next_header_18; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_next_header_19; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_next_header_20; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_next_header_21; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_next_header_22; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_next_header_23; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_next_header_24; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_next_header_25; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_next_header_26; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_next_header_27; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_next_header_28; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_next_header_29; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_next_header_30; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_next_header_31; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_next_header_32; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_next_header_33; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_next_header_34; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_next_header_35; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_next_header_36; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_next_header_37; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_next_header_38; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_next_header_39; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_next_header_40; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_next_header_41; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_next_header_42; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_next_header_43; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_next_header_44; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_next_header_45; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_next_header_46; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_next_header_47; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_next_header_48; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_next_header_49; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_next_header_50; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_next_header_51; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_next_header_52; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_next_header_53; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_next_header_54; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_next_header_55; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_next_header_56; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_next_header_57; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_next_header_58; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_next_header_59; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_next_header_60; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_next_header_61; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_next_header_62; // @[controller.scala 29:25]
  wire [7:0] proc_7_io_next_header_63; // @[controller.scala 29:25]
  wire [2:0] proc_7_io_next_proc; // @[controller.scala 29:25]
  wire  next_table_exe__0 = proc_0_io_ready & proc_0_io_next_en & proc_0_io_next_proc == 3'h0; // @[controller.scala 79:62]
  wire  next_table_exe__1 = proc_1_io_ready & proc_1_io_next_en & proc_1_io_next_proc == 3'h0; // @[controller.scala 79:62]
  wire  next_table_exe__2 = proc_2_io_ready & proc_2_io_next_en & proc_2_io_next_proc == 3'h0; // @[controller.scala 79:62]
  wire  next_table_exe__3 = proc_3_io_ready & proc_3_io_next_en & proc_3_io_next_proc == 3'h0; // @[controller.scala 79:62]
  wire  next_table_exe__4 = proc_4_io_ready & proc_4_io_next_en & proc_4_io_next_proc == 3'h0; // @[controller.scala 79:62]
  wire  next_table_exe__5 = proc_5_io_ready & proc_5_io_next_en & proc_5_io_next_proc == 3'h0; // @[controller.scala 79:62]
  wire  next_table_exe__6 = proc_6_io_ready & proc_6_io_next_en & proc_6_io_next_proc == 3'h0; // @[controller.scala 79:62]
  wire  next_table_exe__7 = proc_7_io_ready & proc_7_io_next_en & proc_7_io_next_proc == 3'h0; // @[controller.scala 79:62]
  wire [3:0] next_table_lo = {next_table_exe__3,next_table_exe__2,next_table_exe__1,next_table_exe__0}; // @[Cat.scala 30:58]
  wire [3:0] next_table_hi = {next_table_exe__7,next_table_exe__6,next_table_exe__5,next_table_exe__4}; // @[Cat.scala 30:58]
  wire  next_table_exe_1_0 = proc_0_io_ready & proc_0_io_next_en & proc_0_io_next_proc == 3'h1; // @[controller.scala 79:62]
  wire  next_table_exe_1_1 = proc_1_io_ready & proc_1_io_next_en & proc_1_io_next_proc == 3'h1; // @[controller.scala 79:62]
  wire  next_table_exe_1_2 = proc_2_io_ready & proc_2_io_next_en & proc_2_io_next_proc == 3'h1; // @[controller.scala 79:62]
  wire  next_table_exe_1_3 = proc_3_io_ready & proc_3_io_next_en & proc_3_io_next_proc == 3'h1; // @[controller.scala 79:62]
  wire  next_table_exe_1_4 = proc_4_io_ready & proc_4_io_next_en & proc_4_io_next_proc == 3'h1; // @[controller.scala 79:62]
  wire  next_table_exe_1_5 = proc_5_io_ready & proc_5_io_next_en & proc_5_io_next_proc == 3'h1; // @[controller.scala 79:62]
  wire  next_table_exe_1_6 = proc_6_io_ready & proc_6_io_next_en & proc_6_io_next_proc == 3'h1; // @[controller.scala 79:62]
  wire  next_table_exe_1_7 = proc_7_io_ready & proc_7_io_next_en & proc_7_io_next_proc == 3'h1; // @[controller.scala 79:62]
  wire [3:0] next_table_lo_1 = {next_table_exe_1_3,next_table_exe_1_2,next_table_exe_1_1,next_table_exe_1_0}; // @[Cat.scala 30:58]
  wire [3:0] next_table_hi_1 = {next_table_exe_1_7,next_table_exe_1_6,next_table_exe_1_5,next_table_exe_1_4}; // @[Cat.scala 30:58]
  wire  next_table_exe_2_0 = proc_0_io_ready & proc_0_io_next_en & proc_0_io_next_proc == 3'h2; // @[controller.scala 79:62]
  wire  next_table_exe_2_1 = proc_1_io_ready & proc_1_io_next_en & proc_1_io_next_proc == 3'h2; // @[controller.scala 79:62]
  wire  next_table_exe_2_2 = proc_2_io_ready & proc_2_io_next_en & proc_2_io_next_proc == 3'h2; // @[controller.scala 79:62]
  wire  next_table_exe_2_3 = proc_3_io_ready & proc_3_io_next_en & proc_3_io_next_proc == 3'h2; // @[controller.scala 79:62]
  wire  next_table_exe_2_4 = proc_4_io_ready & proc_4_io_next_en & proc_4_io_next_proc == 3'h2; // @[controller.scala 79:62]
  wire  next_table_exe_2_5 = proc_5_io_ready & proc_5_io_next_en & proc_5_io_next_proc == 3'h2; // @[controller.scala 79:62]
  wire  next_table_exe_2_6 = proc_6_io_ready & proc_6_io_next_en & proc_6_io_next_proc == 3'h2; // @[controller.scala 79:62]
  wire  next_table_exe_2_7 = proc_7_io_ready & proc_7_io_next_en & proc_7_io_next_proc == 3'h2; // @[controller.scala 79:62]
  wire [3:0] next_table_lo_2 = {next_table_exe_2_3,next_table_exe_2_2,next_table_exe_2_1,next_table_exe_2_0}; // @[Cat.scala 30:58]
  wire [3:0] next_table_hi_2 = {next_table_exe_2_7,next_table_exe_2_6,next_table_exe_2_5,next_table_exe_2_4}; // @[Cat.scala 30:58]
  wire  next_table_exe_3_0 = proc_0_io_ready & proc_0_io_next_en & proc_0_io_next_proc == 3'h3; // @[controller.scala 79:62]
  wire  next_table_exe_3_1 = proc_1_io_ready & proc_1_io_next_en & proc_1_io_next_proc == 3'h3; // @[controller.scala 79:62]
  wire  next_table_exe_3_2 = proc_2_io_ready & proc_2_io_next_en & proc_2_io_next_proc == 3'h3; // @[controller.scala 79:62]
  wire  next_table_exe_3_3 = proc_3_io_ready & proc_3_io_next_en & proc_3_io_next_proc == 3'h3; // @[controller.scala 79:62]
  wire  next_table_exe_3_4 = proc_4_io_ready & proc_4_io_next_en & proc_4_io_next_proc == 3'h3; // @[controller.scala 79:62]
  wire  next_table_exe_3_5 = proc_5_io_ready & proc_5_io_next_en & proc_5_io_next_proc == 3'h3; // @[controller.scala 79:62]
  wire  next_table_exe_3_6 = proc_6_io_ready & proc_6_io_next_en & proc_6_io_next_proc == 3'h3; // @[controller.scala 79:62]
  wire  next_table_exe_3_7 = proc_7_io_ready & proc_7_io_next_en & proc_7_io_next_proc == 3'h3; // @[controller.scala 79:62]
  wire [3:0] next_table_lo_3 = {next_table_exe_3_3,next_table_exe_3_2,next_table_exe_3_1,next_table_exe_3_0}; // @[Cat.scala 30:58]
  wire [3:0] next_table_hi_3 = {next_table_exe_3_7,next_table_exe_3_6,next_table_exe_3_5,next_table_exe_3_4}; // @[Cat.scala 30:58]
  wire  next_table_exe_4_0 = proc_0_io_ready & proc_0_io_next_en & proc_0_io_next_proc == 3'h4; // @[controller.scala 79:62]
  wire  next_table_exe_4_1 = proc_1_io_ready & proc_1_io_next_en & proc_1_io_next_proc == 3'h4; // @[controller.scala 79:62]
  wire  next_table_exe_4_2 = proc_2_io_ready & proc_2_io_next_en & proc_2_io_next_proc == 3'h4; // @[controller.scala 79:62]
  wire  next_table_exe_4_3 = proc_3_io_ready & proc_3_io_next_en & proc_3_io_next_proc == 3'h4; // @[controller.scala 79:62]
  wire  next_table_exe_4_4 = proc_4_io_ready & proc_4_io_next_en & proc_4_io_next_proc == 3'h4; // @[controller.scala 79:62]
  wire  next_table_exe_4_5 = proc_5_io_ready & proc_5_io_next_en & proc_5_io_next_proc == 3'h4; // @[controller.scala 79:62]
  wire  next_table_exe_4_6 = proc_6_io_ready & proc_6_io_next_en & proc_6_io_next_proc == 3'h4; // @[controller.scala 79:62]
  wire  next_table_exe_4_7 = proc_7_io_ready & proc_7_io_next_en & proc_7_io_next_proc == 3'h4; // @[controller.scala 79:62]
  wire [3:0] next_table_lo_4 = {next_table_exe_4_3,next_table_exe_4_2,next_table_exe_4_1,next_table_exe_4_0}; // @[Cat.scala 30:58]
  wire [3:0] next_table_hi_4 = {next_table_exe_4_7,next_table_exe_4_6,next_table_exe_4_5,next_table_exe_4_4}; // @[Cat.scala 30:58]
  wire  next_table_exe_5_0 = proc_0_io_ready & proc_0_io_next_en & proc_0_io_next_proc == 3'h5; // @[controller.scala 79:62]
  wire  next_table_exe_5_1 = proc_1_io_ready & proc_1_io_next_en & proc_1_io_next_proc == 3'h5; // @[controller.scala 79:62]
  wire  next_table_exe_5_2 = proc_2_io_ready & proc_2_io_next_en & proc_2_io_next_proc == 3'h5; // @[controller.scala 79:62]
  wire  next_table_exe_5_3 = proc_3_io_ready & proc_3_io_next_en & proc_3_io_next_proc == 3'h5; // @[controller.scala 79:62]
  wire  next_table_exe_5_4 = proc_4_io_ready & proc_4_io_next_en & proc_4_io_next_proc == 3'h5; // @[controller.scala 79:62]
  wire  next_table_exe_5_5 = proc_5_io_ready & proc_5_io_next_en & proc_5_io_next_proc == 3'h5; // @[controller.scala 79:62]
  wire  next_table_exe_5_6 = proc_6_io_ready & proc_6_io_next_en & proc_6_io_next_proc == 3'h5; // @[controller.scala 79:62]
  wire  next_table_exe_5_7 = proc_7_io_ready & proc_7_io_next_en & proc_7_io_next_proc == 3'h5; // @[controller.scala 79:62]
  wire [3:0] next_table_lo_5 = {next_table_exe_5_3,next_table_exe_5_2,next_table_exe_5_1,next_table_exe_5_0}; // @[Cat.scala 30:58]
  wire [3:0] next_table_hi_5 = {next_table_exe_5_7,next_table_exe_5_6,next_table_exe_5_5,next_table_exe_5_4}; // @[Cat.scala 30:58]
  wire  next_table_exe_6_0 = proc_0_io_ready & proc_0_io_next_en & proc_0_io_next_proc == 3'h6; // @[controller.scala 79:62]
  wire  next_table_exe_6_1 = proc_1_io_ready & proc_1_io_next_en & proc_1_io_next_proc == 3'h6; // @[controller.scala 79:62]
  wire  next_table_exe_6_2 = proc_2_io_ready & proc_2_io_next_en & proc_2_io_next_proc == 3'h6; // @[controller.scala 79:62]
  wire  next_table_exe_6_3 = proc_3_io_ready & proc_3_io_next_en & proc_3_io_next_proc == 3'h6; // @[controller.scala 79:62]
  wire  next_table_exe_6_4 = proc_4_io_ready & proc_4_io_next_en & proc_4_io_next_proc == 3'h6; // @[controller.scala 79:62]
  wire  next_table_exe_6_5 = proc_5_io_ready & proc_5_io_next_en & proc_5_io_next_proc == 3'h6; // @[controller.scala 79:62]
  wire  next_table_exe_6_6 = proc_6_io_ready & proc_6_io_next_en & proc_6_io_next_proc == 3'h6; // @[controller.scala 79:62]
  wire  next_table_exe_6_7 = proc_7_io_ready & proc_7_io_next_en & proc_7_io_next_proc == 3'h6; // @[controller.scala 79:62]
  wire [3:0] next_table_lo_6 = {next_table_exe_6_3,next_table_exe_6_2,next_table_exe_6_1,next_table_exe_6_0}; // @[Cat.scala 30:58]
  wire [3:0] next_table_hi_6 = {next_table_exe_6_7,next_table_exe_6_6,next_table_exe_6_5,next_table_exe_6_4}; // @[Cat.scala 30:58]
  wire  next_table_exe_7_0 = proc_0_io_ready & proc_0_io_next_en & proc_0_io_next_proc == 3'h7; // @[controller.scala 79:62]
  wire  next_table_exe_7_1 = proc_1_io_ready & proc_1_io_next_en & proc_1_io_next_proc == 3'h7; // @[controller.scala 79:62]
  wire  next_table_exe_7_2 = proc_2_io_ready & proc_2_io_next_en & proc_2_io_next_proc == 3'h7; // @[controller.scala 79:62]
  wire  next_table_exe_7_3 = proc_3_io_ready & proc_3_io_next_en & proc_3_io_next_proc == 3'h7; // @[controller.scala 79:62]
  wire  next_table_exe_7_4 = proc_4_io_ready & proc_4_io_next_en & proc_4_io_next_proc == 3'h7; // @[controller.scala 79:62]
  wire  next_table_exe_7_5 = proc_5_io_ready & proc_5_io_next_en & proc_5_io_next_proc == 3'h7; // @[controller.scala 79:62]
  wire  next_table_exe_7_6 = proc_6_io_ready & proc_6_io_next_en & proc_6_io_next_proc == 3'h7; // @[controller.scala 79:62]
  wire  next_table_exe_7_7 = proc_7_io_ready & proc_7_io_next_en & proc_7_io_next_proc == 3'h7; // @[controller.scala 79:62]
  wire [3:0] next_table_lo_7 = {next_table_exe_7_3,next_table_exe_7_2,next_table_exe_7_1,next_table_exe_7_0}; // @[Cat.scala 30:58]
  wire [3:0] next_table_hi_7 = {next_table_exe_7_7,next_table_exe_7_6,next_table_exe_7_5,next_table_exe_7_4}; // @[Cat.scala 30:58]
  wire [7:0] _GEN_256 = 3'h0 == encoders_0_io_output ? proc_0_io_next_header_0 : io_packet_header_0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 38:34]
  wire [7:0] _GEN_257 = 3'h0 == encoders_0_io_output ? proc_0_io_next_header_1 : io_packet_header_1; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 38:34]
  wire [7:0] _GEN_258 = 3'h0 == encoders_0_io_output ? proc_0_io_next_header_2 : io_packet_header_2; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 38:34]
  wire [7:0] _GEN_259 = 3'h0 == encoders_0_io_output ? proc_0_io_next_header_3 : io_packet_header_3; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 38:34]
  wire [7:0] _GEN_260 = 3'h0 == encoders_0_io_output ? proc_0_io_next_header_4 : io_packet_header_4; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 38:34]
  wire [7:0] _GEN_261 = 3'h0 == encoders_0_io_output ? proc_0_io_next_header_5 : io_packet_header_5; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 38:34]
  wire [7:0] _GEN_262 = 3'h0 == encoders_0_io_output ? proc_0_io_next_header_6 : io_packet_header_6; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 38:34]
  wire [7:0] _GEN_263 = 3'h0 == encoders_0_io_output ? proc_0_io_next_header_7 : io_packet_header_7; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 38:34]
  wire [7:0] _GEN_264 = 3'h0 == encoders_0_io_output ? proc_0_io_next_header_8 : io_packet_header_8; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 38:34]
  wire [7:0] _GEN_265 = 3'h0 == encoders_0_io_output ? proc_0_io_next_header_9 : io_packet_header_9; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 38:34]
  wire [7:0] _GEN_266 = 3'h0 == encoders_0_io_output ? proc_0_io_next_header_10 : io_packet_header_10; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 38:34]
  wire [7:0] _GEN_267 = 3'h0 == encoders_0_io_output ? proc_0_io_next_header_11 : io_packet_header_11; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 38:34]
  wire [7:0] _GEN_268 = 3'h0 == encoders_0_io_output ? proc_0_io_next_header_12 : io_packet_header_12; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 38:34]
  wire [7:0] _GEN_269 = 3'h0 == encoders_0_io_output ? proc_0_io_next_header_13 : io_packet_header_13; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 38:34]
  wire [7:0] _GEN_270 = 3'h0 == encoders_0_io_output ? proc_0_io_next_header_14 : io_packet_header_14; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 38:34]
  wire [7:0] _GEN_271 = 3'h0 == encoders_0_io_output ? proc_0_io_next_header_15 : io_packet_header_15; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 38:34]
  wire [7:0] _GEN_272 = 3'h0 == encoders_0_io_output ? proc_0_io_next_header_16 : io_packet_header_16; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 38:34]
  wire [7:0] _GEN_273 = 3'h0 == encoders_0_io_output ? proc_0_io_next_header_17 : io_packet_header_17; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 38:34]
  wire [7:0] _GEN_274 = 3'h0 == encoders_0_io_output ? proc_0_io_next_header_18 : io_packet_header_18; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 38:34]
  wire [7:0] _GEN_275 = 3'h0 == encoders_0_io_output ? proc_0_io_next_header_19 : io_packet_header_19; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 38:34]
  wire [7:0] _GEN_276 = 3'h0 == encoders_0_io_output ? proc_0_io_next_header_20 : io_packet_header_20; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 38:34]
  wire [7:0] _GEN_277 = 3'h0 == encoders_0_io_output ? proc_0_io_next_header_21 : io_packet_header_21; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 38:34]
  wire [7:0] _GEN_278 = 3'h0 == encoders_0_io_output ? proc_0_io_next_header_22 : io_packet_header_22; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 38:34]
  wire [7:0] _GEN_279 = 3'h0 == encoders_0_io_output ? proc_0_io_next_header_23 : io_packet_header_23; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 38:34]
  wire [7:0] _GEN_280 = 3'h0 == encoders_0_io_output ? proc_0_io_next_header_24 : io_packet_header_24; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 38:34]
  wire [7:0] _GEN_281 = 3'h0 == encoders_0_io_output ? proc_0_io_next_header_25 : io_packet_header_25; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 38:34]
  wire [7:0] _GEN_282 = 3'h0 == encoders_0_io_output ? proc_0_io_next_header_26 : io_packet_header_26; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 38:34]
  wire [7:0] _GEN_283 = 3'h0 == encoders_0_io_output ? proc_0_io_next_header_27 : io_packet_header_27; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 38:34]
  wire [7:0] _GEN_284 = 3'h0 == encoders_0_io_output ? proc_0_io_next_header_28 : io_packet_header_28; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 38:34]
  wire [7:0] _GEN_285 = 3'h0 == encoders_0_io_output ? proc_0_io_next_header_29 : io_packet_header_29; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 38:34]
  wire [7:0] _GEN_286 = 3'h0 == encoders_0_io_output ? proc_0_io_next_header_30 : io_packet_header_30; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 38:34]
  wire [7:0] _GEN_287 = 3'h0 == encoders_0_io_output ? proc_0_io_next_header_31 : io_packet_header_31; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 38:34]
  wire [7:0] _GEN_288 = 3'h0 == encoders_0_io_output ? proc_0_io_next_header_32 : io_packet_header_32; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 38:34]
  wire [7:0] _GEN_289 = 3'h0 == encoders_0_io_output ? proc_0_io_next_header_33 : io_packet_header_33; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 38:34]
  wire [7:0] _GEN_290 = 3'h0 == encoders_0_io_output ? proc_0_io_next_header_34 : io_packet_header_34; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 38:34]
  wire [7:0] _GEN_291 = 3'h0 == encoders_0_io_output ? proc_0_io_next_header_35 : io_packet_header_35; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 38:34]
  wire [7:0] _GEN_292 = 3'h0 == encoders_0_io_output ? proc_0_io_next_header_36 : io_packet_header_36; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 38:34]
  wire [7:0] _GEN_293 = 3'h0 == encoders_0_io_output ? proc_0_io_next_header_37 : io_packet_header_37; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 38:34]
  wire [7:0] _GEN_294 = 3'h0 == encoders_0_io_output ? proc_0_io_next_header_38 : io_packet_header_38; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 38:34]
  wire [7:0] _GEN_295 = 3'h0 == encoders_0_io_output ? proc_0_io_next_header_39 : io_packet_header_39; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 38:34]
  wire [7:0] _GEN_296 = 3'h0 == encoders_0_io_output ? proc_0_io_next_header_40 : io_packet_header_40; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 38:34]
  wire [7:0] _GEN_297 = 3'h0 == encoders_0_io_output ? proc_0_io_next_header_41 : io_packet_header_41; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 38:34]
  wire [7:0] _GEN_298 = 3'h0 == encoders_0_io_output ? proc_0_io_next_header_42 : io_packet_header_42; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 38:34]
  wire [7:0] _GEN_299 = 3'h0 == encoders_0_io_output ? proc_0_io_next_header_43 : io_packet_header_43; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 38:34]
  wire [7:0] _GEN_300 = 3'h0 == encoders_0_io_output ? proc_0_io_next_header_44 : io_packet_header_44; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 38:34]
  wire [7:0] _GEN_301 = 3'h0 == encoders_0_io_output ? proc_0_io_next_header_45 : io_packet_header_45; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 38:34]
  wire [7:0] _GEN_302 = 3'h0 == encoders_0_io_output ? proc_0_io_next_header_46 : io_packet_header_46; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 38:34]
  wire [7:0] _GEN_303 = 3'h0 == encoders_0_io_output ? proc_0_io_next_header_47 : io_packet_header_47; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 38:34]
  wire [7:0] _GEN_304 = 3'h0 == encoders_0_io_output ? proc_0_io_next_header_48 : io_packet_header_48; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 38:34]
  wire [7:0] _GEN_305 = 3'h0 == encoders_0_io_output ? proc_0_io_next_header_49 : io_packet_header_49; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 38:34]
  wire [7:0] _GEN_306 = 3'h0 == encoders_0_io_output ? proc_0_io_next_header_50 : io_packet_header_50; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 38:34]
  wire [7:0] _GEN_307 = 3'h0 == encoders_0_io_output ? proc_0_io_next_header_51 : io_packet_header_51; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 38:34]
  wire [7:0] _GEN_308 = 3'h0 == encoders_0_io_output ? proc_0_io_next_header_52 : io_packet_header_52; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 38:34]
  wire [7:0] _GEN_309 = 3'h0 == encoders_0_io_output ? proc_0_io_next_header_53 : io_packet_header_53; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 38:34]
  wire [7:0] _GEN_310 = 3'h0 == encoders_0_io_output ? proc_0_io_next_header_54 : io_packet_header_54; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 38:34]
  wire [7:0] _GEN_311 = 3'h0 == encoders_0_io_output ? proc_0_io_next_header_55 : io_packet_header_55; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 38:34]
  wire [7:0] _GEN_312 = 3'h0 == encoders_0_io_output ? proc_0_io_next_header_56 : io_packet_header_56; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 38:34]
  wire [7:0] _GEN_313 = 3'h0 == encoders_0_io_output ? proc_0_io_next_header_57 : io_packet_header_57; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 38:34]
  wire [7:0] _GEN_314 = 3'h0 == encoders_0_io_output ? proc_0_io_next_header_58 : io_packet_header_58; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 38:34]
  wire [7:0] _GEN_315 = 3'h0 == encoders_0_io_output ? proc_0_io_next_header_59 : io_packet_header_59; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 38:34]
  wire [7:0] _GEN_316 = 3'h0 == encoders_0_io_output ? proc_0_io_next_header_60 : io_packet_header_60; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 38:34]
  wire [7:0] _GEN_317 = 3'h0 == encoders_0_io_output ? proc_0_io_next_header_61 : io_packet_header_61; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 38:34]
  wire [7:0] _GEN_318 = 3'h0 == encoders_0_io_output ? proc_0_io_next_header_62 : io_packet_header_62; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 38:34]
  wire [7:0] _GEN_319 = 3'h0 == encoders_0_io_output ? proc_0_io_next_header_63 : io_packet_header_63; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 38:34]
  wire [7:0] _GEN_320 = 3'h1 == encoders_0_io_output ? proc_1_io_next_header_0 : _GEN_256; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_321 = 3'h1 == encoders_0_io_output ? proc_1_io_next_header_1 : _GEN_257; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_322 = 3'h1 == encoders_0_io_output ? proc_1_io_next_header_2 : _GEN_258; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_323 = 3'h1 == encoders_0_io_output ? proc_1_io_next_header_3 : _GEN_259; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_324 = 3'h1 == encoders_0_io_output ? proc_1_io_next_header_4 : _GEN_260; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_325 = 3'h1 == encoders_0_io_output ? proc_1_io_next_header_5 : _GEN_261; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_326 = 3'h1 == encoders_0_io_output ? proc_1_io_next_header_6 : _GEN_262; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_327 = 3'h1 == encoders_0_io_output ? proc_1_io_next_header_7 : _GEN_263; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_328 = 3'h1 == encoders_0_io_output ? proc_1_io_next_header_8 : _GEN_264; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_329 = 3'h1 == encoders_0_io_output ? proc_1_io_next_header_9 : _GEN_265; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_330 = 3'h1 == encoders_0_io_output ? proc_1_io_next_header_10 : _GEN_266; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_331 = 3'h1 == encoders_0_io_output ? proc_1_io_next_header_11 : _GEN_267; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_332 = 3'h1 == encoders_0_io_output ? proc_1_io_next_header_12 : _GEN_268; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_333 = 3'h1 == encoders_0_io_output ? proc_1_io_next_header_13 : _GEN_269; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_334 = 3'h1 == encoders_0_io_output ? proc_1_io_next_header_14 : _GEN_270; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_335 = 3'h1 == encoders_0_io_output ? proc_1_io_next_header_15 : _GEN_271; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_336 = 3'h1 == encoders_0_io_output ? proc_1_io_next_header_16 : _GEN_272; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_337 = 3'h1 == encoders_0_io_output ? proc_1_io_next_header_17 : _GEN_273; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_338 = 3'h1 == encoders_0_io_output ? proc_1_io_next_header_18 : _GEN_274; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_339 = 3'h1 == encoders_0_io_output ? proc_1_io_next_header_19 : _GEN_275; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_340 = 3'h1 == encoders_0_io_output ? proc_1_io_next_header_20 : _GEN_276; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_341 = 3'h1 == encoders_0_io_output ? proc_1_io_next_header_21 : _GEN_277; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_342 = 3'h1 == encoders_0_io_output ? proc_1_io_next_header_22 : _GEN_278; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_343 = 3'h1 == encoders_0_io_output ? proc_1_io_next_header_23 : _GEN_279; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_344 = 3'h1 == encoders_0_io_output ? proc_1_io_next_header_24 : _GEN_280; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_345 = 3'h1 == encoders_0_io_output ? proc_1_io_next_header_25 : _GEN_281; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_346 = 3'h1 == encoders_0_io_output ? proc_1_io_next_header_26 : _GEN_282; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_347 = 3'h1 == encoders_0_io_output ? proc_1_io_next_header_27 : _GEN_283; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_348 = 3'h1 == encoders_0_io_output ? proc_1_io_next_header_28 : _GEN_284; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_349 = 3'h1 == encoders_0_io_output ? proc_1_io_next_header_29 : _GEN_285; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_350 = 3'h1 == encoders_0_io_output ? proc_1_io_next_header_30 : _GEN_286; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_351 = 3'h1 == encoders_0_io_output ? proc_1_io_next_header_31 : _GEN_287; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_352 = 3'h1 == encoders_0_io_output ? proc_1_io_next_header_32 : _GEN_288; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_353 = 3'h1 == encoders_0_io_output ? proc_1_io_next_header_33 : _GEN_289; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_354 = 3'h1 == encoders_0_io_output ? proc_1_io_next_header_34 : _GEN_290; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_355 = 3'h1 == encoders_0_io_output ? proc_1_io_next_header_35 : _GEN_291; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_356 = 3'h1 == encoders_0_io_output ? proc_1_io_next_header_36 : _GEN_292; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_357 = 3'h1 == encoders_0_io_output ? proc_1_io_next_header_37 : _GEN_293; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_358 = 3'h1 == encoders_0_io_output ? proc_1_io_next_header_38 : _GEN_294; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_359 = 3'h1 == encoders_0_io_output ? proc_1_io_next_header_39 : _GEN_295; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_360 = 3'h1 == encoders_0_io_output ? proc_1_io_next_header_40 : _GEN_296; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_361 = 3'h1 == encoders_0_io_output ? proc_1_io_next_header_41 : _GEN_297; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_362 = 3'h1 == encoders_0_io_output ? proc_1_io_next_header_42 : _GEN_298; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_363 = 3'h1 == encoders_0_io_output ? proc_1_io_next_header_43 : _GEN_299; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_364 = 3'h1 == encoders_0_io_output ? proc_1_io_next_header_44 : _GEN_300; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_365 = 3'h1 == encoders_0_io_output ? proc_1_io_next_header_45 : _GEN_301; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_366 = 3'h1 == encoders_0_io_output ? proc_1_io_next_header_46 : _GEN_302; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_367 = 3'h1 == encoders_0_io_output ? proc_1_io_next_header_47 : _GEN_303; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_368 = 3'h1 == encoders_0_io_output ? proc_1_io_next_header_48 : _GEN_304; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_369 = 3'h1 == encoders_0_io_output ? proc_1_io_next_header_49 : _GEN_305; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_370 = 3'h1 == encoders_0_io_output ? proc_1_io_next_header_50 : _GEN_306; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_371 = 3'h1 == encoders_0_io_output ? proc_1_io_next_header_51 : _GEN_307; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_372 = 3'h1 == encoders_0_io_output ? proc_1_io_next_header_52 : _GEN_308; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_373 = 3'h1 == encoders_0_io_output ? proc_1_io_next_header_53 : _GEN_309; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_374 = 3'h1 == encoders_0_io_output ? proc_1_io_next_header_54 : _GEN_310; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_375 = 3'h1 == encoders_0_io_output ? proc_1_io_next_header_55 : _GEN_311; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_376 = 3'h1 == encoders_0_io_output ? proc_1_io_next_header_56 : _GEN_312; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_377 = 3'h1 == encoders_0_io_output ? proc_1_io_next_header_57 : _GEN_313; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_378 = 3'h1 == encoders_0_io_output ? proc_1_io_next_header_58 : _GEN_314; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_379 = 3'h1 == encoders_0_io_output ? proc_1_io_next_header_59 : _GEN_315; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_380 = 3'h1 == encoders_0_io_output ? proc_1_io_next_header_60 : _GEN_316; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_381 = 3'h1 == encoders_0_io_output ? proc_1_io_next_header_61 : _GEN_317; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_382 = 3'h1 == encoders_0_io_output ? proc_1_io_next_header_62 : _GEN_318; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_383 = 3'h1 == encoders_0_io_output ? proc_1_io_next_header_63 : _GEN_319; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_384 = 3'h2 == encoders_0_io_output ? proc_2_io_next_header_0 : _GEN_320; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_385 = 3'h2 == encoders_0_io_output ? proc_2_io_next_header_1 : _GEN_321; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_386 = 3'h2 == encoders_0_io_output ? proc_2_io_next_header_2 : _GEN_322; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_387 = 3'h2 == encoders_0_io_output ? proc_2_io_next_header_3 : _GEN_323; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_388 = 3'h2 == encoders_0_io_output ? proc_2_io_next_header_4 : _GEN_324; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_389 = 3'h2 == encoders_0_io_output ? proc_2_io_next_header_5 : _GEN_325; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_390 = 3'h2 == encoders_0_io_output ? proc_2_io_next_header_6 : _GEN_326; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_391 = 3'h2 == encoders_0_io_output ? proc_2_io_next_header_7 : _GEN_327; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_392 = 3'h2 == encoders_0_io_output ? proc_2_io_next_header_8 : _GEN_328; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_393 = 3'h2 == encoders_0_io_output ? proc_2_io_next_header_9 : _GEN_329; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_394 = 3'h2 == encoders_0_io_output ? proc_2_io_next_header_10 : _GEN_330; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_395 = 3'h2 == encoders_0_io_output ? proc_2_io_next_header_11 : _GEN_331; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_396 = 3'h2 == encoders_0_io_output ? proc_2_io_next_header_12 : _GEN_332; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_397 = 3'h2 == encoders_0_io_output ? proc_2_io_next_header_13 : _GEN_333; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_398 = 3'h2 == encoders_0_io_output ? proc_2_io_next_header_14 : _GEN_334; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_399 = 3'h2 == encoders_0_io_output ? proc_2_io_next_header_15 : _GEN_335; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_400 = 3'h2 == encoders_0_io_output ? proc_2_io_next_header_16 : _GEN_336; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_401 = 3'h2 == encoders_0_io_output ? proc_2_io_next_header_17 : _GEN_337; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_402 = 3'h2 == encoders_0_io_output ? proc_2_io_next_header_18 : _GEN_338; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_403 = 3'h2 == encoders_0_io_output ? proc_2_io_next_header_19 : _GEN_339; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_404 = 3'h2 == encoders_0_io_output ? proc_2_io_next_header_20 : _GEN_340; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_405 = 3'h2 == encoders_0_io_output ? proc_2_io_next_header_21 : _GEN_341; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_406 = 3'h2 == encoders_0_io_output ? proc_2_io_next_header_22 : _GEN_342; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_407 = 3'h2 == encoders_0_io_output ? proc_2_io_next_header_23 : _GEN_343; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_408 = 3'h2 == encoders_0_io_output ? proc_2_io_next_header_24 : _GEN_344; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_409 = 3'h2 == encoders_0_io_output ? proc_2_io_next_header_25 : _GEN_345; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_410 = 3'h2 == encoders_0_io_output ? proc_2_io_next_header_26 : _GEN_346; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_411 = 3'h2 == encoders_0_io_output ? proc_2_io_next_header_27 : _GEN_347; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_412 = 3'h2 == encoders_0_io_output ? proc_2_io_next_header_28 : _GEN_348; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_413 = 3'h2 == encoders_0_io_output ? proc_2_io_next_header_29 : _GEN_349; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_414 = 3'h2 == encoders_0_io_output ? proc_2_io_next_header_30 : _GEN_350; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_415 = 3'h2 == encoders_0_io_output ? proc_2_io_next_header_31 : _GEN_351; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_416 = 3'h2 == encoders_0_io_output ? proc_2_io_next_header_32 : _GEN_352; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_417 = 3'h2 == encoders_0_io_output ? proc_2_io_next_header_33 : _GEN_353; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_418 = 3'h2 == encoders_0_io_output ? proc_2_io_next_header_34 : _GEN_354; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_419 = 3'h2 == encoders_0_io_output ? proc_2_io_next_header_35 : _GEN_355; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_420 = 3'h2 == encoders_0_io_output ? proc_2_io_next_header_36 : _GEN_356; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_421 = 3'h2 == encoders_0_io_output ? proc_2_io_next_header_37 : _GEN_357; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_422 = 3'h2 == encoders_0_io_output ? proc_2_io_next_header_38 : _GEN_358; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_423 = 3'h2 == encoders_0_io_output ? proc_2_io_next_header_39 : _GEN_359; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_424 = 3'h2 == encoders_0_io_output ? proc_2_io_next_header_40 : _GEN_360; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_425 = 3'h2 == encoders_0_io_output ? proc_2_io_next_header_41 : _GEN_361; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_426 = 3'h2 == encoders_0_io_output ? proc_2_io_next_header_42 : _GEN_362; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_427 = 3'h2 == encoders_0_io_output ? proc_2_io_next_header_43 : _GEN_363; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_428 = 3'h2 == encoders_0_io_output ? proc_2_io_next_header_44 : _GEN_364; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_429 = 3'h2 == encoders_0_io_output ? proc_2_io_next_header_45 : _GEN_365; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_430 = 3'h2 == encoders_0_io_output ? proc_2_io_next_header_46 : _GEN_366; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_431 = 3'h2 == encoders_0_io_output ? proc_2_io_next_header_47 : _GEN_367; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_432 = 3'h2 == encoders_0_io_output ? proc_2_io_next_header_48 : _GEN_368; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_433 = 3'h2 == encoders_0_io_output ? proc_2_io_next_header_49 : _GEN_369; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_434 = 3'h2 == encoders_0_io_output ? proc_2_io_next_header_50 : _GEN_370; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_435 = 3'h2 == encoders_0_io_output ? proc_2_io_next_header_51 : _GEN_371; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_436 = 3'h2 == encoders_0_io_output ? proc_2_io_next_header_52 : _GEN_372; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_437 = 3'h2 == encoders_0_io_output ? proc_2_io_next_header_53 : _GEN_373; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_438 = 3'h2 == encoders_0_io_output ? proc_2_io_next_header_54 : _GEN_374; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_439 = 3'h2 == encoders_0_io_output ? proc_2_io_next_header_55 : _GEN_375; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_440 = 3'h2 == encoders_0_io_output ? proc_2_io_next_header_56 : _GEN_376; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_441 = 3'h2 == encoders_0_io_output ? proc_2_io_next_header_57 : _GEN_377; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_442 = 3'h2 == encoders_0_io_output ? proc_2_io_next_header_58 : _GEN_378; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_443 = 3'h2 == encoders_0_io_output ? proc_2_io_next_header_59 : _GEN_379; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_444 = 3'h2 == encoders_0_io_output ? proc_2_io_next_header_60 : _GEN_380; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_445 = 3'h2 == encoders_0_io_output ? proc_2_io_next_header_61 : _GEN_381; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_446 = 3'h2 == encoders_0_io_output ? proc_2_io_next_header_62 : _GEN_382; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_447 = 3'h2 == encoders_0_io_output ? proc_2_io_next_header_63 : _GEN_383; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_448 = 3'h3 == encoders_0_io_output ? proc_3_io_next_header_0 : _GEN_384; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_449 = 3'h3 == encoders_0_io_output ? proc_3_io_next_header_1 : _GEN_385; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_450 = 3'h3 == encoders_0_io_output ? proc_3_io_next_header_2 : _GEN_386; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_451 = 3'h3 == encoders_0_io_output ? proc_3_io_next_header_3 : _GEN_387; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_452 = 3'h3 == encoders_0_io_output ? proc_3_io_next_header_4 : _GEN_388; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_453 = 3'h3 == encoders_0_io_output ? proc_3_io_next_header_5 : _GEN_389; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_454 = 3'h3 == encoders_0_io_output ? proc_3_io_next_header_6 : _GEN_390; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_455 = 3'h3 == encoders_0_io_output ? proc_3_io_next_header_7 : _GEN_391; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_456 = 3'h3 == encoders_0_io_output ? proc_3_io_next_header_8 : _GEN_392; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_457 = 3'h3 == encoders_0_io_output ? proc_3_io_next_header_9 : _GEN_393; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_458 = 3'h3 == encoders_0_io_output ? proc_3_io_next_header_10 : _GEN_394; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_459 = 3'h3 == encoders_0_io_output ? proc_3_io_next_header_11 : _GEN_395; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_460 = 3'h3 == encoders_0_io_output ? proc_3_io_next_header_12 : _GEN_396; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_461 = 3'h3 == encoders_0_io_output ? proc_3_io_next_header_13 : _GEN_397; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_462 = 3'h3 == encoders_0_io_output ? proc_3_io_next_header_14 : _GEN_398; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_463 = 3'h3 == encoders_0_io_output ? proc_3_io_next_header_15 : _GEN_399; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_464 = 3'h3 == encoders_0_io_output ? proc_3_io_next_header_16 : _GEN_400; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_465 = 3'h3 == encoders_0_io_output ? proc_3_io_next_header_17 : _GEN_401; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_466 = 3'h3 == encoders_0_io_output ? proc_3_io_next_header_18 : _GEN_402; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_467 = 3'h3 == encoders_0_io_output ? proc_3_io_next_header_19 : _GEN_403; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_468 = 3'h3 == encoders_0_io_output ? proc_3_io_next_header_20 : _GEN_404; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_469 = 3'h3 == encoders_0_io_output ? proc_3_io_next_header_21 : _GEN_405; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_470 = 3'h3 == encoders_0_io_output ? proc_3_io_next_header_22 : _GEN_406; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_471 = 3'h3 == encoders_0_io_output ? proc_3_io_next_header_23 : _GEN_407; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_472 = 3'h3 == encoders_0_io_output ? proc_3_io_next_header_24 : _GEN_408; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_473 = 3'h3 == encoders_0_io_output ? proc_3_io_next_header_25 : _GEN_409; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_474 = 3'h3 == encoders_0_io_output ? proc_3_io_next_header_26 : _GEN_410; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_475 = 3'h3 == encoders_0_io_output ? proc_3_io_next_header_27 : _GEN_411; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_476 = 3'h3 == encoders_0_io_output ? proc_3_io_next_header_28 : _GEN_412; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_477 = 3'h3 == encoders_0_io_output ? proc_3_io_next_header_29 : _GEN_413; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_478 = 3'h3 == encoders_0_io_output ? proc_3_io_next_header_30 : _GEN_414; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_479 = 3'h3 == encoders_0_io_output ? proc_3_io_next_header_31 : _GEN_415; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_480 = 3'h3 == encoders_0_io_output ? proc_3_io_next_header_32 : _GEN_416; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_481 = 3'h3 == encoders_0_io_output ? proc_3_io_next_header_33 : _GEN_417; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_482 = 3'h3 == encoders_0_io_output ? proc_3_io_next_header_34 : _GEN_418; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_483 = 3'h3 == encoders_0_io_output ? proc_3_io_next_header_35 : _GEN_419; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_484 = 3'h3 == encoders_0_io_output ? proc_3_io_next_header_36 : _GEN_420; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_485 = 3'h3 == encoders_0_io_output ? proc_3_io_next_header_37 : _GEN_421; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_486 = 3'h3 == encoders_0_io_output ? proc_3_io_next_header_38 : _GEN_422; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_487 = 3'h3 == encoders_0_io_output ? proc_3_io_next_header_39 : _GEN_423; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_488 = 3'h3 == encoders_0_io_output ? proc_3_io_next_header_40 : _GEN_424; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_489 = 3'h3 == encoders_0_io_output ? proc_3_io_next_header_41 : _GEN_425; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_490 = 3'h3 == encoders_0_io_output ? proc_3_io_next_header_42 : _GEN_426; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_491 = 3'h3 == encoders_0_io_output ? proc_3_io_next_header_43 : _GEN_427; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_492 = 3'h3 == encoders_0_io_output ? proc_3_io_next_header_44 : _GEN_428; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_493 = 3'h3 == encoders_0_io_output ? proc_3_io_next_header_45 : _GEN_429; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_494 = 3'h3 == encoders_0_io_output ? proc_3_io_next_header_46 : _GEN_430; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_495 = 3'h3 == encoders_0_io_output ? proc_3_io_next_header_47 : _GEN_431; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_496 = 3'h3 == encoders_0_io_output ? proc_3_io_next_header_48 : _GEN_432; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_497 = 3'h3 == encoders_0_io_output ? proc_3_io_next_header_49 : _GEN_433; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_498 = 3'h3 == encoders_0_io_output ? proc_3_io_next_header_50 : _GEN_434; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_499 = 3'h3 == encoders_0_io_output ? proc_3_io_next_header_51 : _GEN_435; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_500 = 3'h3 == encoders_0_io_output ? proc_3_io_next_header_52 : _GEN_436; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_501 = 3'h3 == encoders_0_io_output ? proc_3_io_next_header_53 : _GEN_437; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_502 = 3'h3 == encoders_0_io_output ? proc_3_io_next_header_54 : _GEN_438; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_503 = 3'h3 == encoders_0_io_output ? proc_3_io_next_header_55 : _GEN_439; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_504 = 3'h3 == encoders_0_io_output ? proc_3_io_next_header_56 : _GEN_440; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_505 = 3'h3 == encoders_0_io_output ? proc_3_io_next_header_57 : _GEN_441; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_506 = 3'h3 == encoders_0_io_output ? proc_3_io_next_header_58 : _GEN_442; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_507 = 3'h3 == encoders_0_io_output ? proc_3_io_next_header_59 : _GEN_443; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_508 = 3'h3 == encoders_0_io_output ? proc_3_io_next_header_60 : _GEN_444; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_509 = 3'h3 == encoders_0_io_output ? proc_3_io_next_header_61 : _GEN_445; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_510 = 3'h3 == encoders_0_io_output ? proc_3_io_next_header_62 : _GEN_446; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_511 = 3'h3 == encoders_0_io_output ? proc_3_io_next_header_63 : _GEN_447; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_512 = 3'h4 == encoders_0_io_output ? proc_4_io_next_header_0 : _GEN_448; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_513 = 3'h4 == encoders_0_io_output ? proc_4_io_next_header_1 : _GEN_449; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_514 = 3'h4 == encoders_0_io_output ? proc_4_io_next_header_2 : _GEN_450; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_515 = 3'h4 == encoders_0_io_output ? proc_4_io_next_header_3 : _GEN_451; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_516 = 3'h4 == encoders_0_io_output ? proc_4_io_next_header_4 : _GEN_452; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_517 = 3'h4 == encoders_0_io_output ? proc_4_io_next_header_5 : _GEN_453; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_518 = 3'h4 == encoders_0_io_output ? proc_4_io_next_header_6 : _GEN_454; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_519 = 3'h4 == encoders_0_io_output ? proc_4_io_next_header_7 : _GEN_455; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_520 = 3'h4 == encoders_0_io_output ? proc_4_io_next_header_8 : _GEN_456; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_521 = 3'h4 == encoders_0_io_output ? proc_4_io_next_header_9 : _GEN_457; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_522 = 3'h4 == encoders_0_io_output ? proc_4_io_next_header_10 : _GEN_458; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_523 = 3'h4 == encoders_0_io_output ? proc_4_io_next_header_11 : _GEN_459; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_524 = 3'h4 == encoders_0_io_output ? proc_4_io_next_header_12 : _GEN_460; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_525 = 3'h4 == encoders_0_io_output ? proc_4_io_next_header_13 : _GEN_461; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_526 = 3'h4 == encoders_0_io_output ? proc_4_io_next_header_14 : _GEN_462; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_527 = 3'h4 == encoders_0_io_output ? proc_4_io_next_header_15 : _GEN_463; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_528 = 3'h4 == encoders_0_io_output ? proc_4_io_next_header_16 : _GEN_464; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_529 = 3'h4 == encoders_0_io_output ? proc_4_io_next_header_17 : _GEN_465; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_530 = 3'h4 == encoders_0_io_output ? proc_4_io_next_header_18 : _GEN_466; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_531 = 3'h4 == encoders_0_io_output ? proc_4_io_next_header_19 : _GEN_467; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_532 = 3'h4 == encoders_0_io_output ? proc_4_io_next_header_20 : _GEN_468; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_533 = 3'h4 == encoders_0_io_output ? proc_4_io_next_header_21 : _GEN_469; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_534 = 3'h4 == encoders_0_io_output ? proc_4_io_next_header_22 : _GEN_470; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_535 = 3'h4 == encoders_0_io_output ? proc_4_io_next_header_23 : _GEN_471; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_536 = 3'h4 == encoders_0_io_output ? proc_4_io_next_header_24 : _GEN_472; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_537 = 3'h4 == encoders_0_io_output ? proc_4_io_next_header_25 : _GEN_473; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_538 = 3'h4 == encoders_0_io_output ? proc_4_io_next_header_26 : _GEN_474; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_539 = 3'h4 == encoders_0_io_output ? proc_4_io_next_header_27 : _GEN_475; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_540 = 3'h4 == encoders_0_io_output ? proc_4_io_next_header_28 : _GEN_476; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_541 = 3'h4 == encoders_0_io_output ? proc_4_io_next_header_29 : _GEN_477; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_542 = 3'h4 == encoders_0_io_output ? proc_4_io_next_header_30 : _GEN_478; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_543 = 3'h4 == encoders_0_io_output ? proc_4_io_next_header_31 : _GEN_479; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_544 = 3'h4 == encoders_0_io_output ? proc_4_io_next_header_32 : _GEN_480; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_545 = 3'h4 == encoders_0_io_output ? proc_4_io_next_header_33 : _GEN_481; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_546 = 3'h4 == encoders_0_io_output ? proc_4_io_next_header_34 : _GEN_482; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_547 = 3'h4 == encoders_0_io_output ? proc_4_io_next_header_35 : _GEN_483; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_548 = 3'h4 == encoders_0_io_output ? proc_4_io_next_header_36 : _GEN_484; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_549 = 3'h4 == encoders_0_io_output ? proc_4_io_next_header_37 : _GEN_485; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_550 = 3'h4 == encoders_0_io_output ? proc_4_io_next_header_38 : _GEN_486; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_551 = 3'h4 == encoders_0_io_output ? proc_4_io_next_header_39 : _GEN_487; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_552 = 3'h4 == encoders_0_io_output ? proc_4_io_next_header_40 : _GEN_488; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_553 = 3'h4 == encoders_0_io_output ? proc_4_io_next_header_41 : _GEN_489; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_554 = 3'h4 == encoders_0_io_output ? proc_4_io_next_header_42 : _GEN_490; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_555 = 3'h4 == encoders_0_io_output ? proc_4_io_next_header_43 : _GEN_491; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_556 = 3'h4 == encoders_0_io_output ? proc_4_io_next_header_44 : _GEN_492; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_557 = 3'h4 == encoders_0_io_output ? proc_4_io_next_header_45 : _GEN_493; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_558 = 3'h4 == encoders_0_io_output ? proc_4_io_next_header_46 : _GEN_494; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_559 = 3'h4 == encoders_0_io_output ? proc_4_io_next_header_47 : _GEN_495; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_560 = 3'h4 == encoders_0_io_output ? proc_4_io_next_header_48 : _GEN_496; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_561 = 3'h4 == encoders_0_io_output ? proc_4_io_next_header_49 : _GEN_497; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_562 = 3'h4 == encoders_0_io_output ? proc_4_io_next_header_50 : _GEN_498; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_563 = 3'h4 == encoders_0_io_output ? proc_4_io_next_header_51 : _GEN_499; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_564 = 3'h4 == encoders_0_io_output ? proc_4_io_next_header_52 : _GEN_500; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_565 = 3'h4 == encoders_0_io_output ? proc_4_io_next_header_53 : _GEN_501; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_566 = 3'h4 == encoders_0_io_output ? proc_4_io_next_header_54 : _GEN_502; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_567 = 3'h4 == encoders_0_io_output ? proc_4_io_next_header_55 : _GEN_503; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_568 = 3'h4 == encoders_0_io_output ? proc_4_io_next_header_56 : _GEN_504; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_569 = 3'h4 == encoders_0_io_output ? proc_4_io_next_header_57 : _GEN_505; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_570 = 3'h4 == encoders_0_io_output ? proc_4_io_next_header_58 : _GEN_506; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_571 = 3'h4 == encoders_0_io_output ? proc_4_io_next_header_59 : _GEN_507; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_572 = 3'h4 == encoders_0_io_output ? proc_4_io_next_header_60 : _GEN_508; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_573 = 3'h4 == encoders_0_io_output ? proc_4_io_next_header_61 : _GEN_509; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_574 = 3'h4 == encoders_0_io_output ? proc_4_io_next_header_62 : _GEN_510; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_575 = 3'h4 == encoders_0_io_output ? proc_4_io_next_header_63 : _GEN_511; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_576 = 3'h5 == encoders_0_io_output ? proc_5_io_next_header_0 : _GEN_512; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_577 = 3'h5 == encoders_0_io_output ? proc_5_io_next_header_1 : _GEN_513; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_578 = 3'h5 == encoders_0_io_output ? proc_5_io_next_header_2 : _GEN_514; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_579 = 3'h5 == encoders_0_io_output ? proc_5_io_next_header_3 : _GEN_515; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_580 = 3'h5 == encoders_0_io_output ? proc_5_io_next_header_4 : _GEN_516; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_581 = 3'h5 == encoders_0_io_output ? proc_5_io_next_header_5 : _GEN_517; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_582 = 3'h5 == encoders_0_io_output ? proc_5_io_next_header_6 : _GEN_518; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_583 = 3'h5 == encoders_0_io_output ? proc_5_io_next_header_7 : _GEN_519; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_584 = 3'h5 == encoders_0_io_output ? proc_5_io_next_header_8 : _GEN_520; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_585 = 3'h5 == encoders_0_io_output ? proc_5_io_next_header_9 : _GEN_521; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_586 = 3'h5 == encoders_0_io_output ? proc_5_io_next_header_10 : _GEN_522; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_587 = 3'h5 == encoders_0_io_output ? proc_5_io_next_header_11 : _GEN_523; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_588 = 3'h5 == encoders_0_io_output ? proc_5_io_next_header_12 : _GEN_524; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_589 = 3'h5 == encoders_0_io_output ? proc_5_io_next_header_13 : _GEN_525; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_590 = 3'h5 == encoders_0_io_output ? proc_5_io_next_header_14 : _GEN_526; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_591 = 3'h5 == encoders_0_io_output ? proc_5_io_next_header_15 : _GEN_527; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_592 = 3'h5 == encoders_0_io_output ? proc_5_io_next_header_16 : _GEN_528; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_593 = 3'h5 == encoders_0_io_output ? proc_5_io_next_header_17 : _GEN_529; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_594 = 3'h5 == encoders_0_io_output ? proc_5_io_next_header_18 : _GEN_530; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_595 = 3'h5 == encoders_0_io_output ? proc_5_io_next_header_19 : _GEN_531; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_596 = 3'h5 == encoders_0_io_output ? proc_5_io_next_header_20 : _GEN_532; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_597 = 3'h5 == encoders_0_io_output ? proc_5_io_next_header_21 : _GEN_533; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_598 = 3'h5 == encoders_0_io_output ? proc_5_io_next_header_22 : _GEN_534; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_599 = 3'h5 == encoders_0_io_output ? proc_5_io_next_header_23 : _GEN_535; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_600 = 3'h5 == encoders_0_io_output ? proc_5_io_next_header_24 : _GEN_536; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_601 = 3'h5 == encoders_0_io_output ? proc_5_io_next_header_25 : _GEN_537; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_602 = 3'h5 == encoders_0_io_output ? proc_5_io_next_header_26 : _GEN_538; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_603 = 3'h5 == encoders_0_io_output ? proc_5_io_next_header_27 : _GEN_539; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_604 = 3'h5 == encoders_0_io_output ? proc_5_io_next_header_28 : _GEN_540; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_605 = 3'h5 == encoders_0_io_output ? proc_5_io_next_header_29 : _GEN_541; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_606 = 3'h5 == encoders_0_io_output ? proc_5_io_next_header_30 : _GEN_542; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_607 = 3'h5 == encoders_0_io_output ? proc_5_io_next_header_31 : _GEN_543; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_608 = 3'h5 == encoders_0_io_output ? proc_5_io_next_header_32 : _GEN_544; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_609 = 3'h5 == encoders_0_io_output ? proc_5_io_next_header_33 : _GEN_545; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_610 = 3'h5 == encoders_0_io_output ? proc_5_io_next_header_34 : _GEN_546; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_611 = 3'h5 == encoders_0_io_output ? proc_5_io_next_header_35 : _GEN_547; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_612 = 3'h5 == encoders_0_io_output ? proc_5_io_next_header_36 : _GEN_548; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_613 = 3'h5 == encoders_0_io_output ? proc_5_io_next_header_37 : _GEN_549; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_614 = 3'h5 == encoders_0_io_output ? proc_5_io_next_header_38 : _GEN_550; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_615 = 3'h5 == encoders_0_io_output ? proc_5_io_next_header_39 : _GEN_551; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_616 = 3'h5 == encoders_0_io_output ? proc_5_io_next_header_40 : _GEN_552; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_617 = 3'h5 == encoders_0_io_output ? proc_5_io_next_header_41 : _GEN_553; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_618 = 3'h5 == encoders_0_io_output ? proc_5_io_next_header_42 : _GEN_554; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_619 = 3'h5 == encoders_0_io_output ? proc_5_io_next_header_43 : _GEN_555; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_620 = 3'h5 == encoders_0_io_output ? proc_5_io_next_header_44 : _GEN_556; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_621 = 3'h5 == encoders_0_io_output ? proc_5_io_next_header_45 : _GEN_557; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_622 = 3'h5 == encoders_0_io_output ? proc_5_io_next_header_46 : _GEN_558; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_623 = 3'h5 == encoders_0_io_output ? proc_5_io_next_header_47 : _GEN_559; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_624 = 3'h5 == encoders_0_io_output ? proc_5_io_next_header_48 : _GEN_560; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_625 = 3'h5 == encoders_0_io_output ? proc_5_io_next_header_49 : _GEN_561; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_626 = 3'h5 == encoders_0_io_output ? proc_5_io_next_header_50 : _GEN_562; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_627 = 3'h5 == encoders_0_io_output ? proc_5_io_next_header_51 : _GEN_563; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_628 = 3'h5 == encoders_0_io_output ? proc_5_io_next_header_52 : _GEN_564; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_629 = 3'h5 == encoders_0_io_output ? proc_5_io_next_header_53 : _GEN_565; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_630 = 3'h5 == encoders_0_io_output ? proc_5_io_next_header_54 : _GEN_566; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_631 = 3'h5 == encoders_0_io_output ? proc_5_io_next_header_55 : _GEN_567; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_632 = 3'h5 == encoders_0_io_output ? proc_5_io_next_header_56 : _GEN_568; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_633 = 3'h5 == encoders_0_io_output ? proc_5_io_next_header_57 : _GEN_569; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_634 = 3'h5 == encoders_0_io_output ? proc_5_io_next_header_58 : _GEN_570; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_635 = 3'h5 == encoders_0_io_output ? proc_5_io_next_header_59 : _GEN_571; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_636 = 3'h5 == encoders_0_io_output ? proc_5_io_next_header_60 : _GEN_572; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_637 = 3'h5 == encoders_0_io_output ? proc_5_io_next_header_61 : _GEN_573; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_638 = 3'h5 == encoders_0_io_output ? proc_5_io_next_header_62 : _GEN_574; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_639 = 3'h5 == encoders_0_io_output ? proc_5_io_next_header_63 : _GEN_575; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_640 = 3'h6 == encoders_0_io_output ? proc_6_io_next_header_0 : _GEN_576; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_641 = 3'h6 == encoders_0_io_output ? proc_6_io_next_header_1 : _GEN_577; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_642 = 3'h6 == encoders_0_io_output ? proc_6_io_next_header_2 : _GEN_578; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_643 = 3'h6 == encoders_0_io_output ? proc_6_io_next_header_3 : _GEN_579; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_644 = 3'h6 == encoders_0_io_output ? proc_6_io_next_header_4 : _GEN_580; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_645 = 3'h6 == encoders_0_io_output ? proc_6_io_next_header_5 : _GEN_581; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_646 = 3'h6 == encoders_0_io_output ? proc_6_io_next_header_6 : _GEN_582; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_647 = 3'h6 == encoders_0_io_output ? proc_6_io_next_header_7 : _GEN_583; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_648 = 3'h6 == encoders_0_io_output ? proc_6_io_next_header_8 : _GEN_584; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_649 = 3'h6 == encoders_0_io_output ? proc_6_io_next_header_9 : _GEN_585; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_650 = 3'h6 == encoders_0_io_output ? proc_6_io_next_header_10 : _GEN_586; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_651 = 3'h6 == encoders_0_io_output ? proc_6_io_next_header_11 : _GEN_587; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_652 = 3'h6 == encoders_0_io_output ? proc_6_io_next_header_12 : _GEN_588; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_653 = 3'h6 == encoders_0_io_output ? proc_6_io_next_header_13 : _GEN_589; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_654 = 3'h6 == encoders_0_io_output ? proc_6_io_next_header_14 : _GEN_590; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_655 = 3'h6 == encoders_0_io_output ? proc_6_io_next_header_15 : _GEN_591; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_656 = 3'h6 == encoders_0_io_output ? proc_6_io_next_header_16 : _GEN_592; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_657 = 3'h6 == encoders_0_io_output ? proc_6_io_next_header_17 : _GEN_593; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_658 = 3'h6 == encoders_0_io_output ? proc_6_io_next_header_18 : _GEN_594; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_659 = 3'h6 == encoders_0_io_output ? proc_6_io_next_header_19 : _GEN_595; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_660 = 3'h6 == encoders_0_io_output ? proc_6_io_next_header_20 : _GEN_596; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_661 = 3'h6 == encoders_0_io_output ? proc_6_io_next_header_21 : _GEN_597; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_662 = 3'h6 == encoders_0_io_output ? proc_6_io_next_header_22 : _GEN_598; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_663 = 3'h6 == encoders_0_io_output ? proc_6_io_next_header_23 : _GEN_599; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_664 = 3'h6 == encoders_0_io_output ? proc_6_io_next_header_24 : _GEN_600; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_665 = 3'h6 == encoders_0_io_output ? proc_6_io_next_header_25 : _GEN_601; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_666 = 3'h6 == encoders_0_io_output ? proc_6_io_next_header_26 : _GEN_602; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_667 = 3'h6 == encoders_0_io_output ? proc_6_io_next_header_27 : _GEN_603; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_668 = 3'h6 == encoders_0_io_output ? proc_6_io_next_header_28 : _GEN_604; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_669 = 3'h6 == encoders_0_io_output ? proc_6_io_next_header_29 : _GEN_605; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_670 = 3'h6 == encoders_0_io_output ? proc_6_io_next_header_30 : _GEN_606; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_671 = 3'h6 == encoders_0_io_output ? proc_6_io_next_header_31 : _GEN_607; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_672 = 3'h6 == encoders_0_io_output ? proc_6_io_next_header_32 : _GEN_608; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_673 = 3'h6 == encoders_0_io_output ? proc_6_io_next_header_33 : _GEN_609; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_674 = 3'h6 == encoders_0_io_output ? proc_6_io_next_header_34 : _GEN_610; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_675 = 3'h6 == encoders_0_io_output ? proc_6_io_next_header_35 : _GEN_611; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_676 = 3'h6 == encoders_0_io_output ? proc_6_io_next_header_36 : _GEN_612; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_677 = 3'h6 == encoders_0_io_output ? proc_6_io_next_header_37 : _GEN_613; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_678 = 3'h6 == encoders_0_io_output ? proc_6_io_next_header_38 : _GEN_614; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_679 = 3'h6 == encoders_0_io_output ? proc_6_io_next_header_39 : _GEN_615; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_680 = 3'h6 == encoders_0_io_output ? proc_6_io_next_header_40 : _GEN_616; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_681 = 3'h6 == encoders_0_io_output ? proc_6_io_next_header_41 : _GEN_617; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_682 = 3'h6 == encoders_0_io_output ? proc_6_io_next_header_42 : _GEN_618; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_683 = 3'h6 == encoders_0_io_output ? proc_6_io_next_header_43 : _GEN_619; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_684 = 3'h6 == encoders_0_io_output ? proc_6_io_next_header_44 : _GEN_620; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_685 = 3'h6 == encoders_0_io_output ? proc_6_io_next_header_45 : _GEN_621; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_686 = 3'h6 == encoders_0_io_output ? proc_6_io_next_header_46 : _GEN_622; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_687 = 3'h6 == encoders_0_io_output ? proc_6_io_next_header_47 : _GEN_623; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_688 = 3'h6 == encoders_0_io_output ? proc_6_io_next_header_48 : _GEN_624; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_689 = 3'h6 == encoders_0_io_output ? proc_6_io_next_header_49 : _GEN_625; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_690 = 3'h6 == encoders_0_io_output ? proc_6_io_next_header_50 : _GEN_626; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_691 = 3'h6 == encoders_0_io_output ? proc_6_io_next_header_51 : _GEN_627; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_692 = 3'h6 == encoders_0_io_output ? proc_6_io_next_header_52 : _GEN_628; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_693 = 3'h6 == encoders_0_io_output ? proc_6_io_next_header_53 : _GEN_629; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_694 = 3'h6 == encoders_0_io_output ? proc_6_io_next_header_54 : _GEN_630; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_695 = 3'h6 == encoders_0_io_output ? proc_6_io_next_header_55 : _GEN_631; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_696 = 3'h6 == encoders_0_io_output ? proc_6_io_next_header_56 : _GEN_632; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_697 = 3'h6 == encoders_0_io_output ? proc_6_io_next_header_57 : _GEN_633; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_698 = 3'h6 == encoders_0_io_output ? proc_6_io_next_header_58 : _GEN_634; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_699 = 3'h6 == encoders_0_io_output ? proc_6_io_next_header_59 : _GEN_635; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_700 = 3'h6 == encoders_0_io_output ? proc_6_io_next_header_60 : _GEN_636; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_701 = 3'h6 == encoders_0_io_output ? proc_6_io_next_header_61 : _GEN_637; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_702 = 3'h6 == encoders_0_io_output ? proc_6_io_next_header_62 : _GEN_638; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_703 = 3'h6 == encoders_0_io_output ? proc_6_io_next_header_63 : _GEN_639; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_704 = 3'h7 == encoders_0_io_output ? proc_7_io_next_header_0 : _GEN_640; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_705 = 3'h7 == encoders_0_io_output ? proc_7_io_next_header_1 : _GEN_641; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_706 = 3'h7 == encoders_0_io_output ? proc_7_io_next_header_2 : _GEN_642; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_707 = 3'h7 == encoders_0_io_output ? proc_7_io_next_header_3 : _GEN_643; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_708 = 3'h7 == encoders_0_io_output ? proc_7_io_next_header_4 : _GEN_644; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_709 = 3'h7 == encoders_0_io_output ? proc_7_io_next_header_5 : _GEN_645; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_710 = 3'h7 == encoders_0_io_output ? proc_7_io_next_header_6 : _GEN_646; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_711 = 3'h7 == encoders_0_io_output ? proc_7_io_next_header_7 : _GEN_647; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_712 = 3'h7 == encoders_0_io_output ? proc_7_io_next_header_8 : _GEN_648; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_713 = 3'h7 == encoders_0_io_output ? proc_7_io_next_header_9 : _GEN_649; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_714 = 3'h7 == encoders_0_io_output ? proc_7_io_next_header_10 : _GEN_650; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_715 = 3'h7 == encoders_0_io_output ? proc_7_io_next_header_11 : _GEN_651; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_716 = 3'h7 == encoders_0_io_output ? proc_7_io_next_header_12 : _GEN_652; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_717 = 3'h7 == encoders_0_io_output ? proc_7_io_next_header_13 : _GEN_653; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_718 = 3'h7 == encoders_0_io_output ? proc_7_io_next_header_14 : _GEN_654; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_719 = 3'h7 == encoders_0_io_output ? proc_7_io_next_header_15 : _GEN_655; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_720 = 3'h7 == encoders_0_io_output ? proc_7_io_next_header_16 : _GEN_656; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_721 = 3'h7 == encoders_0_io_output ? proc_7_io_next_header_17 : _GEN_657; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_722 = 3'h7 == encoders_0_io_output ? proc_7_io_next_header_18 : _GEN_658; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_723 = 3'h7 == encoders_0_io_output ? proc_7_io_next_header_19 : _GEN_659; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_724 = 3'h7 == encoders_0_io_output ? proc_7_io_next_header_20 : _GEN_660; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_725 = 3'h7 == encoders_0_io_output ? proc_7_io_next_header_21 : _GEN_661; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_726 = 3'h7 == encoders_0_io_output ? proc_7_io_next_header_22 : _GEN_662; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_727 = 3'h7 == encoders_0_io_output ? proc_7_io_next_header_23 : _GEN_663; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_728 = 3'h7 == encoders_0_io_output ? proc_7_io_next_header_24 : _GEN_664; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_729 = 3'h7 == encoders_0_io_output ? proc_7_io_next_header_25 : _GEN_665; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_730 = 3'h7 == encoders_0_io_output ? proc_7_io_next_header_26 : _GEN_666; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_731 = 3'h7 == encoders_0_io_output ? proc_7_io_next_header_27 : _GEN_667; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_732 = 3'h7 == encoders_0_io_output ? proc_7_io_next_header_28 : _GEN_668; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_733 = 3'h7 == encoders_0_io_output ? proc_7_io_next_header_29 : _GEN_669; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_734 = 3'h7 == encoders_0_io_output ? proc_7_io_next_header_30 : _GEN_670; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_735 = 3'h7 == encoders_0_io_output ? proc_7_io_next_header_31 : _GEN_671; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_736 = 3'h7 == encoders_0_io_output ? proc_7_io_next_header_32 : _GEN_672; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_737 = 3'h7 == encoders_0_io_output ? proc_7_io_next_header_33 : _GEN_673; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_738 = 3'h7 == encoders_0_io_output ? proc_7_io_next_header_34 : _GEN_674; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_739 = 3'h7 == encoders_0_io_output ? proc_7_io_next_header_35 : _GEN_675; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_740 = 3'h7 == encoders_0_io_output ? proc_7_io_next_header_36 : _GEN_676; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_741 = 3'h7 == encoders_0_io_output ? proc_7_io_next_header_37 : _GEN_677; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_742 = 3'h7 == encoders_0_io_output ? proc_7_io_next_header_38 : _GEN_678; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_743 = 3'h7 == encoders_0_io_output ? proc_7_io_next_header_39 : _GEN_679; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_744 = 3'h7 == encoders_0_io_output ? proc_7_io_next_header_40 : _GEN_680; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_745 = 3'h7 == encoders_0_io_output ? proc_7_io_next_header_41 : _GEN_681; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_746 = 3'h7 == encoders_0_io_output ? proc_7_io_next_header_42 : _GEN_682; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_747 = 3'h7 == encoders_0_io_output ? proc_7_io_next_header_43 : _GEN_683; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_748 = 3'h7 == encoders_0_io_output ? proc_7_io_next_header_44 : _GEN_684; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_749 = 3'h7 == encoders_0_io_output ? proc_7_io_next_header_45 : _GEN_685; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_750 = 3'h7 == encoders_0_io_output ? proc_7_io_next_header_46 : _GEN_686; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_751 = 3'h7 == encoders_0_io_output ? proc_7_io_next_header_47 : _GEN_687; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_752 = 3'h7 == encoders_0_io_output ? proc_7_io_next_header_48 : _GEN_688; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_753 = 3'h7 == encoders_0_io_output ? proc_7_io_next_header_49 : _GEN_689; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_754 = 3'h7 == encoders_0_io_output ? proc_7_io_next_header_50 : _GEN_690; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_755 = 3'h7 == encoders_0_io_output ? proc_7_io_next_header_51 : _GEN_691; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_756 = 3'h7 == encoders_0_io_output ? proc_7_io_next_header_52 : _GEN_692; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_757 = 3'h7 == encoders_0_io_output ? proc_7_io_next_header_53 : _GEN_693; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_758 = 3'h7 == encoders_0_io_output ? proc_7_io_next_header_54 : _GEN_694; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_759 = 3'h7 == encoders_0_io_output ? proc_7_io_next_header_55 : _GEN_695; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_760 = 3'h7 == encoders_0_io_output ? proc_7_io_next_header_56 : _GEN_696; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_761 = 3'h7 == encoders_0_io_output ? proc_7_io_next_header_57 : _GEN_697; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_762 = 3'h7 == encoders_0_io_output ? proc_7_io_next_header_58 : _GEN_698; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_763 = 3'h7 == encoders_0_io_output ? proc_7_io_next_header_59 : _GEN_699; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_764 = 3'h7 == encoders_0_io_output ? proc_7_io_next_header_60 : _GEN_700; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_765 = 3'h7 == encoders_0_io_output ? proc_7_io_next_header_61 : _GEN_701; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_766 = 3'h7 == encoders_0_io_output ? proc_7_io_next_header_62 : _GEN_702; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_767 = 3'h7 == encoders_0_io_output ? proc_7_io_next_header_63 : _GEN_703; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_834 = 3'h0 == encoders_1_io_output ? proc_0_io_next_header_0 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_835 = 3'h0 == encoders_1_io_output ? proc_0_io_next_header_1 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_836 = 3'h0 == encoders_1_io_output ? proc_0_io_next_header_2 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_837 = 3'h0 == encoders_1_io_output ? proc_0_io_next_header_3 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_838 = 3'h0 == encoders_1_io_output ? proc_0_io_next_header_4 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_839 = 3'h0 == encoders_1_io_output ? proc_0_io_next_header_5 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_840 = 3'h0 == encoders_1_io_output ? proc_0_io_next_header_6 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_841 = 3'h0 == encoders_1_io_output ? proc_0_io_next_header_7 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_842 = 3'h0 == encoders_1_io_output ? proc_0_io_next_header_8 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_843 = 3'h0 == encoders_1_io_output ? proc_0_io_next_header_9 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_844 = 3'h0 == encoders_1_io_output ? proc_0_io_next_header_10 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_845 = 3'h0 == encoders_1_io_output ? proc_0_io_next_header_11 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_846 = 3'h0 == encoders_1_io_output ? proc_0_io_next_header_12 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_847 = 3'h0 == encoders_1_io_output ? proc_0_io_next_header_13 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_848 = 3'h0 == encoders_1_io_output ? proc_0_io_next_header_14 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_849 = 3'h0 == encoders_1_io_output ? proc_0_io_next_header_15 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_850 = 3'h0 == encoders_1_io_output ? proc_0_io_next_header_16 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_851 = 3'h0 == encoders_1_io_output ? proc_0_io_next_header_17 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_852 = 3'h0 == encoders_1_io_output ? proc_0_io_next_header_18 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_853 = 3'h0 == encoders_1_io_output ? proc_0_io_next_header_19 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_854 = 3'h0 == encoders_1_io_output ? proc_0_io_next_header_20 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_855 = 3'h0 == encoders_1_io_output ? proc_0_io_next_header_21 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_856 = 3'h0 == encoders_1_io_output ? proc_0_io_next_header_22 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_857 = 3'h0 == encoders_1_io_output ? proc_0_io_next_header_23 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_858 = 3'h0 == encoders_1_io_output ? proc_0_io_next_header_24 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_859 = 3'h0 == encoders_1_io_output ? proc_0_io_next_header_25 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_860 = 3'h0 == encoders_1_io_output ? proc_0_io_next_header_26 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_861 = 3'h0 == encoders_1_io_output ? proc_0_io_next_header_27 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_862 = 3'h0 == encoders_1_io_output ? proc_0_io_next_header_28 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_863 = 3'h0 == encoders_1_io_output ? proc_0_io_next_header_29 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_864 = 3'h0 == encoders_1_io_output ? proc_0_io_next_header_30 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_865 = 3'h0 == encoders_1_io_output ? proc_0_io_next_header_31 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_866 = 3'h0 == encoders_1_io_output ? proc_0_io_next_header_32 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_867 = 3'h0 == encoders_1_io_output ? proc_0_io_next_header_33 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_868 = 3'h0 == encoders_1_io_output ? proc_0_io_next_header_34 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_869 = 3'h0 == encoders_1_io_output ? proc_0_io_next_header_35 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_870 = 3'h0 == encoders_1_io_output ? proc_0_io_next_header_36 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_871 = 3'h0 == encoders_1_io_output ? proc_0_io_next_header_37 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_872 = 3'h0 == encoders_1_io_output ? proc_0_io_next_header_38 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_873 = 3'h0 == encoders_1_io_output ? proc_0_io_next_header_39 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_874 = 3'h0 == encoders_1_io_output ? proc_0_io_next_header_40 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_875 = 3'h0 == encoders_1_io_output ? proc_0_io_next_header_41 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_876 = 3'h0 == encoders_1_io_output ? proc_0_io_next_header_42 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_877 = 3'h0 == encoders_1_io_output ? proc_0_io_next_header_43 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_878 = 3'h0 == encoders_1_io_output ? proc_0_io_next_header_44 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_879 = 3'h0 == encoders_1_io_output ? proc_0_io_next_header_45 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_880 = 3'h0 == encoders_1_io_output ? proc_0_io_next_header_46 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_881 = 3'h0 == encoders_1_io_output ? proc_0_io_next_header_47 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_882 = 3'h0 == encoders_1_io_output ? proc_0_io_next_header_48 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_883 = 3'h0 == encoders_1_io_output ? proc_0_io_next_header_49 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_884 = 3'h0 == encoders_1_io_output ? proc_0_io_next_header_50 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_885 = 3'h0 == encoders_1_io_output ? proc_0_io_next_header_51 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_886 = 3'h0 == encoders_1_io_output ? proc_0_io_next_header_52 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_887 = 3'h0 == encoders_1_io_output ? proc_0_io_next_header_53 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_888 = 3'h0 == encoders_1_io_output ? proc_0_io_next_header_54 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_889 = 3'h0 == encoders_1_io_output ? proc_0_io_next_header_55 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_890 = 3'h0 == encoders_1_io_output ? proc_0_io_next_header_56 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_891 = 3'h0 == encoders_1_io_output ? proc_0_io_next_header_57 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_892 = 3'h0 == encoders_1_io_output ? proc_0_io_next_header_58 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_893 = 3'h0 == encoders_1_io_output ? proc_0_io_next_header_59 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_894 = 3'h0 == encoders_1_io_output ? proc_0_io_next_header_60 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_895 = 3'h0 == encoders_1_io_output ? proc_0_io_next_header_61 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_896 = 3'h0 == encoders_1_io_output ? proc_0_io_next_header_62 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_897 = 3'h0 == encoders_1_io_output ? proc_0_io_next_header_63 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_898 = 3'h1 == encoders_1_io_output ? proc_1_io_next_header_0 : _GEN_834; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_899 = 3'h1 == encoders_1_io_output ? proc_1_io_next_header_1 : _GEN_835; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_900 = 3'h1 == encoders_1_io_output ? proc_1_io_next_header_2 : _GEN_836; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_901 = 3'h1 == encoders_1_io_output ? proc_1_io_next_header_3 : _GEN_837; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_902 = 3'h1 == encoders_1_io_output ? proc_1_io_next_header_4 : _GEN_838; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_903 = 3'h1 == encoders_1_io_output ? proc_1_io_next_header_5 : _GEN_839; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_904 = 3'h1 == encoders_1_io_output ? proc_1_io_next_header_6 : _GEN_840; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_905 = 3'h1 == encoders_1_io_output ? proc_1_io_next_header_7 : _GEN_841; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_906 = 3'h1 == encoders_1_io_output ? proc_1_io_next_header_8 : _GEN_842; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_907 = 3'h1 == encoders_1_io_output ? proc_1_io_next_header_9 : _GEN_843; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_908 = 3'h1 == encoders_1_io_output ? proc_1_io_next_header_10 : _GEN_844; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_909 = 3'h1 == encoders_1_io_output ? proc_1_io_next_header_11 : _GEN_845; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_910 = 3'h1 == encoders_1_io_output ? proc_1_io_next_header_12 : _GEN_846; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_911 = 3'h1 == encoders_1_io_output ? proc_1_io_next_header_13 : _GEN_847; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_912 = 3'h1 == encoders_1_io_output ? proc_1_io_next_header_14 : _GEN_848; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_913 = 3'h1 == encoders_1_io_output ? proc_1_io_next_header_15 : _GEN_849; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_914 = 3'h1 == encoders_1_io_output ? proc_1_io_next_header_16 : _GEN_850; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_915 = 3'h1 == encoders_1_io_output ? proc_1_io_next_header_17 : _GEN_851; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_916 = 3'h1 == encoders_1_io_output ? proc_1_io_next_header_18 : _GEN_852; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_917 = 3'h1 == encoders_1_io_output ? proc_1_io_next_header_19 : _GEN_853; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_918 = 3'h1 == encoders_1_io_output ? proc_1_io_next_header_20 : _GEN_854; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_919 = 3'h1 == encoders_1_io_output ? proc_1_io_next_header_21 : _GEN_855; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_920 = 3'h1 == encoders_1_io_output ? proc_1_io_next_header_22 : _GEN_856; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_921 = 3'h1 == encoders_1_io_output ? proc_1_io_next_header_23 : _GEN_857; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_922 = 3'h1 == encoders_1_io_output ? proc_1_io_next_header_24 : _GEN_858; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_923 = 3'h1 == encoders_1_io_output ? proc_1_io_next_header_25 : _GEN_859; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_924 = 3'h1 == encoders_1_io_output ? proc_1_io_next_header_26 : _GEN_860; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_925 = 3'h1 == encoders_1_io_output ? proc_1_io_next_header_27 : _GEN_861; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_926 = 3'h1 == encoders_1_io_output ? proc_1_io_next_header_28 : _GEN_862; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_927 = 3'h1 == encoders_1_io_output ? proc_1_io_next_header_29 : _GEN_863; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_928 = 3'h1 == encoders_1_io_output ? proc_1_io_next_header_30 : _GEN_864; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_929 = 3'h1 == encoders_1_io_output ? proc_1_io_next_header_31 : _GEN_865; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_930 = 3'h1 == encoders_1_io_output ? proc_1_io_next_header_32 : _GEN_866; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_931 = 3'h1 == encoders_1_io_output ? proc_1_io_next_header_33 : _GEN_867; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_932 = 3'h1 == encoders_1_io_output ? proc_1_io_next_header_34 : _GEN_868; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_933 = 3'h1 == encoders_1_io_output ? proc_1_io_next_header_35 : _GEN_869; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_934 = 3'h1 == encoders_1_io_output ? proc_1_io_next_header_36 : _GEN_870; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_935 = 3'h1 == encoders_1_io_output ? proc_1_io_next_header_37 : _GEN_871; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_936 = 3'h1 == encoders_1_io_output ? proc_1_io_next_header_38 : _GEN_872; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_937 = 3'h1 == encoders_1_io_output ? proc_1_io_next_header_39 : _GEN_873; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_938 = 3'h1 == encoders_1_io_output ? proc_1_io_next_header_40 : _GEN_874; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_939 = 3'h1 == encoders_1_io_output ? proc_1_io_next_header_41 : _GEN_875; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_940 = 3'h1 == encoders_1_io_output ? proc_1_io_next_header_42 : _GEN_876; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_941 = 3'h1 == encoders_1_io_output ? proc_1_io_next_header_43 : _GEN_877; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_942 = 3'h1 == encoders_1_io_output ? proc_1_io_next_header_44 : _GEN_878; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_943 = 3'h1 == encoders_1_io_output ? proc_1_io_next_header_45 : _GEN_879; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_944 = 3'h1 == encoders_1_io_output ? proc_1_io_next_header_46 : _GEN_880; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_945 = 3'h1 == encoders_1_io_output ? proc_1_io_next_header_47 : _GEN_881; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_946 = 3'h1 == encoders_1_io_output ? proc_1_io_next_header_48 : _GEN_882; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_947 = 3'h1 == encoders_1_io_output ? proc_1_io_next_header_49 : _GEN_883; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_948 = 3'h1 == encoders_1_io_output ? proc_1_io_next_header_50 : _GEN_884; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_949 = 3'h1 == encoders_1_io_output ? proc_1_io_next_header_51 : _GEN_885; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_950 = 3'h1 == encoders_1_io_output ? proc_1_io_next_header_52 : _GEN_886; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_951 = 3'h1 == encoders_1_io_output ? proc_1_io_next_header_53 : _GEN_887; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_952 = 3'h1 == encoders_1_io_output ? proc_1_io_next_header_54 : _GEN_888; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_953 = 3'h1 == encoders_1_io_output ? proc_1_io_next_header_55 : _GEN_889; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_954 = 3'h1 == encoders_1_io_output ? proc_1_io_next_header_56 : _GEN_890; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_955 = 3'h1 == encoders_1_io_output ? proc_1_io_next_header_57 : _GEN_891; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_956 = 3'h1 == encoders_1_io_output ? proc_1_io_next_header_58 : _GEN_892; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_957 = 3'h1 == encoders_1_io_output ? proc_1_io_next_header_59 : _GEN_893; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_958 = 3'h1 == encoders_1_io_output ? proc_1_io_next_header_60 : _GEN_894; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_959 = 3'h1 == encoders_1_io_output ? proc_1_io_next_header_61 : _GEN_895; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_960 = 3'h1 == encoders_1_io_output ? proc_1_io_next_header_62 : _GEN_896; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_961 = 3'h1 == encoders_1_io_output ? proc_1_io_next_header_63 : _GEN_897; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_962 = 3'h2 == encoders_1_io_output ? proc_2_io_next_header_0 : _GEN_898; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_963 = 3'h2 == encoders_1_io_output ? proc_2_io_next_header_1 : _GEN_899; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_964 = 3'h2 == encoders_1_io_output ? proc_2_io_next_header_2 : _GEN_900; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_965 = 3'h2 == encoders_1_io_output ? proc_2_io_next_header_3 : _GEN_901; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_966 = 3'h2 == encoders_1_io_output ? proc_2_io_next_header_4 : _GEN_902; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_967 = 3'h2 == encoders_1_io_output ? proc_2_io_next_header_5 : _GEN_903; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_968 = 3'h2 == encoders_1_io_output ? proc_2_io_next_header_6 : _GEN_904; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_969 = 3'h2 == encoders_1_io_output ? proc_2_io_next_header_7 : _GEN_905; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_970 = 3'h2 == encoders_1_io_output ? proc_2_io_next_header_8 : _GEN_906; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_971 = 3'h2 == encoders_1_io_output ? proc_2_io_next_header_9 : _GEN_907; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_972 = 3'h2 == encoders_1_io_output ? proc_2_io_next_header_10 : _GEN_908; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_973 = 3'h2 == encoders_1_io_output ? proc_2_io_next_header_11 : _GEN_909; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_974 = 3'h2 == encoders_1_io_output ? proc_2_io_next_header_12 : _GEN_910; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_975 = 3'h2 == encoders_1_io_output ? proc_2_io_next_header_13 : _GEN_911; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_976 = 3'h2 == encoders_1_io_output ? proc_2_io_next_header_14 : _GEN_912; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_977 = 3'h2 == encoders_1_io_output ? proc_2_io_next_header_15 : _GEN_913; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_978 = 3'h2 == encoders_1_io_output ? proc_2_io_next_header_16 : _GEN_914; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_979 = 3'h2 == encoders_1_io_output ? proc_2_io_next_header_17 : _GEN_915; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_980 = 3'h2 == encoders_1_io_output ? proc_2_io_next_header_18 : _GEN_916; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_981 = 3'h2 == encoders_1_io_output ? proc_2_io_next_header_19 : _GEN_917; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_982 = 3'h2 == encoders_1_io_output ? proc_2_io_next_header_20 : _GEN_918; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_983 = 3'h2 == encoders_1_io_output ? proc_2_io_next_header_21 : _GEN_919; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_984 = 3'h2 == encoders_1_io_output ? proc_2_io_next_header_22 : _GEN_920; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_985 = 3'h2 == encoders_1_io_output ? proc_2_io_next_header_23 : _GEN_921; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_986 = 3'h2 == encoders_1_io_output ? proc_2_io_next_header_24 : _GEN_922; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_987 = 3'h2 == encoders_1_io_output ? proc_2_io_next_header_25 : _GEN_923; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_988 = 3'h2 == encoders_1_io_output ? proc_2_io_next_header_26 : _GEN_924; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_989 = 3'h2 == encoders_1_io_output ? proc_2_io_next_header_27 : _GEN_925; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_990 = 3'h2 == encoders_1_io_output ? proc_2_io_next_header_28 : _GEN_926; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_991 = 3'h2 == encoders_1_io_output ? proc_2_io_next_header_29 : _GEN_927; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_992 = 3'h2 == encoders_1_io_output ? proc_2_io_next_header_30 : _GEN_928; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_993 = 3'h2 == encoders_1_io_output ? proc_2_io_next_header_31 : _GEN_929; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_994 = 3'h2 == encoders_1_io_output ? proc_2_io_next_header_32 : _GEN_930; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_995 = 3'h2 == encoders_1_io_output ? proc_2_io_next_header_33 : _GEN_931; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_996 = 3'h2 == encoders_1_io_output ? proc_2_io_next_header_34 : _GEN_932; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_997 = 3'h2 == encoders_1_io_output ? proc_2_io_next_header_35 : _GEN_933; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_998 = 3'h2 == encoders_1_io_output ? proc_2_io_next_header_36 : _GEN_934; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_999 = 3'h2 == encoders_1_io_output ? proc_2_io_next_header_37 : _GEN_935; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1000 = 3'h2 == encoders_1_io_output ? proc_2_io_next_header_38 : _GEN_936; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1001 = 3'h2 == encoders_1_io_output ? proc_2_io_next_header_39 : _GEN_937; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1002 = 3'h2 == encoders_1_io_output ? proc_2_io_next_header_40 : _GEN_938; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1003 = 3'h2 == encoders_1_io_output ? proc_2_io_next_header_41 : _GEN_939; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1004 = 3'h2 == encoders_1_io_output ? proc_2_io_next_header_42 : _GEN_940; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1005 = 3'h2 == encoders_1_io_output ? proc_2_io_next_header_43 : _GEN_941; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1006 = 3'h2 == encoders_1_io_output ? proc_2_io_next_header_44 : _GEN_942; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1007 = 3'h2 == encoders_1_io_output ? proc_2_io_next_header_45 : _GEN_943; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1008 = 3'h2 == encoders_1_io_output ? proc_2_io_next_header_46 : _GEN_944; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1009 = 3'h2 == encoders_1_io_output ? proc_2_io_next_header_47 : _GEN_945; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1010 = 3'h2 == encoders_1_io_output ? proc_2_io_next_header_48 : _GEN_946; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1011 = 3'h2 == encoders_1_io_output ? proc_2_io_next_header_49 : _GEN_947; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1012 = 3'h2 == encoders_1_io_output ? proc_2_io_next_header_50 : _GEN_948; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1013 = 3'h2 == encoders_1_io_output ? proc_2_io_next_header_51 : _GEN_949; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1014 = 3'h2 == encoders_1_io_output ? proc_2_io_next_header_52 : _GEN_950; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1015 = 3'h2 == encoders_1_io_output ? proc_2_io_next_header_53 : _GEN_951; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1016 = 3'h2 == encoders_1_io_output ? proc_2_io_next_header_54 : _GEN_952; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1017 = 3'h2 == encoders_1_io_output ? proc_2_io_next_header_55 : _GEN_953; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1018 = 3'h2 == encoders_1_io_output ? proc_2_io_next_header_56 : _GEN_954; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1019 = 3'h2 == encoders_1_io_output ? proc_2_io_next_header_57 : _GEN_955; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1020 = 3'h2 == encoders_1_io_output ? proc_2_io_next_header_58 : _GEN_956; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1021 = 3'h2 == encoders_1_io_output ? proc_2_io_next_header_59 : _GEN_957; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1022 = 3'h2 == encoders_1_io_output ? proc_2_io_next_header_60 : _GEN_958; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1023 = 3'h2 == encoders_1_io_output ? proc_2_io_next_header_61 : _GEN_959; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1024 = 3'h2 == encoders_1_io_output ? proc_2_io_next_header_62 : _GEN_960; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1025 = 3'h2 == encoders_1_io_output ? proc_2_io_next_header_63 : _GEN_961; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1026 = 3'h3 == encoders_1_io_output ? proc_3_io_next_header_0 : _GEN_962; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1027 = 3'h3 == encoders_1_io_output ? proc_3_io_next_header_1 : _GEN_963; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1028 = 3'h3 == encoders_1_io_output ? proc_3_io_next_header_2 : _GEN_964; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1029 = 3'h3 == encoders_1_io_output ? proc_3_io_next_header_3 : _GEN_965; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1030 = 3'h3 == encoders_1_io_output ? proc_3_io_next_header_4 : _GEN_966; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1031 = 3'h3 == encoders_1_io_output ? proc_3_io_next_header_5 : _GEN_967; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1032 = 3'h3 == encoders_1_io_output ? proc_3_io_next_header_6 : _GEN_968; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1033 = 3'h3 == encoders_1_io_output ? proc_3_io_next_header_7 : _GEN_969; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1034 = 3'h3 == encoders_1_io_output ? proc_3_io_next_header_8 : _GEN_970; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1035 = 3'h3 == encoders_1_io_output ? proc_3_io_next_header_9 : _GEN_971; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1036 = 3'h3 == encoders_1_io_output ? proc_3_io_next_header_10 : _GEN_972; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1037 = 3'h3 == encoders_1_io_output ? proc_3_io_next_header_11 : _GEN_973; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1038 = 3'h3 == encoders_1_io_output ? proc_3_io_next_header_12 : _GEN_974; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1039 = 3'h3 == encoders_1_io_output ? proc_3_io_next_header_13 : _GEN_975; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1040 = 3'h3 == encoders_1_io_output ? proc_3_io_next_header_14 : _GEN_976; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1041 = 3'h3 == encoders_1_io_output ? proc_3_io_next_header_15 : _GEN_977; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1042 = 3'h3 == encoders_1_io_output ? proc_3_io_next_header_16 : _GEN_978; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1043 = 3'h3 == encoders_1_io_output ? proc_3_io_next_header_17 : _GEN_979; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1044 = 3'h3 == encoders_1_io_output ? proc_3_io_next_header_18 : _GEN_980; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1045 = 3'h3 == encoders_1_io_output ? proc_3_io_next_header_19 : _GEN_981; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1046 = 3'h3 == encoders_1_io_output ? proc_3_io_next_header_20 : _GEN_982; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1047 = 3'h3 == encoders_1_io_output ? proc_3_io_next_header_21 : _GEN_983; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1048 = 3'h3 == encoders_1_io_output ? proc_3_io_next_header_22 : _GEN_984; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1049 = 3'h3 == encoders_1_io_output ? proc_3_io_next_header_23 : _GEN_985; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1050 = 3'h3 == encoders_1_io_output ? proc_3_io_next_header_24 : _GEN_986; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1051 = 3'h3 == encoders_1_io_output ? proc_3_io_next_header_25 : _GEN_987; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1052 = 3'h3 == encoders_1_io_output ? proc_3_io_next_header_26 : _GEN_988; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1053 = 3'h3 == encoders_1_io_output ? proc_3_io_next_header_27 : _GEN_989; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1054 = 3'h3 == encoders_1_io_output ? proc_3_io_next_header_28 : _GEN_990; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1055 = 3'h3 == encoders_1_io_output ? proc_3_io_next_header_29 : _GEN_991; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1056 = 3'h3 == encoders_1_io_output ? proc_3_io_next_header_30 : _GEN_992; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1057 = 3'h3 == encoders_1_io_output ? proc_3_io_next_header_31 : _GEN_993; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1058 = 3'h3 == encoders_1_io_output ? proc_3_io_next_header_32 : _GEN_994; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1059 = 3'h3 == encoders_1_io_output ? proc_3_io_next_header_33 : _GEN_995; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1060 = 3'h3 == encoders_1_io_output ? proc_3_io_next_header_34 : _GEN_996; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1061 = 3'h3 == encoders_1_io_output ? proc_3_io_next_header_35 : _GEN_997; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1062 = 3'h3 == encoders_1_io_output ? proc_3_io_next_header_36 : _GEN_998; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1063 = 3'h3 == encoders_1_io_output ? proc_3_io_next_header_37 : _GEN_999; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1064 = 3'h3 == encoders_1_io_output ? proc_3_io_next_header_38 : _GEN_1000; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1065 = 3'h3 == encoders_1_io_output ? proc_3_io_next_header_39 : _GEN_1001; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1066 = 3'h3 == encoders_1_io_output ? proc_3_io_next_header_40 : _GEN_1002; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1067 = 3'h3 == encoders_1_io_output ? proc_3_io_next_header_41 : _GEN_1003; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1068 = 3'h3 == encoders_1_io_output ? proc_3_io_next_header_42 : _GEN_1004; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1069 = 3'h3 == encoders_1_io_output ? proc_3_io_next_header_43 : _GEN_1005; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1070 = 3'h3 == encoders_1_io_output ? proc_3_io_next_header_44 : _GEN_1006; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1071 = 3'h3 == encoders_1_io_output ? proc_3_io_next_header_45 : _GEN_1007; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1072 = 3'h3 == encoders_1_io_output ? proc_3_io_next_header_46 : _GEN_1008; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1073 = 3'h3 == encoders_1_io_output ? proc_3_io_next_header_47 : _GEN_1009; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1074 = 3'h3 == encoders_1_io_output ? proc_3_io_next_header_48 : _GEN_1010; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1075 = 3'h3 == encoders_1_io_output ? proc_3_io_next_header_49 : _GEN_1011; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1076 = 3'h3 == encoders_1_io_output ? proc_3_io_next_header_50 : _GEN_1012; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1077 = 3'h3 == encoders_1_io_output ? proc_3_io_next_header_51 : _GEN_1013; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1078 = 3'h3 == encoders_1_io_output ? proc_3_io_next_header_52 : _GEN_1014; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1079 = 3'h3 == encoders_1_io_output ? proc_3_io_next_header_53 : _GEN_1015; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1080 = 3'h3 == encoders_1_io_output ? proc_3_io_next_header_54 : _GEN_1016; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1081 = 3'h3 == encoders_1_io_output ? proc_3_io_next_header_55 : _GEN_1017; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1082 = 3'h3 == encoders_1_io_output ? proc_3_io_next_header_56 : _GEN_1018; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1083 = 3'h3 == encoders_1_io_output ? proc_3_io_next_header_57 : _GEN_1019; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1084 = 3'h3 == encoders_1_io_output ? proc_3_io_next_header_58 : _GEN_1020; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1085 = 3'h3 == encoders_1_io_output ? proc_3_io_next_header_59 : _GEN_1021; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1086 = 3'h3 == encoders_1_io_output ? proc_3_io_next_header_60 : _GEN_1022; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1087 = 3'h3 == encoders_1_io_output ? proc_3_io_next_header_61 : _GEN_1023; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1088 = 3'h3 == encoders_1_io_output ? proc_3_io_next_header_62 : _GEN_1024; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1089 = 3'h3 == encoders_1_io_output ? proc_3_io_next_header_63 : _GEN_1025; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1090 = 3'h4 == encoders_1_io_output ? proc_4_io_next_header_0 : _GEN_1026; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1091 = 3'h4 == encoders_1_io_output ? proc_4_io_next_header_1 : _GEN_1027; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1092 = 3'h4 == encoders_1_io_output ? proc_4_io_next_header_2 : _GEN_1028; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1093 = 3'h4 == encoders_1_io_output ? proc_4_io_next_header_3 : _GEN_1029; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1094 = 3'h4 == encoders_1_io_output ? proc_4_io_next_header_4 : _GEN_1030; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1095 = 3'h4 == encoders_1_io_output ? proc_4_io_next_header_5 : _GEN_1031; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1096 = 3'h4 == encoders_1_io_output ? proc_4_io_next_header_6 : _GEN_1032; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1097 = 3'h4 == encoders_1_io_output ? proc_4_io_next_header_7 : _GEN_1033; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1098 = 3'h4 == encoders_1_io_output ? proc_4_io_next_header_8 : _GEN_1034; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1099 = 3'h4 == encoders_1_io_output ? proc_4_io_next_header_9 : _GEN_1035; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1100 = 3'h4 == encoders_1_io_output ? proc_4_io_next_header_10 : _GEN_1036; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1101 = 3'h4 == encoders_1_io_output ? proc_4_io_next_header_11 : _GEN_1037; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1102 = 3'h4 == encoders_1_io_output ? proc_4_io_next_header_12 : _GEN_1038; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1103 = 3'h4 == encoders_1_io_output ? proc_4_io_next_header_13 : _GEN_1039; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1104 = 3'h4 == encoders_1_io_output ? proc_4_io_next_header_14 : _GEN_1040; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1105 = 3'h4 == encoders_1_io_output ? proc_4_io_next_header_15 : _GEN_1041; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1106 = 3'h4 == encoders_1_io_output ? proc_4_io_next_header_16 : _GEN_1042; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1107 = 3'h4 == encoders_1_io_output ? proc_4_io_next_header_17 : _GEN_1043; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1108 = 3'h4 == encoders_1_io_output ? proc_4_io_next_header_18 : _GEN_1044; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1109 = 3'h4 == encoders_1_io_output ? proc_4_io_next_header_19 : _GEN_1045; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1110 = 3'h4 == encoders_1_io_output ? proc_4_io_next_header_20 : _GEN_1046; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1111 = 3'h4 == encoders_1_io_output ? proc_4_io_next_header_21 : _GEN_1047; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1112 = 3'h4 == encoders_1_io_output ? proc_4_io_next_header_22 : _GEN_1048; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1113 = 3'h4 == encoders_1_io_output ? proc_4_io_next_header_23 : _GEN_1049; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1114 = 3'h4 == encoders_1_io_output ? proc_4_io_next_header_24 : _GEN_1050; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1115 = 3'h4 == encoders_1_io_output ? proc_4_io_next_header_25 : _GEN_1051; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1116 = 3'h4 == encoders_1_io_output ? proc_4_io_next_header_26 : _GEN_1052; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1117 = 3'h4 == encoders_1_io_output ? proc_4_io_next_header_27 : _GEN_1053; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1118 = 3'h4 == encoders_1_io_output ? proc_4_io_next_header_28 : _GEN_1054; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1119 = 3'h4 == encoders_1_io_output ? proc_4_io_next_header_29 : _GEN_1055; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1120 = 3'h4 == encoders_1_io_output ? proc_4_io_next_header_30 : _GEN_1056; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1121 = 3'h4 == encoders_1_io_output ? proc_4_io_next_header_31 : _GEN_1057; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1122 = 3'h4 == encoders_1_io_output ? proc_4_io_next_header_32 : _GEN_1058; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1123 = 3'h4 == encoders_1_io_output ? proc_4_io_next_header_33 : _GEN_1059; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1124 = 3'h4 == encoders_1_io_output ? proc_4_io_next_header_34 : _GEN_1060; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1125 = 3'h4 == encoders_1_io_output ? proc_4_io_next_header_35 : _GEN_1061; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1126 = 3'h4 == encoders_1_io_output ? proc_4_io_next_header_36 : _GEN_1062; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1127 = 3'h4 == encoders_1_io_output ? proc_4_io_next_header_37 : _GEN_1063; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1128 = 3'h4 == encoders_1_io_output ? proc_4_io_next_header_38 : _GEN_1064; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1129 = 3'h4 == encoders_1_io_output ? proc_4_io_next_header_39 : _GEN_1065; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1130 = 3'h4 == encoders_1_io_output ? proc_4_io_next_header_40 : _GEN_1066; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1131 = 3'h4 == encoders_1_io_output ? proc_4_io_next_header_41 : _GEN_1067; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1132 = 3'h4 == encoders_1_io_output ? proc_4_io_next_header_42 : _GEN_1068; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1133 = 3'h4 == encoders_1_io_output ? proc_4_io_next_header_43 : _GEN_1069; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1134 = 3'h4 == encoders_1_io_output ? proc_4_io_next_header_44 : _GEN_1070; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1135 = 3'h4 == encoders_1_io_output ? proc_4_io_next_header_45 : _GEN_1071; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1136 = 3'h4 == encoders_1_io_output ? proc_4_io_next_header_46 : _GEN_1072; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1137 = 3'h4 == encoders_1_io_output ? proc_4_io_next_header_47 : _GEN_1073; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1138 = 3'h4 == encoders_1_io_output ? proc_4_io_next_header_48 : _GEN_1074; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1139 = 3'h4 == encoders_1_io_output ? proc_4_io_next_header_49 : _GEN_1075; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1140 = 3'h4 == encoders_1_io_output ? proc_4_io_next_header_50 : _GEN_1076; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1141 = 3'h4 == encoders_1_io_output ? proc_4_io_next_header_51 : _GEN_1077; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1142 = 3'h4 == encoders_1_io_output ? proc_4_io_next_header_52 : _GEN_1078; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1143 = 3'h4 == encoders_1_io_output ? proc_4_io_next_header_53 : _GEN_1079; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1144 = 3'h4 == encoders_1_io_output ? proc_4_io_next_header_54 : _GEN_1080; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1145 = 3'h4 == encoders_1_io_output ? proc_4_io_next_header_55 : _GEN_1081; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1146 = 3'h4 == encoders_1_io_output ? proc_4_io_next_header_56 : _GEN_1082; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1147 = 3'h4 == encoders_1_io_output ? proc_4_io_next_header_57 : _GEN_1083; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1148 = 3'h4 == encoders_1_io_output ? proc_4_io_next_header_58 : _GEN_1084; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1149 = 3'h4 == encoders_1_io_output ? proc_4_io_next_header_59 : _GEN_1085; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1150 = 3'h4 == encoders_1_io_output ? proc_4_io_next_header_60 : _GEN_1086; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1151 = 3'h4 == encoders_1_io_output ? proc_4_io_next_header_61 : _GEN_1087; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1152 = 3'h4 == encoders_1_io_output ? proc_4_io_next_header_62 : _GEN_1088; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1153 = 3'h4 == encoders_1_io_output ? proc_4_io_next_header_63 : _GEN_1089; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1154 = 3'h5 == encoders_1_io_output ? proc_5_io_next_header_0 : _GEN_1090; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1155 = 3'h5 == encoders_1_io_output ? proc_5_io_next_header_1 : _GEN_1091; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1156 = 3'h5 == encoders_1_io_output ? proc_5_io_next_header_2 : _GEN_1092; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1157 = 3'h5 == encoders_1_io_output ? proc_5_io_next_header_3 : _GEN_1093; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1158 = 3'h5 == encoders_1_io_output ? proc_5_io_next_header_4 : _GEN_1094; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1159 = 3'h5 == encoders_1_io_output ? proc_5_io_next_header_5 : _GEN_1095; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1160 = 3'h5 == encoders_1_io_output ? proc_5_io_next_header_6 : _GEN_1096; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1161 = 3'h5 == encoders_1_io_output ? proc_5_io_next_header_7 : _GEN_1097; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1162 = 3'h5 == encoders_1_io_output ? proc_5_io_next_header_8 : _GEN_1098; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1163 = 3'h5 == encoders_1_io_output ? proc_5_io_next_header_9 : _GEN_1099; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1164 = 3'h5 == encoders_1_io_output ? proc_5_io_next_header_10 : _GEN_1100; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1165 = 3'h5 == encoders_1_io_output ? proc_5_io_next_header_11 : _GEN_1101; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1166 = 3'h5 == encoders_1_io_output ? proc_5_io_next_header_12 : _GEN_1102; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1167 = 3'h5 == encoders_1_io_output ? proc_5_io_next_header_13 : _GEN_1103; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1168 = 3'h5 == encoders_1_io_output ? proc_5_io_next_header_14 : _GEN_1104; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1169 = 3'h5 == encoders_1_io_output ? proc_5_io_next_header_15 : _GEN_1105; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1170 = 3'h5 == encoders_1_io_output ? proc_5_io_next_header_16 : _GEN_1106; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1171 = 3'h5 == encoders_1_io_output ? proc_5_io_next_header_17 : _GEN_1107; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1172 = 3'h5 == encoders_1_io_output ? proc_5_io_next_header_18 : _GEN_1108; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1173 = 3'h5 == encoders_1_io_output ? proc_5_io_next_header_19 : _GEN_1109; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1174 = 3'h5 == encoders_1_io_output ? proc_5_io_next_header_20 : _GEN_1110; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1175 = 3'h5 == encoders_1_io_output ? proc_5_io_next_header_21 : _GEN_1111; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1176 = 3'h5 == encoders_1_io_output ? proc_5_io_next_header_22 : _GEN_1112; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1177 = 3'h5 == encoders_1_io_output ? proc_5_io_next_header_23 : _GEN_1113; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1178 = 3'h5 == encoders_1_io_output ? proc_5_io_next_header_24 : _GEN_1114; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1179 = 3'h5 == encoders_1_io_output ? proc_5_io_next_header_25 : _GEN_1115; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1180 = 3'h5 == encoders_1_io_output ? proc_5_io_next_header_26 : _GEN_1116; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1181 = 3'h5 == encoders_1_io_output ? proc_5_io_next_header_27 : _GEN_1117; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1182 = 3'h5 == encoders_1_io_output ? proc_5_io_next_header_28 : _GEN_1118; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1183 = 3'h5 == encoders_1_io_output ? proc_5_io_next_header_29 : _GEN_1119; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1184 = 3'h5 == encoders_1_io_output ? proc_5_io_next_header_30 : _GEN_1120; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1185 = 3'h5 == encoders_1_io_output ? proc_5_io_next_header_31 : _GEN_1121; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1186 = 3'h5 == encoders_1_io_output ? proc_5_io_next_header_32 : _GEN_1122; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1187 = 3'h5 == encoders_1_io_output ? proc_5_io_next_header_33 : _GEN_1123; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1188 = 3'h5 == encoders_1_io_output ? proc_5_io_next_header_34 : _GEN_1124; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1189 = 3'h5 == encoders_1_io_output ? proc_5_io_next_header_35 : _GEN_1125; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1190 = 3'h5 == encoders_1_io_output ? proc_5_io_next_header_36 : _GEN_1126; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1191 = 3'h5 == encoders_1_io_output ? proc_5_io_next_header_37 : _GEN_1127; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1192 = 3'h5 == encoders_1_io_output ? proc_5_io_next_header_38 : _GEN_1128; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1193 = 3'h5 == encoders_1_io_output ? proc_5_io_next_header_39 : _GEN_1129; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1194 = 3'h5 == encoders_1_io_output ? proc_5_io_next_header_40 : _GEN_1130; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1195 = 3'h5 == encoders_1_io_output ? proc_5_io_next_header_41 : _GEN_1131; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1196 = 3'h5 == encoders_1_io_output ? proc_5_io_next_header_42 : _GEN_1132; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1197 = 3'h5 == encoders_1_io_output ? proc_5_io_next_header_43 : _GEN_1133; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1198 = 3'h5 == encoders_1_io_output ? proc_5_io_next_header_44 : _GEN_1134; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1199 = 3'h5 == encoders_1_io_output ? proc_5_io_next_header_45 : _GEN_1135; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1200 = 3'h5 == encoders_1_io_output ? proc_5_io_next_header_46 : _GEN_1136; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1201 = 3'h5 == encoders_1_io_output ? proc_5_io_next_header_47 : _GEN_1137; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1202 = 3'h5 == encoders_1_io_output ? proc_5_io_next_header_48 : _GEN_1138; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1203 = 3'h5 == encoders_1_io_output ? proc_5_io_next_header_49 : _GEN_1139; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1204 = 3'h5 == encoders_1_io_output ? proc_5_io_next_header_50 : _GEN_1140; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1205 = 3'h5 == encoders_1_io_output ? proc_5_io_next_header_51 : _GEN_1141; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1206 = 3'h5 == encoders_1_io_output ? proc_5_io_next_header_52 : _GEN_1142; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1207 = 3'h5 == encoders_1_io_output ? proc_5_io_next_header_53 : _GEN_1143; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1208 = 3'h5 == encoders_1_io_output ? proc_5_io_next_header_54 : _GEN_1144; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1209 = 3'h5 == encoders_1_io_output ? proc_5_io_next_header_55 : _GEN_1145; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1210 = 3'h5 == encoders_1_io_output ? proc_5_io_next_header_56 : _GEN_1146; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1211 = 3'h5 == encoders_1_io_output ? proc_5_io_next_header_57 : _GEN_1147; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1212 = 3'h5 == encoders_1_io_output ? proc_5_io_next_header_58 : _GEN_1148; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1213 = 3'h5 == encoders_1_io_output ? proc_5_io_next_header_59 : _GEN_1149; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1214 = 3'h5 == encoders_1_io_output ? proc_5_io_next_header_60 : _GEN_1150; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1215 = 3'h5 == encoders_1_io_output ? proc_5_io_next_header_61 : _GEN_1151; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1216 = 3'h5 == encoders_1_io_output ? proc_5_io_next_header_62 : _GEN_1152; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1217 = 3'h5 == encoders_1_io_output ? proc_5_io_next_header_63 : _GEN_1153; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1218 = 3'h6 == encoders_1_io_output ? proc_6_io_next_header_0 : _GEN_1154; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1219 = 3'h6 == encoders_1_io_output ? proc_6_io_next_header_1 : _GEN_1155; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1220 = 3'h6 == encoders_1_io_output ? proc_6_io_next_header_2 : _GEN_1156; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1221 = 3'h6 == encoders_1_io_output ? proc_6_io_next_header_3 : _GEN_1157; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1222 = 3'h6 == encoders_1_io_output ? proc_6_io_next_header_4 : _GEN_1158; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1223 = 3'h6 == encoders_1_io_output ? proc_6_io_next_header_5 : _GEN_1159; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1224 = 3'h6 == encoders_1_io_output ? proc_6_io_next_header_6 : _GEN_1160; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1225 = 3'h6 == encoders_1_io_output ? proc_6_io_next_header_7 : _GEN_1161; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1226 = 3'h6 == encoders_1_io_output ? proc_6_io_next_header_8 : _GEN_1162; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1227 = 3'h6 == encoders_1_io_output ? proc_6_io_next_header_9 : _GEN_1163; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1228 = 3'h6 == encoders_1_io_output ? proc_6_io_next_header_10 : _GEN_1164; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1229 = 3'h6 == encoders_1_io_output ? proc_6_io_next_header_11 : _GEN_1165; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1230 = 3'h6 == encoders_1_io_output ? proc_6_io_next_header_12 : _GEN_1166; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1231 = 3'h6 == encoders_1_io_output ? proc_6_io_next_header_13 : _GEN_1167; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1232 = 3'h6 == encoders_1_io_output ? proc_6_io_next_header_14 : _GEN_1168; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1233 = 3'h6 == encoders_1_io_output ? proc_6_io_next_header_15 : _GEN_1169; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1234 = 3'h6 == encoders_1_io_output ? proc_6_io_next_header_16 : _GEN_1170; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1235 = 3'h6 == encoders_1_io_output ? proc_6_io_next_header_17 : _GEN_1171; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1236 = 3'h6 == encoders_1_io_output ? proc_6_io_next_header_18 : _GEN_1172; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1237 = 3'h6 == encoders_1_io_output ? proc_6_io_next_header_19 : _GEN_1173; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1238 = 3'h6 == encoders_1_io_output ? proc_6_io_next_header_20 : _GEN_1174; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1239 = 3'h6 == encoders_1_io_output ? proc_6_io_next_header_21 : _GEN_1175; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1240 = 3'h6 == encoders_1_io_output ? proc_6_io_next_header_22 : _GEN_1176; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1241 = 3'h6 == encoders_1_io_output ? proc_6_io_next_header_23 : _GEN_1177; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1242 = 3'h6 == encoders_1_io_output ? proc_6_io_next_header_24 : _GEN_1178; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1243 = 3'h6 == encoders_1_io_output ? proc_6_io_next_header_25 : _GEN_1179; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1244 = 3'h6 == encoders_1_io_output ? proc_6_io_next_header_26 : _GEN_1180; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1245 = 3'h6 == encoders_1_io_output ? proc_6_io_next_header_27 : _GEN_1181; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1246 = 3'h6 == encoders_1_io_output ? proc_6_io_next_header_28 : _GEN_1182; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1247 = 3'h6 == encoders_1_io_output ? proc_6_io_next_header_29 : _GEN_1183; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1248 = 3'h6 == encoders_1_io_output ? proc_6_io_next_header_30 : _GEN_1184; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1249 = 3'h6 == encoders_1_io_output ? proc_6_io_next_header_31 : _GEN_1185; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1250 = 3'h6 == encoders_1_io_output ? proc_6_io_next_header_32 : _GEN_1186; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1251 = 3'h6 == encoders_1_io_output ? proc_6_io_next_header_33 : _GEN_1187; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1252 = 3'h6 == encoders_1_io_output ? proc_6_io_next_header_34 : _GEN_1188; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1253 = 3'h6 == encoders_1_io_output ? proc_6_io_next_header_35 : _GEN_1189; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1254 = 3'h6 == encoders_1_io_output ? proc_6_io_next_header_36 : _GEN_1190; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1255 = 3'h6 == encoders_1_io_output ? proc_6_io_next_header_37 : _GEN_1191; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1256 = 3'h6 == encoders_1_io_output ? proc_6_io_next_header_38 : _GEN_1192; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1257 = 3'h6 == encoders_1_io_output ? proc_6_io_next_header_39 : _GEN_1193; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1258 = 3'h6 == encoders_1_io_output ? proc_6_io_next_header_40 : _GEN_1194; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1259 = 3'h6 == encoders_1_io_output ? proc_6_io_next_header_41 : _GEN_1195; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1260 = 3'h6 == encoders_1_io_output ? proc_6_io_next_header_42 : _GEN_1196; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1261 = 3'h6 == encoders_1_io_output ? proc_6_io_next_header_43 : _GEN_1197; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1262 = 3'h6 == encoders_1_io_output ? proc_6_io_next_header_44 : _GEN_1198; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1263 = 3'h6 == encoders_1_io_output ? proc_6_io_next_header_45 : _GEN_1199; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1264 = 3'h6 == encoders_1_io_output ? proc_6_io_next_header_46 : _GEN_1200; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1265 = 3'h6 == encoders_1_io_output ? proc_6_io_next_header_47 : _GEN_1201; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1266 = 3'h6 == encoders_1_io_output ? proc_6_io_next_header_48 : _GEN_1202; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1267 = 3'h6 == encoders_1_io_output ? proc_6_io_next_header_49 : _GEN_1203; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1268 = 3'h6 == encoders_1_io_output ? proc_6_io_next_header_50 : _GEN_1204; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1269 = 3'h6 == encoders_1_io_output ? proc_6_io_next_header_51 : _GEN_1205; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1270 = 3'h6 == encoders_1_io_output ? proc_6_io_next_header_52 : _GEN_1206; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1271 = 3'h6 == encoders_1_io_output ? proc_6_io_next_header_53 : _GEN_1207; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1272 = 3'h6 == encoders_1_io_output ? proc_6_io_next_header_54 : _GEN_1208; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1273 = 3'h6 == encoders_1_io_output ? proc_6_io_next_header_55 : _GEN_1209; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1274 = 3'h6 == encoders_1_io_output ? proc_6_io_next_header_56 : _GEN_1210; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1275 = 3'h6 == encoders_1_io_output ? proc_6_io_next_header_57 : _GEN_1211; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1276 = 3'h6 == encoders_1_io_output ? proc_6_io_next_header_58 : _GEN_1212; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1277 = 3'h6 == encoders_1_io_output ? proc_6_io_next_header_59 : _GEN_1213; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1278 = 3'h6 == encoders_1_io_output ? proc_6_io_next_header_60 : _GEN_1214; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1279 = 3'h6 == encoders_1_io_output ? proc_6_io_next_header_61 : _GEN_1215; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1280 = 3'h6 == encoders_1_io_output ? proc_6_io_next_header_62 : _GEN_1216; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1281 = 3'h6 == encoders_1_io_output ? proc_6_io_next_header_63 : _GEN_1217; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1282 = 3'h7 == encoders_1_io_output ? proc_7_io_next_header_0 : _GEN_1218; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1283 = 3'h7 == encoders_1_io_output ? proc_7_io_next_header_1 : _GEN_1219; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1284 = 3'h7 == encoders_1_io_output ? proc_7_io_next_header_2 : _GEN_1220; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1285 = 3'h7 == encoders_1_io_output ? proc_7_io_next_header_3 : _GEN_1221; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1286 = 3'h7 == encoders_1_io_output ? proc_7_io_next_header_4 : _GEN_1222; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1287 = 3'h7 == encoders_1_io_output ? proc_7_io_next_header_5 : _GEN_1223; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1288 = 3'h7 == encoders_1_io_output ? proc_7_io_next_header_6 : _GEN_1224; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1289 = 3'h7 == encoders_1_io_output ? proc_7_io_next_header_7 : _GEN_1225; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1290 = 3'h7 == encoders_1_io_output ? proc_7_io_next_header_8 : _GEN_1226; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1291 = 3'h7 == encoders_1_io_output ? proc_7_io_next_header_9 : _GEN_1227; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1292 = 3'h7 == encoders_1_io_output ? proc_7_io_next_header_10 : _GEN_1228; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1293 = 3'h7 == encoders_1_io_output ? proc_7_io_next_header_11 : _GEN_1229; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1294 = 3'h7 == encoders_1_io_output ? proc_7_io_next_header_12 : _GEN_1230; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1295 = 3'h7 == encoders_1_io_output ? proc_7_io_next_header_13 : _GEN_1231; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1296 = 3'h7 == encoders_1_io_output ? proc_7_io_next_header_14 : _GEN_1232; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1297 = 3'h7 == encoders_1_io_output ? proc_7_io_next_header_15 : _GEN_1233; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1298 = 3'h7 == encoders_1_io_output ? proc_7_io_next_header_16 : _GEN_1234; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1299 = 3'h7 == encoders_1_io_output ? proc_7_io_next_header_17 : _GEN_1235; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1300 = 3'h7 == encoders_1_io_output ? proc_7_io_next_header_18 : _GEN_1236; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1301 = 3'h7 == encoders_1_io_output ? proc_7_io_next_header_19 : _GEN_1237; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1302 = 3'h7 == encoders_1_io_output ? proc_7_io_next_header_20 : _GEN_1238; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1303 = 3'h7 == encoders_1_io_output ? proc_7_io_next_header_21 : _GEN_1239; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1304 = 3'h7 == encoders_1_io_output ? proc_7_io_next_header_22 : _GEN_1240; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1305 = 3'h7 == encoders_1_io_output ? proc_7_io_next_header_23 : _GEN_1241; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1306 = 3'h7 == encoders_1_io_output ? proc_7_io_next_header_24 : _GEN_1242; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1307 = 3'h7 == encoders_1_io_output ? proc_7_io_next_header_25 : _GEN_1243; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1308 = 3'h7 == encoders_1_io_output ? proc_7_io_next_header_26 : _GEN_1244; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1309 = 3'h7 == encoders_1_io_output ? proc_7_io_next_header_27 : _GEN_1245; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1310 = 3'h7 == encoders_1_io_output ? proc_7_io_next_header_28 : _GEN_1246; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1311 = 3'h7 == encoders_1_io_output ? proc_7_io_next_header_29 : _GEN_1247; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1312 = 3'h7 == encoders_1_io_output ? proc_7_io_next_header_30 : _GEN_1248; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1313 = 3'h7 == encoders_1_io_output ? proc_7_io_next_header_31 : _GEN_1249; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1314 = 3'h7 == encoders_1_io_output ? proc_7_io_next_header_32 : _GEN_1250; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1315 = 3'h7 == encoders_1_io_output ? proc_7_io_next_header_33 : _GEN_1251; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1316 = 3'h7 == encoders_1_io_output ? proc_7_io_next_header_34 : _GEN_1252; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1317 = 3'h7 == encoders_1_io_output ? proc_7_io_next_header_35 : _GEN_1253; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1318 = 3'h7 == encoders_1_io_output ? proc_7_io_next_header_36 : _GEN_1254; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1319 = 3'h7 == encoders_1_io_output ? proc_7_io_next_header_37 : _GEN_1255; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1320 = 3'h7 == encoders_1_io_output ? proc_7_io_next_header_38 : _GEN_1256; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1321 = 3'h7 == encoders_1_io_output ? proc_7_io_next_header_39 : _GEN_1257; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1322 = 3'h7 == encoders_1_io_output ? proc_7_io_next_header_40 : _GEN_1258; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1323 = 3'h7 == encoders_1_io_output ? proc_7_io_next_header_41 : _GEN_1259; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1324 = 3'h7 == encoders_1_io_output ? proc_7_io_next_header_42 : _GEN_1260; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1325 = 3'h7 == encoders_1_io_output ? proc_7_io_next_header_43 : _GEN_1261; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1326 = 3'h7 == encoders_1_io_output ? proc_7_io_next_header_44 : _GEN_1262; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1327 = 3'h7 == encoders_1_io_output ? proc_7_io_next_header_45 : _GEN_1263; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1328 = 3'h7 == encoders_1_io_output ? proc_7_io_next_header_46 : _GEN_1264; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1329 = 3'h7 == encoders_1_io_output ? proc_7_io_next_header_47 : _GEN_1265; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1330 = 3'h7 == encoders_1_io_output ? proc_7_io_next_header_48 : _GEN_1266; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1331 = 3'h7 == encoders_1_io_output ? proc_7_io_next_header_49 : _GEN_1267; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1332 = 3'h7 == encoders_1_io_output ? proc_7_io_next_header_50 : _GEN_1268; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1333 = 3'h7 == encoders_1_io_output ? proc_7_io_next_header_51 : _GEN_1269; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1334 = 3'h7 == encoders_1_io_output ? proc_7_io_next_header_52 : _GEN_1270; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1335 = 3'h7 == encoders_1_io_output ? proc_7_io_next_header_53 : _GEN_1271; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1336 = 3'h7 == encoders_1_io_output ? proc_7_io_next_header_54 : _GEN_1272; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1337 = 3'h7 == encoders_1_io_output ? proc_7_io_next_header_55 : _GEN_1273; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1338 = 3'h7 == encoders_1_io_output ? proc_7_io_next_header_56 : _GEN_1274; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1339 = 3'h7 == encoders_1_io_output ? proc_7_io_next_header_57 : _GEN_1275; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1340 = 3'h7 == encoders_1_io_output ? proc_7_io_next_header_58 : _GEN_1276; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1341 = 3'h7 == encoders_1_io_output ? proc_7_io_next_header_59 : _GEN_1277; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1342 = 3'h7 == encoders_1_io_output ? proc_7_io_next_header_60 : _GEN_1278; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1343 = 3'h7 == encoders_1_io_output ? proc_7_io_next_header_61 : _GEN_1279; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1344 = 3'h7 == encoders_1_io_output ? proc_7_io_next_header_62 : _GEN_1280; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1345 = 3'h7 == encoders_1_io_output ? proc_7_io_next_header_63 : _GEN_1281; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1411 = 3'h0 == encoders_2_io_output ? proc_0_io_next_header_0 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1412 = 3'h0 == encoders_2_io_output ? proc_0_io_next_header_1 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1413 = 3'h0 == encoders_2_io_output ? proc_0_io_next_header_2 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1414 = 3'h0 == encoders_2_io_output ? proc_0_io_next_header_3 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1415 = 3'h0 == encoders_2_io_output ? proc_0_io_next_header_4 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1416 = 3'h0 == encoders_2_io_output ? proc_0_io_next_header_5 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1417 = 3'h0 == encoders_2_io_output ? proc_0_io_next_header_6 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1418 = 3'h0 == encoders_2_io_output ? proc_0_io_next_header_7 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1419 = 3'h0 == encoders_2_io_output ? proc_0_io_next_header_8 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1420 = 3'h0 == encoders_2_io_output ? proc_0_io_next_header_9 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1421 = 3'h0 == encoders_2_io_output ? proc_0_io_next_header_10 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1422 = 3'h0 == encoders_2_io_output ? proc_0_io_next_header_11 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1423 = 3'h0 == encoders_2_io_output ? proc_0_io_next_header_12 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1424 = 3'h0 == encoders_2_io_output ? proc_0_io_next_header_13 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1425 = 3'h0 == encoders_2_io_output ? proc_0_io_next_header_14 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1426 = 3'h0 == encoders_2_io_output ? proc_0_io_next_header_15 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1427 = 3'h0 == encoders_2_io_output ? proc_0_io_next_header_16 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1428 = 3'h0 == encoders_2_io_output ? proc_0_io_next_header_17 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1429 = 3'h0 == encoders_2_io_output ? proc_0_io_next_header_18 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1430 = 3'h0 == encoders_2_io_output ? proc_0_io_next_header_19 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1431 = 3'h0 == encoders_2_io_output ? proc_0_io_next_header_20 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1432 = 3'h0 == encoders_2_io_output ? proc_0_io_next_header_21 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1433 = 3'h0 == encoders_2_io_output ? proc_0_io_next_header_22 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1434 = 3'h0 == encoders_2_io_output ? proc_0_io_next_header_23 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1435 = 3'h0 == encoders_2_io_output ? proc_0_io_next_header_24 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1436 = 3'h0 == encoders_2_io_output ? proc_0_io_next_header_25 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1437 = 3'h0 == encoders_2_io_output ? proc_0_io_next_header_26 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1438 = 3'h0 == encoders_2_io_output ? proc_0_io_next_header_27 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1439 = 3'h0 == encoders_2_io_output ? proc_0_io_next_header_28 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1440 = 3'h0 == encoders_2_io_output ? proc_0_io_next_header_29 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1441 = 3'h0 == encoders_2_io_output ? proc_0_io_next_header_30 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1442 = 3'h0 == encoders_2_io_output ? proc_0_io_next_header_31 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1443 = 3'h0 == encoders_2_io_output ? proc_0_io_next_header_32 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1444 = 3'h0 == encoders_2_io_output ? proc_0_io_next_header_33 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1445 = 3'h0 == encoders_2_io_output ? proc_0_io_next_header_34 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1446 = 3'h0 == encoders_2_io_output ? proc_0_io_next_header_35 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1447 = 3'h0 == encoders_2_io_output ? proc_0_io_next_header_36 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1448 = 3'h0 == encoders_2_io_output ? proc_0_io_next_header_37 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1449 = 3'h0 == encoders_2_io_output ? proc_0_io_next_header_38 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1450 = 3'h0 == encoders_2_io_output ? proc_0_io_next_header_39 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1451 = 3'h0 == encoders_2_io_output ? proc_0_io_next_header_40 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1452 = 3'h0 == encoders_2_io_output ? proc_0_io_next_header_41 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1453 = 3'h0 == encoders_2_io_output ? proc_0_io_next_header_42 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1454 = 3'h0 == encoders_2_io_output ? proc_0_io_next_header_43 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1455 = 3'h0 == encoders_2_io_output ? proc_0_io_next_header_44 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1456 = 3'h0 == encoders_2_io_output ? proc_0_io_next_header_45 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1457 = 3'h0 == encoders_2_io_output ? proc_0_io_next_header_46 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1458 = 3'h0 == encoders_2_io_output ? proc_0_io_next_header_47 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1459 = 3'h0 == encoders_2_io_output ? proc_0_io_next_header_48 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1460 = 3'h0 == encoders_2_io_output ? proc_0_io_next_header_49 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1461 = 3'h0 == encoders_2_io_output ? proc_0_io_next_header_50 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1462 = 3'h0 == encoders_2_io_output ? proc_0_io_next_header_51 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1463 = 3'h0 == encoders_2_io_output ? proc_0_io_next_header_52 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1464 = 3'h0 == encoders_2_io_output ? proc_0_io_next_header_53 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1465 = 3'h0 == encoders_2_io_output ? proc_0_io_next_header_54 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1466 = 3'h0 == encoders_2_io_output ? proc_0_io_next_header_55 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1467 = 3'h0 == encoders_2_io_output ? proc_0_io_next_header_56 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1468 = 3'h0 == encoders_2_io_output ? proc_0_io_next_header_57 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1469 = 3'h0 == encoders_2_io_output ? proc_0_io_next_header_58 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1470 = 3'h0 == encoders_2_io_output ? proc_0_io_next_header_59 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1471 = 3'h0 == encoders_2_io_output ? proc_0_io_next_header_60 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1472 = 3'h0 == encoders_2_io_output ? proc_0_io_next_header_61 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1473 = 3'h0 == encoders_2_io_output ? proc_0_io_next_header_62 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1474 = 3'h0 == encoders_2_io_output ? proc_0_io_next_header_63 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1475 = 3'h1 == encoders_2_io_output ? proc_1_io_next_header_0 : _GEN_1411; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1476 = 3'h1 == encoders_2_io_output ? proc_1_io_next_header_1 : _GEN_1412; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1477 = 3'h1 == encoders_2_io_output ? proc_1_io_next_header_2 : _GEN_1413; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1478 = 3'h1 == encoders_2_io_output ? proc_1_io_next_header_3 : _GEN_1414; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1479 = 3'h1 == encoders_2_io_output ? proc_1_io_next_header_4 : _GEN_1415; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1480 = 3'h1 == encoders_2_io_output ? proc_1_io_next_header_5 : _GEN_1416; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1481 = 3'h1 == encoders_2_io_output ? proc_1_io_next_header_6 : _GEN_1417; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1482 = 3'h1 == encoders_2_io_output ? proc_1_io_next_header_7 : _GEN_1418; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1483 = 3'h1 == encoders_2_io_output ? proc_1_io_next_header_8 : _GEN_1419; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1484 = 3'h1 == encoders_2_io_output ? proc_1_io_next_header_9 : _GEN_1420; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1485 = 3'h1 == encoders_2_io_output ? proc_1_io_next_header_10 : _GEN_1421; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1486 = 3'h1 == encoders_2_io_output ? proc_1_io_next_header_11 : _GEN_1422; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1487 = 3'h1 == encoders_2_io_output ? proc_1_io_next_header_12 : _GEN_1423; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1488 = 3'h1 == encoders_2_io_output ? proc_1_io_next_header_13 : _GEN_1424; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1489 = 3'h1 == encoders_2_io_output ? proc_1_io_next_header_14 : _GEN_1425; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1490 = 3'h1 == encoders_2_io_output ? proc_1_io_next_header_15 : _GEN_1426; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1491 = 3'h1 == encoders_2_io_output ? proc_1_io_next_header_16 : _GEN_1427; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1492 = 3'h1 == encoders_2_io_output ? proc_1_io_next_header_17 : _GEN_1428; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1493 = 3'h1 == encoders_2_io_output ? proc_1_io_next_header_18 : _GEN_1429; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1494 = 3'h1 == encoders_2_io_output ? proc_1_io_next_header_19 : _GEN_1430; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1495 = 3'h1 == encoders_2_io_output ? proc_1_io_next_header_20 : _GEN_1431; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1496 = 3'h1 == encoders_2_io_output ? proc_1_io_next_header_21 : _GEN_1432; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1497 = 3'h1 == encoders_2_io_output ? proc_1_io_next_header_22 : _GEN_1433; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1498 = 3'h1 == encoders_2_io_output ? proc_1_io_next_header_23 : _GEN_1434; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1499 = 3'h1 == encoders_2_io_output ? proc_1_io_next_header_24 : _GEN_1435; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1500 = 3'h1 == encoders_2_io_output ? proc_1_io_next_header_25 : _GEN_1436; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1501 = 3'h1 == encoders_2_io_output ? proc_1_io_next_header_26 : _GEN_1437; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1502 = 3'h1 == encoders_2_io_output ? proc_1_io_next_header_27 : _GEN_1438; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1503 = 3'h1 == encoders_2_io_output ? proc_1_io_next_header_28 : _GEN_1439; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1504 = 3'h1 == encoders_2_io_output ? proc_1_io_next_header_29 : _GEN_1440; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1505 = 3'h1 == encoders_2_io_output ? proc_1_io_next_header_30 : _GEN_1441; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1506 = 3'h1 == encoders_2_io_output ? proc_1_io_next_header_31 : _GEN_1442; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1507 = 3'h1 == encoders_2_io_output ? proc_1_io_next_header_32 : _GEN_1443; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1508 = 3'h1 == encoders_2_io_output ? proc_1_io_next_header_33 : _GEN_1444; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1509 = 3'h1 == encoders_2_io_output ? proc_1_io_next_header_34 : _GEN_1445; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1510 = 3'h1 == encoders_2_io_output ? proc_1_io_next_header_35 : _GEN_1446; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1511 = 3'h1 == encoders_2_io_output ? proc_1_io_next_header_36 : _GEN_1447; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1512 = 3'h1 == encoders_2_io_output ? proc_1_io_next_header_37 : _GEN_1448; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1513 = 3'h1 == encoders_2_io_output ? proc_1_io_next_header_38 : _GEN_1449; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1514 = 3'h1 == encoders_2_io_output ? proc_1_io_next_header_39 : _GEN_1450; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1515 = 3'h1 == encoders_2_io_output ? proc_1_io_next_header_40 : _GEN_1451; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1516 = 3'h1 == encoders_2_io_output ? proc_1_io_next_header_41 : _GEN_1452; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1517 = 3'h1 == encoders_2_io_output ? proc_1_io_next_header_42 : _GEN_1453; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1518 = 3'h1 == encoders_2_io_output ? proc_1_io_next_header_43 : _GEN_1454; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1519 = 3'h1 == encoders_2_io_output ? proc_1_io_next_header_44 : _GEN_1455; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1520 = 3'h1 == encoders_2_io_output ? proc_1_io_next_header_45 : _GEN_1456; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1521 = 3'h1 == encoders_2_io_output ? proc_1_io_next_header_46 : _GEN_1457; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1522 = 3'h1 == encoders_2_io_output ? proc_1_io_next_header_47 : _GEN_1458; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1523 = 3'h1 == encoders_2_io_output ? proc_1_io_next_header_48 : _GEN_1459; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1524 = 3'h1 == encoders_2_io_output ? proc_1_io_next_header_49 : _GEN_1460; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1525 = 3'h1 == encoders_2_io_output ? proc_1_io_next_header_50 : _GEN_1461; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1526 = 3'h1 == encoders_2_io_output ? proc_1_io_next_header_51 : _GEN_1462; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1527 = 3'h1 == encoders_2_io_output ? proc_1_io_next_header_52 : _GEN_1463; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1528 = 3'h1 == encoders_2_io_output ? proc_1_io_next_header_53 : _GEN_1464; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1529 = 3'h1 == encoders_2_io_output ? proc_1_io_next_header_54 : _GEN_1465; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1530 = 3'h1 == encoders_2_io_output ? proc_1_io_next_header_55 : _GEN_1466; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1531 = 3'h1 == encoders_2_io_output ? proc_1_io_next_header_56 : _GEN_1467; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1532 = 3'h1 == encoders_2_io_output ? proc_1_io_next_header_57 : _GEN_1468; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1533 = 3'h1 == encoders_2_io_output ? proc_1_io_next_header_58 : _GEN_1469; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1534 = 3'h1 == encoders_2_io_output ? proc_1_io_next_header_59 : _GEN_1470; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1535 = 3'h1 == encoders_2_io_output ? proc_1_io_next_header_60 : _GEN_1471; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1536 = 3'h1 == encoders_2_io_output ? proc_1_io_next_header_61 : _GEN_1472; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1537 = 3'h1 == encoders_2_io_output ? proc_1_io_next_header_62 : _GEN_1473; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1538 = 3'h1 == encoders_2_io_output ? proc_1_io_next_header_63 : _GEN_1474; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1539 = 3'h2 == encoders_2_io_output ? proc_2_io_next_header_0 : _GEN_1475; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1540 = 3'h2 == encoders_2_io_output ? proc_2_io_next_header_1 : _GEN_1476; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1541 = 3'h2 == encoders_2_io_output ? proc_2_io_next_header_2 : _GEN_1477; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1542 = 3'h2 == encoders_2_io_output ? proc_2_io_next_header_3 : _GEN_1478; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1543 = 3'h2 == encoders_2_io_output ? proc_2_io_next_header_4 : _GEN_1479; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1544 = 3'h2 == encoders_2_io_output ? proc_2_io_next_header_5 : _GEN_1480; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1545 = 3'h2 == encoders_2_io_output ? proc_2_io_next_header_6 : _GEN_1481; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1546 = 3'h2 == encoders_2_io_output ? proc_2_io_next_header_7 : _GEN_1482; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1547 = 3'h2 == encoders_2_io_output ? proc_2_io_next_header_8 : _GEN_1483; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1548 = 3'h2 == encoders_2_io_output ? proc_2_io_next_header_9 : _GEN_1484; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1549 = 3'h2 == encoders_2_io_output ? proc_2_io_next_header_10 : _GEN_1485; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1550 = 3'h2 == encoders_2_io_output ? proc_2_io_next_header_11 : _GEN_1486; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1551 = 3'h2 == encoders_2_io_output ? proc_2_io_next_header_12 : _GEN_1487; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1552 = 3'h2 == encoders_2_io_output ? proc_2_io_next_header_13 : _GEN_1488; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1553 = 3'h2 == encoders_2_io_output ? proc_2_io_next_header_14 : _GEN_1489; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1554 = 3'h2 == encoders_2_io_output ? proc_2_io_next_header_15 : _GEN_1490; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1555 = 3'h2 == encoders_2_io_output ? proc_2_io_next_header_16 : _GEN_1491; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1556 = 3'h2 == encoders_2_io_output ? proc_2_io_next_header_17 : _GEN_1492; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1557 = 3'h2 == encoders_2_io_output ? proc_2_io_next_header_18 : _GEN_1493; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1558 = 3'h2 == encoders_2_io_output ? proc_2_io_next_header_19 : _GEN_1494; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1559 = 3'h2 == encoders_2_io_output ? proc_2_io_next_header_20 : _GEN_1495; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1560 = 3'h2 == encoders_2_io_output ? proc_2_io_next_header_21 : _GEN_1496; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1561 = 3'h2 == encoders_2_io_output ? proc_2_io_next_header_22 : _GEN_1497; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1562 = 3'h2 == encoders_2_io_output ? proc_2_io_next_header_23 : _GEN_1498; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1563 = 3'h2 == encoders_2_io_output ? proc_2_io_next_header_24 : _GEN_1499; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1564 = 3'h2 == encoders_2_io_output ? proc_2_io_next_header_25 : _GEN_1500; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1565 = 3'h2 == encoders_2_io_output ? proc_2_io_next_header_26 : _GEN_1501; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1566 = 3'h2 == encoders_2_io_output ? proc_2_io_next_header_27 : _GEN_1502; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1567 = 3'h2 == encoders_2_io_output ? proc_2_io_next_header_28 : _GEN_1503; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1568 = 3'h2 == encoders_2_io_output ? proc_2_io_next_header_29 : _GEN_1504; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1569 = 3'h2 == encoders_2_io_output ? proc_2_io_next_header_30 : _GEN_1505; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1570 = 3'h2 == encoders_2_io_output ? proc_2_io_next_header_31 : _GEN_1506; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1571 = 3'h2 == encoders_2_io_output ? proc_2_io_next_header_32 : _GEN_1507; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1572 = 3'h2 == encoders_2_io_output ? proc_2_io_next_header_33 : _GEN_1508; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1573 = 3'h2 == encoders_2_io_output ? proc_2_io_next_header_34 : _GEN_1509; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1574 = 3'h2 == encoders_2_io_output ? proc_2_io_next_header_35 : _GEN_1510; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1575 = 3'h2 == encoders_2_io_output ? proc_2_io_next_header_36 : _GEN_1511; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1576 = 3'h2 == encoders_2_io_output ? proc_2_io_next_header_37 : _GEN_1512; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1577 = 3'h2 == encoders_2_io_output ? proc_2_io_next_header_38 : _GEN_1513; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1578 = 3'h2 == encoders_2_io_output ? proc_2_io_next_header_39 : _GEN_1514; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1579 = 3'h2 == encoders_2_io_output ? proc_2_io_next_header_40 : _GEN_1515; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1580 = 3'h2 == encoders_2_io_output ? proc_2_io_next_header_41 : _GEN_1516; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1581 = 3'h2 == encoders_2_io_output ? proc_2_io_next_header_42 : _GEN_1517; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1582 = 3'h2 == encoders_2_io_output ? proc_2_io_next_header_43 : _GEN_1518; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1583 = 3'h2 == encoders_2_io_output ? proc_2_io_next_header_44 : _GEN_1519; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1584 = 3'h2 == encoders_2_io_output ? proc_2_io_next_header_45 : _GEN_1520; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1585 = 3'h2 == encoders_2_io_output ? proc_2_io_next_header_46 : _GEN_1521; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1586 = 3'h2 == encoders_2_io_output ? proc_2_io_next_header_47 : _GEN_1522; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1587 = 3'h2 == encoders_2_io_output ? proc_2_io_next_header_48 : _GEN_1523; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1588 = 3'h2 == encoders_2_io_output ? proc_2_io_next_header_49 : _GEN_1524; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1589 = 3'h2 == encoders_2_io_output ? proc_2_io_next_header_50 : _GEN_1525; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1590 = 3'h2 == encoders_2_io_output ? proc_2_io_next_header_51 : _GEN_1526; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1591 = 3'h2 == encoders_2_io_output ? proc_2_io_next_header_52 : _GEN_1527; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1592 = 3'h2 == encoders_2_io_output ? proc_2_io_next_header_53 : _GEN_1528; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1593 = 3'h2 == encoders_2_io_output ? proc_2_io_next_header_54 : _GEN_1529; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1594 = 3'h2 == encoders_2_io_output ? proc_2_io_next_header_55 : _GEN_1530; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1595 = 3'h2 == encoders_2_io_output ? proc_2_io_next_header_56 : _GEN_1531; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1596 = 3'h2 == encoders_2_io_output ? proc_2_io_next_header_57 : _GEN_1532; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1597 = 3'h2 == encoders_2_io_output ? proc_2_io_next_header_58 : _GEN_1533; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1598 = 3'h2 == encoders_2_io_output ? proc_2_io_next_header_59 : _GEN_1534; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1599 = 3'h2 == encoders_2_io_output ? proc_2_io_next_header_60 : _GEN_1535; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1600 = 3'h2 == encoders_2_io_output ? proc_2_io_next_header_61 : _GEN_1536; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1601 = 3'h2 == encoders_2_io_output ? proc_2_io_next_header_62 : _GEN_1537; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1602 = 3'h2 == encoders_2_io_output ? proc_2_io_next_header_63 : _GEN_1538; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1603 = 3'h3 == encoders_2_io_output ? proc_3_io_next_header_0 : _GEN_1539; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1604 = 3'h3 == encoders_2_io_output ? proc_3_io_next_header_1 : _GEN_1540; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1605 = 3'h3 == encoders_2_io_output ? proc_3_io_next_header_2 : _GEN_1541; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1606 = 3'h3 == encoders_2_io_output ? proc_3_io_next_header_3 : _GEN_1542; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1607 = 3'h3 == encoders_2_io_output ? proc_3_io_next_header_4 : _GEN_1543; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1608 = 3'h3 == encoders_2_io_output ? proc_3_io_next_header_5 : _GEN_1544; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1609 = 3'h3 == encoders_2_io_output ? proc_3_io_next_header_6 : _GEN_1545; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1610 = 3'h3 == encoders_2_io_output ? proc_3_io_next_header_7 : _GEN_1546; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1611 = 3'h3 == encoders_2_io_output ? proc_3_io_next_header_8 : _GEN_1547; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1612 = 3'h3 == encoders_2_io_output ? proc_3_io_next_header_9 : _GEN_1548; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1613 = 3'h3 == encoders_2_io_output ? proc_3_io_next_header_10 : _GEN_1549; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1614 = 3'h3 == encoders_2_io_output ? proc_3_io_next_header_11 : _GEN_1550; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1615 = 3'h3 == encoders_2_io_output ? proc_3_io_next_header_12 : _GEN_1551; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1616 = 3'h3 == encoders_2_io_output ? proc_3_io_next_header_13 : _GEN_1552; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1617 = 3'h3 == encoders_2_io_output ? proc_3_io_next_header_14 : _GEN_1553; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1618 = 3'h3 == encoders_2_io_output ? proc_3_io_next_header_15 : _GEN_1554; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1619 = 3'h3 == encoders_2_io_output ? proc_3_io_next_header_16 : _GEN_1555; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1620 = 3'h3 == encoders_2_io_output ? proc_3_io_next_header_17 : _GEN_1556; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1621 = 3'h3 == encoders_2_io_output ? proc_3_io_next_header_18 : _GEN_1557; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1622 = 3'h3 == encoders_2_io_output ? proc_3_io_next_header_19 : _GEN_1558; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1623 = 3'h3 == encoders_2_io_output ? proc_3_io_next_header_20 : _GEN_1559; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1624 = 3'h3 == encoders_2_io_output ? proc_3_io_next_header_21 : _GEN_1560; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1625 = 3'h3 == encoders_2_io_output ? proc_3_io_next_header_22 : _GEN_1561; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1626 = 3'h3 == encoders_2_io_output ? proc_3_io_next_header_23 : _GEN_1562; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1627 = 3'h3 == encoders_2_io_output ? proc_3_io_next_header_24 : _GEN_1563; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1628 = 3'h3 == encoders_2_io_output ? proc_3_io_next_header_25 : _GEN_1564; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1629 = 3'h3 == encoders_2_io_output ? proc_3_io_next_header_26 : _GEN_1565; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1630 = 3'h3 == encoders_2_io_output ? proc_3_io_next_header_27 : _GEN_1566; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1631 = 3'h3 == encoders_2_io_output ? proc_3_io_next_header_28 : _GEN_1567; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1632 = 3'h3 == encoders_2_io_output ? proc_3_io_next_header_29 : _GEN_1568; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1633 = 3'h3 == encoders_2_io_output ? proc_3_io_next_header_30 : _GEN_1569; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1634 = 3'h3 == encoders_2_io_output ? proc_3_io_next_header_31 : _GEN_1570; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1635 = 3'h3 == encoders_2_io_output ? proc_3_io_next_header_32 : _GEN_1571; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1636 = 3'h3 == encoders_2_io_output ? proc_3_io_next_header_33 : _GEN_1572; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1637 = 3'h3 == encoders_2_io_output ? proc_3_io_next_header_34 : _GEN_1573; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1638 = 3'h3 == encoders_2_io_output ? proc_3_io_next_header_35 : _GEN_1574; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1639 = 3'h3 == encoders_2_io_output ? proc_3_io_next_header_36 : _GEN_1575; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1640 = 3'h3 == encoders_2_io_output ? proc_3_io_next_header_37 : _GEN_1576; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1641 = 3'h3 == encoders_2_io_output ? proc_3_io_next_header_38 : _GEN_1577; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1642 = 3'h3 == encoders_2_io_output ? proc_3_io_next_header_39 : _GEN_1578; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1643 = 3'h3 == encoders_2_io_output ? proc_3_io_next_header_40 : _GEN_1579; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1644 = 3'h3 == encoders_2_io_output ? proc_3_io_next_header_41 : _GEN_1580; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1645 = 3'h3 == encoders_2_io_output ? proc_3_io_next_header_42 : _GEN_1581; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1646 = 3'h3 == encoders_2_io_output ? proc_3_io_next_header_43 : _GEN_1582; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1647 = 3'h3 == encoders_2_io_output ? proc_3_io_next_header_44 : _GEN_1583; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1648 = 3'h3 == encoders_2_io_output ? proc_3_io_next_header_45 : _GEN_1584; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1649 = 3'h3 == encoders_2_io_output ? proc_3_io_next_header_46 : _GEN_1585; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1650 = 3'h3 == encoders_2_io_output ? proc_3_io_next_header_47 : _GEN_1586; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1651 = 3'h3 == encoders_2_io_output ? proc_3_io_next_header_48 : _GEN_1587; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1652 = 3'h3 == encoders_2_io_output ? proc_3_io_next_header_49 : _GEN_1588; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1653 = 3'h3 == encoders_2_io_output ? proc_3_io_next_header_50 : _GEN_1589; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1654 = 3'h3 == encoders_2_io_output ? proc_3_io_next_header_51 : _GEN_1590; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1655 = 3'h3 == encoders_2_io_output ? proc_3_io_next_header_52 : _GEN_1591; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1656 = 3'h3 == encoders_2_io_output ? proc_3_io_next_header_53 : _GEN_1592; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1657 = 3'h3 == encoders_2_io_output ? proc_3_io_next_header_54 : _GEN_1593; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1658 = 3'h3 == encoders_2_io_output ? proc_3_io_next_header_55 : _GEN_1594; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1659 = 3'h3 == encoders_2_io_output ? proc_3_io_next_header_56 : _GEN_1595; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1660 = 3'h3 == encoders_2_io_output ? proc_3_io_next_header_57 : _GEN_1596; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1661 = 3'h3 == encoders_2_io_output ? proc_3_io_next_header_58 : _GEN_1597; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1662 = 3'h3 == encoders_2_io_output ? proc_3_io_next_header_59 : _GEN_1598; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1663 = 3'h3 == encoders_2_io_output ? proc_3_io_next_header_60 : _GEN_1599; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1664 = 3'h3 == encoders_2_io_output ? proc_3_io_next_header_61 : _GEN_1600; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1665 = 3'h3 == encoders_2_io_output ? proc_3_io_next_header_62 : _GEN_1601; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1666 = 3'h3 == encoders_2_io_output ? proc_3_io_next_header_63 : _GEN_1602; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1667 = 3'h4 == encoders_2_io_output ? proc_4_io_next_header_0 : _GEN_1603; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1668 = 3'h4 == encoders_2_io_output ? proc_4_io_next_header_1 : _GEN_1604; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1669 = 3'h4 == encoders_2_io_output ? proc_4_io_next_header_2 : _GEN_1605; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1670 = 3'h4 == encoders_2_io_output ? proc_4_io_next_header_3 : _GEN_1606; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1671 = 3'h4 == encoders_2_io_output ? proc_4_io_next_header_4 : _GEN_1607; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1672 = 3'h4 == encoders_2_io_output ? proc_4_io_next_header_5 : _GEN_1608; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1673 = 3'h4 == encoders_2_io_output ? proc_4_io_next_header_6 : _GEN_1609; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1674 = 3'h4 == encoders_2_io_output ? proc_4_io_next_header_7 : _GEN_1610; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1675 = 3'h4 == encoders_2_io_output ? proc_4_io_next_header_8 : _GEN_1611; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1676 = 3'h4 == encoders_2_io_output ? proc_4_io_next_header_9 : _GEN_1612; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1677 = 3'h4 == encoders_2_io_output ? proc_4_io_next_header_10 : _GEN_1613; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1678 = 3'h4 == encoders_2_io_output ? proc_4_io_next_header_11 : _GEN_1614; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1679 = 3'h4 == encoders_2_io_output ? proc_4_io_next_header_12 : _GEN_1615; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1680 = 3'h4 == encoders_2_io_output ? proc_4_io_next_header_13 : _GEN_1616; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1681 = 3'h4 == encoders_2_io_output ? proc_4_io_next_header_14 : _GEN_1617; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1682 = 3'h4 == encoders_2_io_output ? proc_4_io_next_header_15 : _GEN_1618; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1683 = 3'h4 == encoders_2_io_output ? proc_4_io_next_header_16 : _GEN_1619; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1684 = 3'h4 == encoders_2_io_output ? proc_4_io_next_header_17 : _GEN_1620; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1685 = 3'h4 == encoders_2_io_output ? proc_4_io_next_header_18 : _GEN_1621; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1686 = 3'h4 == encoders_2_io_output ? proc_4_io_next_header_19 : _GEN_1622; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1687 = 3'h4 == encoders_2_io_output ? proc_4_io_next_header_20 : _GEN_1623; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1688 = 3'h4 == encoders_2_io_output ? proc_4_io_next_header_21 : _GEN_1624; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1689 = 3'h4 == encoders_2_io_output ? proc_4_io_next_header_22 : _GEN_1625; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1690 = 3'h4 == encoders_2_io_output ? proc_4_io_next_header_23 : _GEN_1626; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1691 = 3'h4 == encoders_2_io_output ? proc_4_io_next_header_24 : _GEN_1627; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1692 = 3'h4 == encoders_2_io_output ? proc_4_io_next_header_25 : _GEN_1628; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1693 = 3'h4 == encoders_2_io_output ? proc_4_io_next_header_26 : _GEN_1629; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1694 = 3'h4 == encoders_2_io_output ? proc_4_io_next_header_27 : _GEN_1630; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1695 = 3'h4 == encoders_2_io_output ? proc_4_io_next_header_28 : _GEN_1631; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1696 = 3'h4 == encoders_2_io_output ? proc_4_io_next_header_29 : _GEN_1632; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1697 = 3'h4 == encoders_2_io_output ? proc_4_io_next_header_30 : _GEN_1633; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1698 = 3'h4 == encoders_2_io_output ? proc_4_io_next_header_31 : _GEN_1634; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1699 = 3'h4 == encoders_2_io_output ? proc_4_io_next_header_32 : _GEN_1635; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1700 = 3'h4 == encoders_2_io_output ? proc_4_io_next_header_33 : _GEN_1636; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1701 = 3'h4 == encoders_2_io_output ? proc_4_io_next_header_34 : _GEN_1637; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1702 = 3'h4 == encoders_2_io_output ? proc_4_io_next_header_35 : _GEN_1638; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1703 = 3'h4 == encoders_2_io_output ? proc_4_io_next_header_36 : _GEN_1639; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1704 = 3'h4 == encoders_2_io_output ? proc_4_io_next_header_37 : _GEN_1640; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1705 = 3'h4 == encoders_2_io_output ? proc_4_io_next_header_38 : _GEN_1641; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1706 = 3'h4 == encoders_2_io_output ? proc_4_io_next_header_39 : _GEN_1642; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1707 = 3'h4 == encoders_2_io_output ? proc_4_io_next_header_40 : _GEN_1643; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1708 = 3'h4 == encoders_2_io_output ? proc_4_io_next_header_41 : _GEN_1644; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1709 = 3'h4 == encoders_2_io_output ? proc_4_io_next_header_42 : _GEN_1645; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1710 = 3'h4 == encoders_2_io_output ? proc_4_io_next_header_43 : _GEN_1646; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1711 = 3'h4 == encoders_2_io_output ? proc_4_io_next_header_44 : _GEN_1647; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1712 = 3'h4 == encoders_2_io_output ? proc_4_io_next_header_45 : _GEN_1648; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1713 = 3'h4 == encoders_2_io_output ? proc_4_io_next_header_46 : _GEN_1649; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1714 = 3'h4 == encoders_2_io_output ? proc_4_io_next_header_47 : _GEN_1650; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1715 = 3'h4 == encoders_2_io_output ? proc_4_io_next_header_48 : _GEN_1651; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1716 = 3'h4 == encoders_2_io_output ? proc_4_io_next_header_49 : _GEN_1652; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1717 = 3'h4 == encoders_2_io_output ? proc_4_io_next_header_50 : _GEN_1653; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1718 = 3'h4 == encoders_2_io_output ? proc_4_io_next_header_51 : _GEN_1654; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1719 = 3'h4 == encoders_2_io_output ? proc_4_io_next_header_52 : _GEN_1655; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1720 = 3'h4 == encoders_2_io_output ? proc_4_io_next_header_53 : _GEN_1656; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1721 = 3'h4 == encoders_2_io_output ? proc_4_io_next_header_54 : _GEN_1657; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1722 = 3'h4 == encoders_2_io_output ? proc_4_io_next_header_55 : _GEN_1658; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1723 = 3'h4 == encoders_2_io_output ? proc_4_io_next_header_56 : _GEN_1659; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1724 = 3'h4 == encoders_2_io_output ? proc_4_io_next_header_57 : _GEN_1660; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1725 = 3'h4 == encoders_2_io_output ? proc_4_io_next_header_58 : _GEN_1661; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1726 = 3'h4 == encoders_2_io_output ? proc_4_io_next_header_59 : _GEN_1662; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1727 = 3'h4 == encoders_2_io_output ? proc_4_io_next_header_60 : _GEN_1663; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1728 = 3'h4 == encoders_2_io_output ? proc_4_io_next_header_61 : _GEN_1664; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1729 = 3'h4 == encoders_2_io_output ? proc_4_io_next_header_62 : _GEN_1665; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1730 = 3'h4 == encoders_2_io_output ? proc_4_io_next_header_63 : _GEN_1666; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1731 = 3'h5 == encoders_2_io_output ? proc_5_io_next_header_0 : _GEN_1667; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1732 = 3'h5 == encoders_2_io_output ? proc_5_io_next_header_1 : _GEN_1668; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1733 = 3'h5 == encoders_2_io_output ? proc_5_io_next_header_2 : _GEN_1669; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1734 = 3'h5 == encoders_2_io_output ? proc_5_io_next_header_3 : _GEN_1670; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1735 = 3'h5 == encoders_2_io_output ? proc_5_io_next_header_4 : _GEN_1671; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1736 = 3'h5 == encoders_2_io_output ? proc_5_io_next_header_5 : _GEN_1672; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1737 = 3'h5 == encoders_2_io_output ? proc_5_io_next_header_6 : _GEN_1673; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1738 = 3'h5 == encoders_2_io_output ? proc_5_io_next_header_7 : _GEN_1674; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1739 = 3'h5 == encoders_2_io_output ? proc_5_io_next_header_8 : _GEN_1675; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1740 = 3'h5 == encoders_2_io_output ? proc_5_io_next_header_9 : _GEN_1676; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1741 = 3'h5 == encoders_2_io_output ? proc_5_io_next_header_10 : _GEN_1677; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1742 = 3'h5 == encoders_2_io_output ? proc_5_io_next_header_11 : _GEN_1678; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1743 = 3'h5 == encoders_2_io_output ? proc_5_io_next_header_12 : _GEN_1679; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1744 = 3'h5 == encoders_2_io_output ? proc_5_io_next_header_13 : _GEN_1680; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1745 = 3'h5 == encoders_2_io_output ? proc_5_io_next_header_14 : _GEN_1681; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1746 = 3'h5 == encoders_2_io_output ? proc_5_io_next_header_15 : _GEN_1682; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1747 = 3'h5 == encoders_2_io_output ? proc_5_io_next_header_16 : _GEN_1683; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1748 = 3'h5 == encoders_2_io_output ? proc_5_io_next_header_17 : _GEN_1684; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1749 = 3'h5 == encoders_2_io_output ? proc_5_io_next_header_18 : _GEN_1685; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1750 = 3'h5 == encoders_2_io_output ? proc_5_io_next_header_19 : _GEN_1686; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1751 = 3'h5 == encoders_2_io_output ? proc_5_io_next_header_20 : _GEN_1687; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1752 = 3'h5 == encoders_2_io_output ? proc_5_io_next_header_21 : _GEN_1688; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1753 = 3'h5 == encoders_2_io_output ? proc_5_io_next_header_22 : _GEN_1689; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1754 = 3'h5 == encoders_2_io_output ? proc_5_io_next_header_23 : _GEN_1690; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1755 = 3'h5 == encoders_2_io_output ? proc_5_io_next_header_24 : _GEN_1691; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1756 = 3'h5 == encoders_2_io_output ? proc_5_io_next_header_25 : _GEN_1692; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1757 = 3'h5 == encoders_2_io_output ? proc_5_io_next_header_26 : _GEN_1693; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1758 = 3'h5 == encoders_2_io_output ? proc_5_io_next_header_27 : _GEN_1694; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1759 = 3'h5 == encoders_2_io_output ? proc_5_io_next_header_28 : _GEN_1695; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1760 = 3'h5 == encoders_2_io_output ? proc_5_io_next_header_29 : _GEN_1696; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1761 = 3'h5 == encoders_2_io_output ? proc_5_io_next_header_30 : _GEN_1697; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1762 = 3'h5 == encoders_2_io_output ? proc_5_io_next_header_31 : _GEN_1698; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1763 = 3'h5 == encoders_2_io_output ? proc_5_io_next_header_32 : _GEN_1699; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1764 = 3'h5 == encoders_2_io_output ? proc_5_io_next_header_33 : _GEN_1700; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1765 = 3'h5 == encoders_2_io_output ? proc_5_io_next_header_34 : _GEN_1701; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1766 = 3'h5 == encoders_2_io_output ? proc_5_io_next_header_35 : _GEN_1702; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1767 = 3'h5 == encoders_2_io_output ? proc_5_io_next_header_36 : _GEN_1703; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1768 = 3'h5 == encoders_2_io_output ? proc_5_io_next_header_37 : _GEN_1704; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1769 = 3'h5 == encoders_2_io_output ? proc_5_io_next_header_38 : _GEN_1705; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1770 = 3'h5 == encoders_2_io_output ? proc_5_io_next_header_39 : _GEN_1706; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1771 = 3'h5 == encoders_2_io_output ? proc_5_io_next_header_40 : _GEN_1707; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1772 = 3'h5 == encoders_2_io_output ? proc_5_io_next_header_41 : _GEN_1708; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1773 = 3'h5 == encoders_2_io_output ? proc_5_io_next_header_42 : _GEN_1709; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1774 = 3'h5 == encoders_2_io_output ? proc_5_io_next_header_43 : _GEN_1710; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1775 = 3'h5 == encoders_2_io_output ? proc_5_io_next_header_44 : _GEN_1711; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1776 = 3'h5 == encoders_2_io_output ? proc_5_io_next_header_45 : _GEN_1712; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1777 = 3'h5 == encoders_2_io_output ? proc_5_io_next_header_46 : _GEN_1713; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1778 = 3'h5 == encoders_2_io_output ? proc_5_io_next_header_47 : _GEN_1714; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1779 = 3'h5 == encoders_2_io_output ? proc_5_io_next_header_48 : _GEN_1715; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1780 = 3'h5 == encoders_2_io_output ? proc_5_io_next_header_49 : _GEN_1716; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1781 = 3'h5 == encoders_2_io_output ? proc_5_io_next_header_50 : _GEN_1717; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1782 = 3'h5 == encoders_2_io_output ? proc_5_io_next_header_51 : _GEN_1718; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1783 = 3'h5 == encoders_2_io_output ? proc_5_io_next_header_52 : _GEN_1719; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1784 = 3'h5 == encoders_2_io_output ? proc_5_io_next_header_53 : _GEN_1720; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1785 = 3'h5 == encoders_2_io_output ? proc_5_io_next_header_54 : _GEN_1721; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1786 = 3'h5 == encoders_2_io_output ? proc_5_io_next_header_55 : _GEN_1722; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1787 = 3'h5 == encoders_2_io_output ? proc_5_io_next_header_56 : _GEN_1723; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1788 = 3'h5 == encoders_2_io_output ? proc_5_io_next_header_57 : _GEN_1724; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1789 = 3'h5 == encoders_2_io_output ? proc_5_io_next_header_58 : _GEN_1725; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1790 = 3'h5 == encoders_2_io_output ? proc_5_io_next_header_59 : _GEN_1726; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1791 = 3'h5 == encoders_2_io_output ? proc_5_io_next_header_60 : _GEN_1727; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1792 = 3'h5 == encoders_2_io_output ? proc_5_io_next_header_61 : _GEN_1728; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1793 = 3'h5 == encoders_2_io_output ? proc_5_io_next_header_62 : _GEN_1729; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1794 = 3'h5 == encoders_2_io_output ? proc_5_io_next_header_63 : _GEN_1730; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1795 = 3'h6 == encoders_2_io_output ? proc_6_io_next_header_0 : _GEN_1731; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1796 = 3'h6 == encoders_2_io_output ? proc_6_io_next_header_1 : _GEN_1732; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1797 = 3'h6 == encoders_2_io_output ? proc_6_io_next_header_2 : _GEN_1733; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1798 = 3'h6 == encoders_2_io_output ? proc_6_io_next_header_3 : _GEN_1734; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1799 = 3'h6 == encoders_2_io_output ? proc_6_io_next_header_4 : _GEN_1735; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1800 = 3'h6 == encoders_2_io_output ? proc_6_io_next_header_5 : _GEN_1736; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1801 = 3'h6 == encoders_2_io_output ? proc_6_io_next_header_6 : _GEN_1737; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1802 = 3'h6 == encoders_2_io_output ? proc_6_io_next_header_7 : _GEN_1738; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1803 = 3'h6 == encoders_2_io_output ? proc_6_io_next_header_8 : _GEN_1739; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1804 = 3'h6 == encoders_2_io_output ? proc_6_io_next_header_9 : _GEN_1740; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1805 = 3'h6 == encoders_2_io_output ? proc_6_io_next_header_10 : _GEN_1741; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1806 = 3'h6 == encoders_2_io_output ? proc_6_io_next_header_11 : _GEN_1742; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1807 = 3'h6 == encoders_2_io_output ? proc_6_io_next_header_12 : _GEN_1743; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1808 = 3'h6 == encoders_2_io_output ? proc_6_io_next_header_13 : _GEN_1744; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1809 = 3'h6 == encoders_2_io_output ? proc_6_io_next_header_14 : _GEN_1745; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1810 = 3'h6 == encoders_2_io_output ? proc_6_io_next_header_15 : _GEN_1746; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1811 = 3'h6 == encoders_2_io_output ? proc_6_io_next_header_16 : _GEN_1747; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1812 = 3'h6 == encoders_2_io_output ? proc_6_io_next_header_17 : _GEN_1748; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1813 = 3'h6 == encoders_2_io_output ? proc_6_io_next_header_18 : _GEN_1749; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1814 = 3'h6 == encoders_2_io_output ? proc_6_io_next_header_19 : _GEN_1750; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1815 = 3'h6 == encoders_2_io_output ? proc_6_io_next_header_20 : _GEN_1751; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1816 = 3'h6 == encoders_2_io_output ? proc_6_io_next_header_21 : _GEN_1752; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1817 = 3'h6 == encoders_2_io_output ? proc_6_io_next_header_22 : _GEN_1753; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1818 = 3'h6 == encoders_2_io_output ? proc_6_io_next_header_23 : _GEN_1754; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1819 = 3'h6 == encoders_2_io_output ? proc_6_io_next_header_24 : _GEN_1755; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1820 = 3'h6 == encoders_2_io_output ? proc_6_io_next_header_25 : _GEN_1756; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1821 = 3'h6 == encoders_2_io_output ? proc_6_io_next_header_26 : _GEN_1757; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1822 = 3'h6 == encoders_2_io_output ? proc_6_io_next_header_27 : _GEN_1758; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1823 = 3'h6 == encoders_2_io_output ? proc_6_io_next_header_28 : _GEN_1759; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1824 = 3'h6 == encoders_2_io_output ? proc_6_io_next_header_29 : _GEN_1760; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1825 = 3'h6 == encoders_2_io_output ? proc_6_io_next_header_30 : _GEN_1761; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1826 = 3'h6 == encoders_2_io_output ? proc_6_io_next_header_31 : _GEN_1762; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1827 = 3'h6 == encoders_2_io_output ? proc_6_io_next_header_32 : _GEN_1763; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1828 = 3'h6 == encoders_2_io_output ? proc_6_io_next_header_33 : _GEN_1764; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1829 = 3'h6 == encoders_2_io_output ? proc_6_io_next_header_34 : _GEN_1765; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1830 = 3'h6 == encoders_2_io_output ? proc_6_io_next_header_35 : _GEN_1766; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1831 = 3'h6 == encoders_2_io_output ? proc_6_io_next_header_36 : _GEN_1767; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1832 = 3'h6 == encoders_2_io_output ? proc_6_io_next_header_37 : _GEN_1768; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1833 = 3'h6 == encoders_2_io_output ? proc_6_io_next_header_38 : _GEN_1769; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1834 = 3'h6 == encoders_2_io_output ? proc_6_io_next_header_39 : _GEN_1770; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1835 = 3'h6 == encoders_2_io_output ? proc_6_io_next_header_40 : _GEN_1771; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1836 = 3'h6 == encoders_2_io_output ? proc_6_io_next_header_41 : _GEN_1772; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1837 = 3'h6 == encoders_2_io_output ? proc_6_io_next_header_42 : _GEN_1773; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1838 = 3'h6 == encoders_2_io_output ? proc_6_io_next_header_43 : _GEN_1774; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1839 = 3'h6 == encoders_2_io_output ? proc_6_io_next_header_44 : _GEN_1775; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1840 = 3'h6 == encoders_2_io_output ? proc_6_io_next_header_45 : _GEN_1776; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1841 = 3'h6 == encoders_2_io_output ? proc_6_io_next_header_46 : _GEN_1777; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1842 = 3'h6 == encoders_2_io_output ? proc_6_io_next_header_47 : _GEN_1778; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1843 = 3'h6 == encoders_2_io_output ? proc_6_io_next_header_48 : _GEN_1779; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1844 = 3'h6 == encoders_2_io_output ? proc_6_io_next_header_49 : _GEN_1780; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1845 = 3'h6 == encoders_2_io_output ? proc_6_io_next_header_50 : _GEN_1781; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1846 = 3'h6 == encoders_2_io_output ? proc_6_io_next_header_51 : _GEN_1782; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1847 = 3'h6 == encoders_2_io_output ? proc_6_io_next_header_52 : _GEN_1783; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1848 = 3'h6 == encoders_2_io_output ? proc_6_io_next_header_53 : _GEN_1784; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1849 = 3'h6 == encoders_2_io_output ? proc_6_io_next_header_54 : _GEN_1785; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1850 = 3'h6 == encoders_2_io_output ? proc_6_io_next_header_55 : _GEN_1786; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1851 = 3'h6 == encoders_2_io_output ? proc_6_io_next_header_56 : _GEN_1787; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1852 = 3'h6 == encoders_2_io_output ? proc_6_io_next_header_57 : _GEN_1788; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1853 = 3'h6 == encoders_2_io_output ? proc_6_io_next_header_58 : _GEN_1789; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1854 = 3'h6 == encoders_2_io_output ? proc_6_io_next_header_59 : _GEN_1790; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1855 = 3'h6 == encoders_2_io_output ? proc_6_io_next_header_60 : _GEN_1791; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1856 = 3'h6 == encoders_2_io_output ? proc_6_io_next_header_61 : _GEN_1792; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1857 = 3'h6 == encoders_2_io_output ? proc_6_io_next_header_62 : _GEN_1793; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1858 = 3'h6 == encoders_2_io_output ? proc_6_io_next_header_63 : _GEN_1794; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1859 = 3'h7 == encoders_2_io_output ? proc_7_io_next_header_0 : _GEN_1795; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1860 = 3'h7 == encoders_2_io_output ? proc_7_io_next_header_1 : _GEN_1796; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1861 = 3'h7 == encoders_2_io_output ? proc_7_io_next_header_2 : _GEN_1797; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1862 = 3'h7 == encoders_2_io_output ? proc_7_io_next_header_3 : _GEN_1798; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1863 = 3'h7 == encoders_2_io_output ? proc_7_io_next_header_4 : _GEN_1799; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1864 = 3'h7 == encoders_2_io_output ? proc_7_io_next_header_5 : _GEN_1800; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1865 = 3'h7 == encoders_2_io_output ? proc_7_io_next_header_6 : _GEN_1801; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1866 = 3'h7 == encoders_2_io_output ? proc_7_io_next_header_7 : _GEN_1802; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1867 = 3'h7 == encoders_2_io_output ? proc_7_io_next_header_8 : _GEN_1803; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1868 = 3'h7 == encoders_2_io_output ? proc_7_io_next_header_9 : _GEN_1804; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1869 = 3'h7 == encoders_2_io_output ? proc_7_io_next_header_10 : _GEN_1805; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1870 = 3'h7 == encoders_2_io_output ? proc_7_io_next_header_11 : _GEN_1806; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1871 = 3'h7 == encoders_2_io_output ? proc_7_io_next_header_12 : _GEN_1807; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1872 = 3'h7 == encoders_2_io_output ? proc_7_io_next_header_13 : _GEN_1808; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1873 = 3'h7 == encoders_2_io_output ? proc_7_io_next_header_14 : _GEN_1809; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1874 = 3'h7 == encoders_2_io_output ? proc_7_io_next_header_15 : _GEN_1810; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1875 = 3'h7 == encoders_2_io_output ? proc_7_io_next_header_16 : _GEN_1811; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1876 = 3'h7 == encoders_2_io_output ? proc_7_io_next_header_17 : _GEN_1812; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1877 = 3'h7 == encoders_2_io_output ? proc_7_io_next_header_18 : _GEN_1813; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1878 = 3'h7 == encoders_2_io_output ? proc_7_io_next_header_19 : _GEN_1814; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1879 = 3'h7 == encoders_2_io_output ? proc_7_io_next_header_20 : _GEN_1815; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1880 = 3'h7 == encoders_2_io_output ? proc_7_io_next_header_21 : _GEN_1816; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1881 = 3'h7 == encoders_2_io_output ? proc_7_io_next_header_22 : _GEN_1817; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1882 = 3'h7 == encoders_2_io_output ? proc_7_io_next_header_23 : _GEN_1818; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1883 = 3'h7 == encoders_2_io_output ? proc_7_io_next_header_24 : _GEN_1819; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1884 = 3'h7 == encoders_2_io_output ? proc_7_io_next_header_25 : _GEN_1820; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1885 = 3'h7 == encoders_2_io_output ? proc_7_io_next_header_26 : _GEN_1821; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1886 = 3'h7 == encoders_2_io_output ? proc_7_io_next_header_27 : _GEN_1822; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1887 = 3'h7 == encoders_2_io_output ? proc_7_io_next_header_28 : _GEN_1823; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1888 = 3'h7 == encoders_2_io_output ? proc_7_io_next_header_29 : _GEN_1824; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1889 = 3'h7 == encoders_2_io_output ? proc_7_io_next_header_30 : _GEN_1825; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1890 = 3'h7 == encoders_2_io_output ? proc_7_io_next_header_31 : _GEN_1826; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1891 = 3'h7 == encoders_2_io_output ? proc_7_io_next_header_32 : _GEN_1827; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1892 = 3'h7 == encoders_2_io_output ? proc_7_io_next_header_33 : _GEN_1828; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1893 = 3'h7 == encoders_2_io_output ? proc_7_io_next_header_34 : _GEN_1829; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1894 = 3'h7 == encoders_2_io_output ? proc_7_io_next_header_35 : _GEN_1830; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1895 = 3'h7 == encoders_2_io_output ? proc_7_io_next_header_36 : _GEN_1831; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1896 = 3'h7 == encoders_2_io_output ? proc_7_io_next_header_37 : _GEN_1832; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1897 = 3'h7 == encoders_2_io_output ? proc_7_io_next_header_38 : _GEN_1833; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1898 = 3'h7 == encoders_2_io_output ? proc_7_io_next_header_39 : _GEN_1834; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1899 = 3'h7 == encoders_2_io_output ? proc_7_io_next_header_40 : _GEN_1835; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1900 = 3'h7 == encoders_2_io_output ? proc_7_io_next_header_41 : _GEN_1836; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1901 = 3'h7 == encoders_2_io_output ? proc_7_io_next_header_42 : _GEN_1837; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1902 = 3'h7 == encoders_2_io_output ? proc_7_io_next_header_43 : _GEN_1838; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1903 = 3'h7 == encoders_2_io_output ? proc_7_io_next_header_44 : _GEN_1839; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1904 = 3'h7 == encoders_2_io_output ? proc_7_io_next_header_45 : _GEN_1840; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1905 = 3'h7 == encoders_2_io_output ? proc_7_io_next_header_46 : _GEN_1841; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1906 = 3'h7 == encoders_2_io_output ? proc_7_io_next_header_47 : _GEN_1842; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1907 = 3'h7 == encoders_2_io_output ? proc_7_io_next_header_48 : _GEN_1843; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1908 = 3'h7 == encoders_2_io_output ? proc_7_io_next_header_49 : _GEN_1844; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1909 = 3'h7 == encoders_2_io_output ? proc_7_io_next_header_50 : _GEN_1845; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1910 = 3'h7 == encoders_2_io_output ? proc_7_io_next_header_51 : _GEN_1846; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1911 = 3'h7 == encoders_2_io_output ? proc_7_io_next_header_52 : _GEN_1847; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1912 = 3'h7 == encoders_2_io_output ? proc_7_io_next_header_53 : _GEN_1848; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1913 = 3'h7 == encoders_2_io_output ? proc_7_io_next_header_54 : _GEN_1849; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1914 = 3'h7 == encoders_2_io_output ? proc_7_io_next_header_55 : _GEN_1850; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1915 = 3'h7 == encoders_2_io_output ? proc_7_io_next_header_56 : _GEN_1851; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1916 = 3'h7 == encoders_2_io_output ? proc_7_io_next_header_57 : _GEN_1852; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1917 = 3'h7 == encoders_2_io_output ? proc_7_io_next_header_58 : _GEN_1853; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1918 = 3'h7 == encoders_2_io_output ? proc_7_io_next_header_59 : _GEN_1854; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1919 = 3'h7 == encoders_2_io_output ? proc_7_io_next_header_60 : _GEN_1855; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1920 = 3'h7 == encoders_2_io_output ? proc_7_io_next_header_61 : _GEN_1856; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1921 = 3'h7 == encoders_2_io_output ? proc_7_io_next_header_62 : _GEN_1857; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1922 = 3'h7 == encoders_2_io_output ? proc_7_io_next_header_63 : _GEN_1858; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_1988 = 3'h0 == encoders_3_io_output ? proc_0_io_next_header_0 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1989 = 3'h0 == encoders_3_io_output ? proc_0_io_next_header_1 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1990 = 3'h0 == encoders_3_io_output ? proc_0_io_next_header_2 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1991 = 3'h0 == encoders_3_io_output ? proc_0_io_next_header_3 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1992 = 3'h0 == encoders_3_io_output ? proc_0_io_next_header_4 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1993 = 3'h0 == encoders_3_io_output ? proc_0_io_next_header_5 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1994 = 3'h0 == encoders_3_io_output ? proc_0_io_next_header_6 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1995 = 3'h0 == encoders_3_io_output ? proc_0_io_next_header_7 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1996 = 3'h0 == encoders_3_io_output ? proc_0_io_next_header_8 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1997 = 3'h0 == encoders_3_io_output ? proc_0_io_next_header_9 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1998 = 3'h0 == encoders_3_io_output ? proc_0_io_next_header_10 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_1999 = 3'h0 == encoders_3_io_output ? proc_0_io_next_header_11 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2000 = 3'h0 == encoders_3_io_output ? proc_0_io_next_header_12 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2001 = 3'h0 == encoders_3_io_output ? proc_0_io_next_header_13 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2002 = 3'h0 == encoders_3_io_output ? proc_0_io_next_header_14 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2003 = 3'h0 == encoders_3_io_output ? proc_0_io_next_header_15 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2004 = 3'h0 == encoders_3_io_output ? proc_0_io_next_header_16 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2005 = 3'h0 == encoders_3_io_output ? proc_0_io_next_header_17 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2006 = 3'h0 == encoders_3_io_output ? proc_0_io_next_header_18 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2007 = 3'h0 == encoders_3_io_output ? proc_0_io_next_header_19 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2008 = 3'h0 == encoders_3_io_output ? proc_0_io_next_header_20 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2009 = 3'h0 == encoders_3_io_output ? proc_0_io_next_header_21 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2010 = 3'h0 == encoders_3_io_output ? proc_0_io_next_header_22 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2011 = 3'h0 == encoders_3_io_output ? proc_0_io_next_header_23 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2012 = 3'h0 == encoders_3_io_output ? proc_0_io_next_header_24 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2013 = 3'h0 == encoders_3_io_output ? proc_0_io_next_header_25 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2014 = 3'h0 == encoders_3_io_output ? proc_0_io_next_header_26 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2015 = 3'h0 == encoders_3_io_output ? proc_0_io_next_header_27 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2016 = 3'h0 == encoders_3_io_output ? proc_0_io_next_header_28 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2017 = 3'h0 == encoders_3_io_output ? proc_0_io_next_header_29 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2018 = 3'h0 == encoders_3_io_output ? proc_0_io_next_header_30 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2019 = 3'h0 == encoders_3_io_output ? proc_0_io_next_header_31 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2020 = 3'h0 == encoders_3_io_output ? proc_0_io_next_header_32 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2021 = 3'h0 == encoders_3_io_output ? proc_0_io_next_header_33 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2022 = 3'h0 == encoders_3_io_output ? proc_0_io_next_header_34 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2023 = 3'h0 == encoders_3_io_output ? proc_0_io_next_header_35 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2024 = 3'h0 == encoders_3_io_output ? proc_0_io_next_header_36 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2025 = 3'h0 == encoders_3_io_output ? proc_0_io_next_header_37 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2026 = 3'h0 == encoders_3_io_output ? proc_0_io_next_header_38 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2027 = 3'h0 == encoders_3_io_output ? proc_0_io_next_header_39 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2028 = 3'h0 == encoders_3_io_output ? proc_0_io_next_header_40 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2029 = 3'h0 == encoders_3_io_output ? proc_0_io_next_header_41 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2030 = 3'h0 == encoders_3_io_output ? proc_0_io_next_header_42 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2031 = 3'h0 == encoders_3_io_output ? proc_0_io_next_header_43 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2032 = 3'h0 == encoders_3_io_output ? proc_0_io_next_header_44 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2033 = 3'h0 == encoders_3_io_output ? proc_0_io_next_header_45 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2034 = 3'h0 == encoders_3_io_output ? proc_0_io_next_header_46 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2035 = 3'h0 == encoders_3_io_output ? proc_0_io_next_header_47 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2036 = 3'h0 == encoders_3_io_output ? proc_0_io_next_header_48 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2037 = 3'h0 == encoders_3_io_output ? proc_0_io_next_header_49 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2038 = 3'h0 == encoders_3_io_output ? proc_0_io_next_header_50 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2039 = 3'h0 == encoders_3_io_output ? proc_0_io_next_header_51 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2040 = 3'h0 == encoders_3_io_output ? proc_0_io_next_header_52 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2041 = 3'h0 == encoders_3_io_output ? proc_0_io_next_header_53 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2042 = 3'h0 == encoders_3_io_output ? proc_0_io_next_header_54 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2043 = 3'h0 == encoders_3_io_output ? proc_0_io_next_header_55 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2044 = 3'h0 == encoders_3_io_output ? proc_0_io_next_header_56 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2045 = 3'h0 == encoders_3_io_output ? proc_0_io_next_header_57 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2046 = 3'h0 == encoders_3_io_output ? proc_0_io_next_header_58 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2047 = 3'h0 == encoders_3_io_output ? proc_0_io_next_header_59 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2048 = 3'h0 == encoders_3_io_output ? proc_0_io_next_header_60 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2049 = 3'h0 == encoders_3_io_output ? proc_0_io_next_header_61 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2050 = 3'h0 == encoders_3_io_output ? proc_0_io_next_header_62 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2051 = 3'h0 == encoders_3_io_output ? proc_0_io_next_header_63 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2052 = 3'h1 == encoders_3_io_output ? proc_1_io_next_header_0 : _GEN_1988; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2053 = 3'h1 == encoders_3_io_output ? proc_1_io_next_header_1 : _GEN_1989; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2054 = 3'h1 == encoders_3_io_output ? proc_1_io_next_header_2 : _GEN_1990; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2055 = 3'h1 == encoders_3_io_output ? proc_1_io_next_header_3 : _GEN_1991; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2056 = 3'h1 == encoders_3_io_output ? proc_1_io_next_header_4 : _GEN_1992; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2057 = 3'h1 == encoders_3_io_output ? proc_1_io_next_header_5 : _GEN_1993; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2058 = 3'h1 == encoders_3_io_output ? proc_1_io_next_header_6 : _GEN_1994; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2059 = 3'h1 == encoders_3_io_output ? proc_1_io_next_header_7 : _GEN_1995; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2060 = 3'h1 == encoders_3_io_output ? proc_1_io_next_header_8 : _GEN_1996; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2061 = 3'h1 == encoders_3_io_output ? proc_1_io_next_header_9 : _GEN_1997; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2062 = 3'h1 == encoders_3_io_output ? proc_1_io_next_header_10 : _GEN_1998; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2063 = 3'h1 == encoders_3_io_output ? proc_1_io_next_header_11 : _GEN_1999; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2064 = 3'h1 == encoders_3_io_output ? proc_1_io_next_header_12 : _GEN_2000; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2065 = 3'h1 == encoders_3_io_output ? proc_1_io_next_header_13 : _GEN_2001; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2066 = 3'h1 == encoders_3_io_output ? proc_1_io_next_header_14 : _GEN_2002; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2067 = 3'h1 == encoders_3_io_output ? proc_1_io_next_header_15 : _GEN_2003; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2068 = 3'h1 == encoders_3_io_output ? proc_1_io_next_header_16 : _GEN_2004; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2069 = 3'h1 == encoders_3_io_output ? proc_1_io_next_header_17 : _GEN_2005; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2070 = 3'h1 == encoders_3_io_output ? proc_1_io_next_header_18 : _GEN_2006; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2071 = 3'h1 == encoders_3_io_output ? proc_1_io_next_header_19 : _GEN_2007; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2072 = 3'h1 == encoders_3_io_output ? proc_1_io_next_header_20 : _GEN_2008; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2073 = 3'h1 == encoders_3_io_output ? proc_1_io_next_header_21 : _GEN_2009; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2074 = 3'h1 == encoders_3_io_output ? proc_1_io_next_header_22 : _GEN_2010; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2075 = 3'h1 == encoders_3_io_output ? proc_1_io_next_header_23 : _GEN_2011; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2076 = 3'h1 == encoders_3_io_output ? proc_1_io_next_header_24 : _GEN_2012; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2077 = 3'h1 == encoders_3_io_output ? proc_1_io_next_header_25 : _GEN_2013; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2078 = 3'h1 == encoders_3_io_output ? proc_1_io_next_header_26 : _GEN_2014; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2079 = 3'h1 == encoders_3_io_output ? proc_1_io_next_header_27 : _GEN_2015; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2080 = 3'h1 == encoders_3_io_output ? proc_1_io_next_header_28 : _GEN_2016; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2081 = 3'h1 == encoders_3_io_output ? proc_1_io_next_header_29 : _GEN_2017; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2082 = 3'h1 == encoders_3_io_output ? proc_1_io_next_header_30 : _GEN_2018; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2083 = 3'h1 == encoders_3_io_output ? proc_1_io_next_header_31 : _GEN_2019; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2084 = 3'h1 == encoders_3_io_output ? proc_1_io_next_header_32 : _GEN_2020; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2085 = 3'h1 == encoders_3_io_output ? proc_1_io_next_header_33 : _GEN_2021; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2086 = 3'h1 == encoders_3_io_output ? proc_1_io_next_header_34 : _GEN_2022; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2087 = 3'h1 == encoders_3_io_output ? proc_1_io_next_header_35 : _GEN_2023; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2088 = 3'h1 == encoders_3_io_output ? proc_1_io_next_header_36 : _GEN_2024; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2089 = 3'h1 == encoders_3_io_output ? proc_1_io_next_header_37 : _GEN_2025; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2090 = 3'h1 == encoders_3_io_output ? proc_1_io_next_header_38 : _GEN_2026; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2091 = 3'h1 == encoders_3_io_output ? proc_1_io_next_header_39 : _GEN_2027; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2092 = 3'h1 == encoders_3_io_output ? proc_1_io_next_header_40 : _GEN_2028; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2093 = 3'h1 == encoders_3_io_output ? proc_1_io_next_header_41 : _GEN_2029; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2094 = 3'h1 == encoders_3_io_output ? proc_1_io_next_header_42 : _GEN_2030; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2095 = 3'h1 == encoders_3_io_output ? proc_1_io_next_header_43 : _GEN_2031; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2096 = 3'h1 == encoders_3_io_output ? proc_1_io_next_header_44 : _GEN_2032; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2097 = 3'h1 == encoders_3_io_output ? proc_1_io_next_header_45 : _GEN_2033; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2098 = 3'h1 == encoders_3_io_output ? proc_1_io_next_header_46 : _GEN_2034; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2099 = 3'h1 == encoders_3_io_output ? proc_1_io_next_header_47 : _GEN_2035; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2100 = 3'h1 == encoders_3_io_output ? proc_1_io_next_header_48 : _GEN_2036; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2101 = 3'h1 == encoders_3_io_output ? proc_1_io_next_header_49 : _GEN_2037; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2102 = 3'h1 == encoders_3_io_output ? proc_1_io_next_header_50 : _GEN_2038; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2103 = 3'h1 == encoders_3_io_output ? proc_1_io_next_header_51 : _GEN_2039; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2104 = 3'h1 == encoders_3_io_output ? proc_1_io_next_header_52 : _GEN_2040; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2105 = 3'h1 == encoders_3_io_output ? proc_1_io_next_header_53 : _GEN_2041; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2106 = 3'h1 == encoders_3_io_output ? proc_1_io_next_header_54 : _GEN_2042; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2107 = 3'h1 == encoders_3_io_output ? proc_1_io_next_header_55 : _GEN_2043; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2108 = 3'h1 == encoders_3_io_output ? proc_1_io_next_header_56 : _GEN_2044; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2109 = 3'h1 == encoders_3_io_output ? proc_1_io_next_header_57 : _GEN_2045; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2110 = 3'h1 == encoders_3_io_output ? proc_1_io_next_header_58 : _GEN_2046; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2111 = 3'h1 == encoders_3_io_output ? proc_1_io_next_header_59 : _GEN_2047; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2112 = 3'h1 == encoders_3_io_output ? proc_1_io_next_header_60 : _GEN_2048; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2113 = 3'h1 == encoders_3_io_output ? proc_1_io_next_header_61 : _GEN_2049; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2114 = 3'h1 == encoders_3_io_output ? proc_1_io_next_header_62 : _GEN_2050; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2115 = 3'h1 == encoders_3_io_output ? proc_1_io_next_header_63 : _GEN_2051; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2116 = 3'h2 == encoders_3_io_output ? proc_2_io_next_header_0 : _GEN_2052; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2117 = 3'h2 == encoders_3_io_output ? proc_2_io_next_header_1 : _GEN_2053; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2118 = 3'h2 == encoders_3_io_output ? proc_2_io_next_header_2 : _GEN_2054; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2119 = 3'h2 == encoders_3_io_output ? proc_2_io_next_header_3 : _GEN_2055; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2120 = 3'h2 == encoders_3_io_output ? proc_2_io_next_header_4 : _GEN_2056; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2121 = 3'h2 == encoders_3_io_output ? proc_2_io_next_header_5 : _GEN_2057; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2122 = 3'h2 == encoders_3_io_output ? proc_2_io_next_header_6 : _GEN_2058; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2123 = 3'h2 == encoders_3_io_output ? proc_2_io_next_header_7 : _GEN_2059; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2124 = 3'h2 == encoders_3_io_output ? proc_2_io_next_header_8 : _GEN_2060; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2125 = 3'h2 == encoders_3_io_output ? proc_2_io_next_header_9 : _GEN_2061; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2126 = 3'h2 == encoders_3_io_output ? proc_2_io_next_header_10 : _GEN_2062; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2127 = 3'h2 == encoders_3_io_output ? proc_2_io_next_header_11 : _GEN_2063; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2128 = 3'h2 == encoders_3_io_output ? proc_2_io_next_header_12 : _GEN_2064; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2129 = 3'h2 == encoders_3_io_output ? proc_2_io_next_header_13 : _GEN_2065; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2130 = 3'h2 == encoders_3_io_output ? proc_2_io_next_header_14 : _GEN_2066; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2131 = 3'h2 == encoders_3_io_output ? proc_2_io_next_header_15 : _GEN_2067; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2132 = 3'h2 == encoders_3_io_output ? proc_2_io_next_header_16 : _GEN_2068; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2133 = 3'h2 == encoders_3_io_output ? proc_2_io_next_header_17 : _GEN_2069; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2134 = 3'h2 == encoders_3_io_output ? proc_2_io_next_header_18 : _GEN_2070; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2135 = 3'h2 == encoders_3_io_output ? proc_2_io_next_header_19 : _GEN_2071; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2136 = 3'h2 == encoders_3_io_output ? proc_2_io_next_header_20 : _GEN_2072; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2137 = 3'h2 == encoders_3_io_output ? proc_2_io_next_header_21 : _GEN_2073; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2138 = 3'h2 == encoders_3_io_output ? proc_2_io_next_header_22 : _GEN_2074; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2139 = 3'h2 == encoders_3_io_output ? proc_2_io_next_header_23 : _GEN_2075; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2140 = 3'h2 == encoders_3_io_output ? proc_2_io_next_header_24 : _GEN_2076; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2141 = 3'h2 == encoders_3_io_output ? proc_2_io_next_header_25 : _GEN_2077; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2142 = 3'h2 == encoders_3_io_output ? proc_2_io_next_header_26 : _GEN_2078; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2143 = 3'h2 == encoders_3_io_output ? proc_2_io_next_header_27 : _GEN_2079; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2144 = 3'h2 == encoders_3_io_output ? proc_2_io_next_header_28 : _GEN_2080; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2145 = 3'h2 == encoders_3_io_output ? proc_2_io_next_header_29 : _GEN_2081; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2146 = 3'h2 == encoders_3_io_output ? proc_2_io_next_header_30 : _GEN_2082; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2147 = 3'h2 == encoders_3_io_output ? proc_2_io_next_header_31 : _GEN_2083; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2148 = 3'h2 == encoders_3_io_output ? proc_2_io_next_header_32 : _GEN_2084; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2149 = 3'h2 == encoders_3_io_output ? proc_2_io_next_header_33 : _GEN_2085; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2150 = 3'h2 == encoders_3_io_output ? proc_2_io_next_header_34 : _GEN_2086; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2151 = 3'h2 == encoders_3_io_output ? proc_2_io_next_header_35 : _GEN_2087; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2152 = 3'h2 == encoders_3_io_output ? proc_2_io_next_header_36 : _GEN_2088; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2153 = 3'h2 == encoders_3_io_output ? proc_2_io_next_header_37 : _GEN_2089; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2154 = 3'h2 == encoders_3_io_output ? proc_2_io_next_header_38 : _GEN_2090; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2155 = 3'h2 == encoders_3_io_output ? proc_2_io_next_header_39 : _GEN_2091; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2156 = 3'h2 == encoders_3_io_output ? proc_2_io_next_header_40 : _GEN_2092; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2157 = 3'h2 == encoders_3_io_output ? proc_2_io_next_header_41 : _GEN_2093; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2158 = 3'h2 == encoders_3_io_output ? proc_2_io_next_header_42 : _GEN_2094; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2159 = 3'h2 == encoders_3_io_output ? proc_2_io_next_header_43 : _GEN_2095; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2160 = 3'h2 == encoders_3_io_output ? proc_2_io_next_header_44 : _GEN_2096; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2161 = 3'h2 == encoders_3_io_output ? proc_2_io_next_header_45 : _GEN_2097; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2162 = 3'h2 == encoders_3_io_output ? proc_2_io_next_header_46 : _GEN_2098; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2163 = 3'h2 == encoders_3_io_output ? proc_2_io_next_header_47 : _GEN_2099; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2164 = 3'h2 == encoders_3_io_output ? proc_2_io_next_header_48 : _GEN_2100; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2165 = 3'h2 == encoders_3_io_output ? proc_2_io_next_header_49 : _GEN_2101; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2166 = 3'h2 == encoders_3_io_output ? proc_2_io_next_header_50 : _GEN_2102; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2167 = 3'h2 == encoders_3_io_output ? proc_2_io_next_header_51 : _GEN_2103; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2168 = 3'h2 == encoders_3_io_output ? proc_2_io_next_header_52 : _GEN_2104; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2169 = 3'h2 == encoders_3_io_output ? proc_2_io_next_header_53 : _GEN_2105; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2170 = 3'h2 == encoders_3_io_output ? proc_2_io_next_header_54 : _GEN_2106; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2171 = 3'h2 == encoders_3_io_output ? proc_2_io_next_header_55 : _GEN_2107; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2172 = 3'h2 == encoders_3_io_output ? proc_2_io_next_header_56 : _GEN_2108; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2173 = 3'h2 == encoders_3_io_output ? proc_2_io_next_header_57 : _GEN_2109; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2174 = 3'h2 == encoders_3_io_output ? proc_2_io_next_header_58 : _GEN_2110; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2175 = 3'h2 == encoders_3_io_output ? proc_2_io_next_header_59 : _GEN_2111; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2176 = 3'h2 == encoders_3_io_output ? proc_2_io_next_header_60 : _GEN_2112; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2177 = 3'h2 == encoders_3_io_output ? proc_2_io_next_header_61 : _GEN_2113; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2178 = 3'h2 == encoders_3_io_output ? proc_2_io_next_header_62 : _GEN_2114; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2179 = 3'h2 == encoders_3_io_output ? proc_2_io_next_header_63 : _GEN_2115; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2180 = 3'h3 == encoders_3_io_output ? proc_3_io_next_header_0 : _GEN_2116; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2181 = 3'h3 == encoders_3_io_output ? proc_3_io_next_header_1 : _GEN_2117; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2182 = 3'h3 == encoders_3_io_output ? proc_3_io_next_header_2 : _GEN_2118; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2183 = 3'h3 == encoders_3_io_output ? proc_3_io_next_header_3 : _GEN_2119; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2184 = 3'h3 == encoders_3_io_output ? proc_3_io_next_header_4 : _GEN_2120; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2185 = 3'h3 == encoders_3_io_output ? proc_3_io_next_header_5 : _GEN_2121; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2186 = 3'h3 == encoders_3_io_output ? proc_3_io_next_header_6 : _GEN_2122; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2187 = 3'h3 == encoders_3_io_output ? proc_3_io_next_header_7 : _GEN_2123; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2188 = 3'h3 == encoders_3_io_output ? proc_3_io_next_header_8 : _GEN_2124; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2189 = 3'h3 == encoders_3_io_output ? proc_3_io_next_header_9 : _GEN_2125; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2190 = 3'h3 == encoders_3_io_output ? proc_3_io_next_header_10 : _GEN_2126; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2191 = 3'h3 == encoders_3_io_output ? proc_3_io_next_header_11 : _GEN_2127; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2192 = 3'h3 == encoders_3_io_output ? proc_3_io_next_header_12 : _GEN_2128; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2193 = 3'h3 == encoders_3_io_output ? proc_3_io_next_header_13 : _GEN_2129; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2194 = 3'h3 == encoders_3_io_output ? proc_3_io_next_header_14 : _GEN_2130; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2195 = 3'h3 == encoders_3_io_output ? proc_3_io_next_header_15 : _GEN_2131; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2196 = 3'h3 == encoders_3_io_output ? proc_3_io_next_header_16 : _GEN_2132; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2197 = 3'h3 == encoders_3_io_output ? proc_3_io_next_header_17 : _GEN_2133; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2198 = 3'h3 == encoders_3_io_output ? proc_3_io_next_header_18 : _GEN_2134; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2199 = 3'h3 == encoders_3_io_output ? proc_3_io_next_header_19 : _GEN_2135; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2200 = 3'h3 == encoders_3_io_output ? proc_3_io_next_header_20 : _GEN_2136; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2201 = 3'h3 == encoders_3_io_output ? proc_3_io_next_header_21 : _GEN_2137; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2202 = 3'h3 == encoders_3_io_output ? proc_3_io_next_header_22 : _GEN_2138; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2203 = 3'h3 == encoders_3_io_output ? proc_3_io_next_header_23 : _GEN_2139; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2204 = 3'h3 == encoders_3_io_output ? proc_3_io_next_header_24 : _GEN_2140; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2205 = 3'h3 == encoders_3_io_output ? proc_3_io_next_header_25 : _GEN_2141; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2206 = 3'h3 == encoders_3_io_output ? proc_3_io_next_header_26 : _GEN_2142; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2207 = 3'h3 == encoders_3_io_output ? proc_3_io_next_header_27 : _GEN_2143; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2208 = 3'h3 == encoders_3_io_output ? proc_3_io_next_header_28 : _GEN_2144; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2209 = 3'h3 == encoders_3_io_output ? proc_3_io_next_header_29 : _GEN_2145; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2210 = 3'h3 == encoders_3_io_output ? proc_3_io_next_header_30 : _GEN_2146; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2211 = 3'h3 == encoders_3_io_output ? proc_3_io_next_header_31 : _GEN_2147; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2212 = 3'h3 == encoders_3_io_output ? proc_3_io_next_header_32 : _GEN_2148; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2213 = 3'h3 == encoders_3_io_output ? proc_3_io_next_header_33 : _GEN_2149; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2214 = 3'h3 == encoders_3_io_output ? proc_3_io_next_header_34 : _GEN_2150; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2215 = 3'h3 == encoders_3_io_output ? proc_3_io_next_header_35 : _GEN_2151; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2216 = 3'h3 == encoders_3_io_output ? proc_3_io_next_header_36 : _GEN_2152; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2217 = 3'h3 == encoders_3_io_output ? proc_3_io_next_header_37 : _GEN_2153; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2218 = 3'h3 == encoders_3_io_output ? proc_3_io_next_header_38 : _GEN_2154; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2219 = 3'h3 == encoders_3_io_output ? proc_3_io_next_header_39 : _GEN_2155; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2220 = 3'h3 == encoders_3_io_output ? proc_3_io_next_header_40 : _GEN_2156; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2221 = 3'h3 == encoders_3_io_output ? proc_3_io_next_header_41 : _GEN_2157; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2222 = 3'h3 == encoders_3_io_output ? proc_3_io_next_header_42 : _GEN_2158; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2223 = 3'h3 == encoders_3_io_output ? proc_3_io_next_header_43 : _GEN_2159; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2224 = 3'h3 == encoders_3_io_output ? proc_3_io_next_header_44 : _GEN_2160; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2225 = 3'h3 == encoders_3_io_output ? proc_3_io_next_header_45 : _GEN_2161; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2226 = 3'h3 == encoders_3_io_output ? proc_3_io_next_header_46 : _GEN_2162; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2227 = 3'h3 == encoders_3_io_output ? proc_3_io_next_header_47 : _GEN_2163; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2228 = 3'h3 == encoders_3_io_output ? proc_3_io_next_header_48 : _GEN_2164; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2229 = 3'h3 == encoders_3_io_output ? proc_3_io_next_header_49 : _GEN_2165; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2230 = 3'h3 == encoders_3_io_output ? proc_3_io_next_header_50 : _GEN_2166; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2231 = 3'h3 == encoders_3_io_output ? proc_3_io_next_header_51 : _GEN_2167; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2232 = 3'h3 == encoders_3_io_output ? proc_3_io_next_header_52 : _GEN_2168; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2233 = 3'h3 == encoders_3_io_output ? proc_3_io_next_header_53 : _GEN_2169; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2234 = 3'h3 == encoders_3_io_output ? proc_3_io_next_header_54 : _GEN_2170; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2235 = 3'h3 == encoders_3_io_output ? proc_3_io_next_header_55 : _GEN_2171; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2236 = 3'h3 == encoders_3_io_output ? proc_3_io_next_header_56 : _GEN_2172; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2237 = 3'h3 == encoders_3_io_output ? proc_3_io_next_header_57 : _GEN_2173; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2238 = 3'h3 == encoders_3_io_output ? proc_3_io_next_header_58 : _GEN_2174; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2239 = 3'h3 == encoders_3_io_output ? proc_3_io_next_header_59 : _GEN_2175; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2240 = 3'h3 == encoders_3_io_output ? proc_3_io_next_header_60 : _GEN_2176; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2241 = 3'h3 == encoders_3_io_output ? proc_3_io_next_header_61 : _GEN_2177; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2242 = 3'h3 == encoders_3_io_output ? proc_3_io_next_header_62 : _GEN_2178; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2243 = 3'h3 == encoders_3_io_output ? proc_3_io_next_header_63 : _GEN_2179; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2244 = 3'h4 == encoders_3_io_output ? proc_4_io_next_header_0 : _GEN_2180; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2245 = 3'h4 == encoders_3_io_output ? proc_4_io_next_header_1 : _GEN_2181; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2246 = 3'h4 == encoders_3_io_output ? proc_4_io_next_header_2 : _GEN_2182; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2247 = 3'h4 == encoders_3_io_output ? proc_4_io_next_header_3 : _GEN_2183; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2248 = 3'h4 == encoders_3_io_output ? proc_4_io_next_header_4 : _GEN_2184; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2249 = 3'h4 == encoders_3_io_output ? proc_4_io_next_header_5 : _GEN_2185; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2250 = 3'h4 == encoders_3_io_output ? proc_4_io_next_header_6 : _GEN_2186; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2251 = 3'h4 == encoders_3_io_output ? proc_4_io_next_header_7 : _GEN_2187; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2252 = 3'h4 == encoders_3_io_output ? proc_4_io_next_header_8 : _GEN_2188; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2253 = 3'h4 == encoders_3_io_output ? proc_4_io_next_header_9 : _GEN_2189; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2254 = 3'h4 == encoders_3_io_output ? proc_4_io_next_header_10 : _GEN_2190; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2255 = 3'h4 == encoders_3_io_output ? proc_4_io_next_header_11 : _GEN_2191; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2256 = 3'h4 == encoders_3_io_output ? proc_4_io_next_header_12 : _GEN_2192; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2257 = 3'h4 == encoders_3_io_output ? proc_4_io_next_header_13 : _GEN_2193; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2258 = 3'h4 == encoders_3_io_output ? proc_4_io_next_header_14 : _GEN_2194; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2259 = 3'h4 == encoders_3_io_output ? proc_4_io_next_header_15 : _GEN_2195; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2260 = 3'h4 == encoders_3_io_output ? proc_4_io_next_header_16 : _GEN_2196; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2261 = 3'h4 == encoders_3_io_output ? proc_4_io_next_header_17 : _GEN_2197; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2262 = 3'h4 == encoders_3_io_output ? proc_4_io_next_header_18 : _GEN_2198; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2263 = 3'h4 == encoders_3_io_output ? proc_4_io_next_header_19 : _GEN_2199; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2264 = 3'h4 == encoders_3_io_output ? proc_4_io_next_header_20 : _GEN_2200; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2265 = 3'h4 == encoders_3_io_output ? proc_4_io_next_header_21 : _GEN_2201; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2266 = 3'h4 == encoders_3_io_output ? proc_4_io_next_header_22 : _GEN_2202; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2267 = 3'h4 == encoders_3_io_output ? proc_4_io_next_header_23 : _GEN_2203; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2268 = 3'h4 == encoders_3_io_output ? proc_4_io_next_header_24 : _GEN_2204; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2269 = 3'h4 == encoders_3_io_output ? proc_4_io_next_header_25 : _GEN_2205; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2270 = 3'h4 == encoders_3_io_output ? proc_4_io_next_header_26 : _GEN_2206; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2271 = 3'h4 == encoders_3_io_output ? proc_4_io_next_header_27 : _GEN_2207; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2272 = 3'h4 == encoders_3_io_output ? proc_4_io_next_header_28 : _GEN_2208; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2273 = 3'h4 == encoders_3_io_output ? proc_4_io_next_header_29 : _GEN_2209; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2274 = 3'h4 == encoders_3_io_output ? proc_4_io_next_header_30 : _GEN_2210; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2275 = 3'h4 == encoders_3_io_output ? proc_4_io_next_header_31 : _GEN_2211; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2276 = 3'h4 == encoders_3_io_output ? proc_4_io_next_header_32 : _GEN_2212; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2277 = 3'h4 == encoders_3_io_output ? proc_4_io_next_header_33 : _GEN_2213; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2278 = 3'h4 == encoders_3_io_output ? proc_4_io_next_header_34 : _GEN_2214; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2279 = 3'h4 == encoders_3_io_output ? proc_4_io_next_header_35 : _GEN_2215; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2280 = 3'h4 == encoders_3_io_output ? proc_4_io_next_header_36 : _GEN_2216; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2281 = 3'h4 == encoders_3_io_output ? proc_4_io_next_header_37 : _GEN_2217; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2282 = 3'h4 == encoders_3_io_output ? proc_4_io_next_header_38 : _GEN_2218; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2283 = 3'h4 == encoders_3_io_output ? proc_4_io_next_header_39 : _GEN_2219; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2284 = 3'h4 == encoders_3_io_output ? proc_4_io_next_header_40 : _GEN_2220; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2285 = 3'h4 == encoders_3_io_output ? proc_4_io_next_header_41 : _GEN_2221; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2286 = 3'h4 == encoders_3_io_output ? proc_4_io_next_header_42 : _GEN_2222; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2287 = 3'h4 == encoders_3_io_output ? proc_4_io_next_header_43 : _GEN_2223; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2288 = 3'h4 == encoders_3_io_output ? proc_4_io_next_header_44 : _GEN_2224; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2289 = 3'h4 == encoders_3_io_output ? proc_4_io_next_header_45 : _GEN_2225; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2290 = 3'h4 == encoders_3_io_output ? proc_4_io_next_header_46 : _GEN_2226; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2291 = 3'h4 == encoders_3_io_output ? proc_4_io_next_header_47 : _GEN_2227; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2292 = 3'h4 == encoders_3_io_output ? proc_4_io_next_header_48 : _GEN_2228; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2293 = 3'h4 == encoders_3_io_output ? proc_4_io_next_header_49 : _GEN_2229; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2294 = 3'h4 == encoders_3_io_output ? proc_4_io_next_header_50 : _GEN_2230; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2295 = 3'h4 == encoders_3_io_output ? proc_4_io_next_header_51 : _GEN_2231; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2296 = 3'h4 == encoders_3_io_output ? proc_4_io_next_header_52 : _GEN_2232; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2297 = 3'h4 == encoders_3_io_output ? proc_4_io_next_header_53 : _GEN_2233; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2298 = 3'h4 == encoders_3_io_output ? proc_4_io_next_header_54 : _GEN_2234; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2299 = 3'h4 == encoders_3_io_output ? proc_4_io_next_header_55 : _GEN_2235; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2300 = 3'h4 == encoders_3_io_output ? proc_4_io_next_header_56 : _GEN_2236; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2301 = 3'h4 == encoders_3_io_output ? proc_4_io_next_header_57 : _GEN_2237; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2302 = 3'h4 == encoders_3_io_output ? proc_4_io_next_header_58 : _GEN_2238; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2303 = 3'h4 == encoders_3_io_output ? proc_4_io_next_header_59 : _GEN_2239; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2304 = 3'h4 == encoders_3_io_output ? proc_4_io_next_header_60 : _GEN_2240; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2305 = 3'h4 == encoders_3_io_output ? proc_4_io_next_header_61 : _GEN_2241; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2306 = 3'h4 == encoders_3_io_output ? proc_4_io_next_header_62 : _GEN_2242; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2307 = 3'h4 == encoders_3_io_output ? proc_4_io_next_header_63 : _GEN_2243; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2308 = 3'h5 == encoders_3_io_output ? proc_5_io_next_header_0 : _GEN_2244; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2309 = 3'h5 == encoders_3_io_output ? proc_5_io_next_header_1 : _GEN_2245; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2310 = 3'h5 == encoders_3_io_output ? proc_5_io_next_header_2 : _GEN_2246; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2311 = 3'h5 == encoders_3_io_output ? proc_5_io_next_header_3 : _GEN_2247; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2312 = 3'h5 == encoders_3_io_output ? proc_5_io_next_header_4 : _GEN_2248; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2313 = 3'h5 == encoders_3_io_output ? proc_5_io_next_header_5 : _GEN_2249; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2314 = 3'h5 == encoders_3_io_output ? proc_5_io_next_header_6 : _GEN_2250; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2315 = 3'h5 == encoders_3_io_output ? proc_5_io_next_header_7 : _GEN_2251; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2316 = 3'h5 == encoders_3_io_output ? proc_5_io_next_header_8 : _GEN_2252; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2317 = 3'h5 == encoders_3_io_output ? proc_5_io_next_header_9 : _GEN_2253; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2318 = 3'h5 == encoders_3_io_output ? proc_5_io_next_header_10 : _GEN_2254; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2319 = 3'h5 == encoders_3_io_output ? proc_5_io_next_header_11 : _GEN_2255; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2320 = 3'h5 == encoders_3_io_output ? proc_5_io_next_header_12 : _GEN_2256; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2321 = 3'h5 == encoders_3_io_output ? proc_5_io_next_header_13 : _GEN_2257; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2322 = 3'h5 == encoders_3_io_output ? proc_5_io_next_header_14 : _GEN_2258; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2323 = 3'h5 == encoders_3_io_output ? proc_5_io_next_header_15 : _GEN_2259; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2324 = 3'h5 == encoders_3_io_output ? proc_5_io_next_header_16 : _GEN_2260; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2325 = 3'h5 == encoders_3_io_output ? proc_5_io_next_header_17 : _GEN_2261; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2326 = 3'h5 == encoders_3_io_output ? proc_5_io_next_header_18 : _GEN_2262; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2327 = 3'h5 == encoders_3_io_output ? proc_5_io_next_header_19 : _GEN_2263; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2328 = 3'h5 == encoders_3_io_output ? proc_5_io_next_header_20 : _GEN_2264; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2329 = 3'h5 == encoders_3_io_output ? proc_5_io_next_header_21 : _GEN_2265; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2330 = 3'h5 == encoders_3_io_output ? proc_5_io_next_header_22 : _GEN_2266; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2331 = 3'h5 == encoders_3_io_output ? proc_5_io_next_header_23 : _GEN_2267; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2332 = 3'h5 == encoders_3_io_output ? proc_5_io_next_header_24 : _GEN_2268; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2333 = 3'h5 == encoders_3_io_output ? proc_5_io_next_header_25 : _GEN_2269; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2334 = 3'h5 == encoders_3_io_output ? proc_5_io_next_header_26 : _GEN_2270; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2335 = 3'h5 == encoders_3_io_output ? proc_5_io_next_header_27 : _GEN_2271; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2336 = 3'h5 == encoders_3_io_output ? proc_5_io_next_header_28 : _GEN_2272; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2337 = 3'h5 == encoders_3_io_output ? proc_5_io_next_header_29 : _GEN_2273; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2338 = 3'h5 == encoders_3_io_output ? proc_5_io_next_header_30 : _GEN_2274; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2339 = 3'h5 == encoders_3_io_output ? proc_5_io_next_header_31 : _GEN_2275; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2340 = 3'h5 == encoders_3_io_output ? proc_5_io_next_header_32 : _GEN_2276; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2341 = 3'h5 == encoders_3_io_output ? proc_5_io_next_header_33 : _GEN_2277; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2342 = 3'h5 == encoders_3_io_output ? proc_5_io_next_header_34 : _GEN_2278; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2343 = 3'h5 == encoders_3_io_output ? proc_5_io_next_header_35 : _GEN_2279; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2344 = 3'h5 == encoders_3_io_output ? proc_5_io_next_header_36 : _GEN_2280; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2345 = 3'h5 == encoders_3_io_output ? proc_5_io_next_header_37 : _GEN_2281; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2346 = 3'h5 == encoders_3_io_output ? proc_5_io_next_header_38 : _GEN_2282; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2347 = 3'h5 == encoders_3_io_output ? proc_5_io_next_header_39 : _GEN_2283; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2348 = 3'h5 == encoders_3_io_output ? proc_5_io_next_header_40 : _GEN_2284; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2349 = 3'h5 == encoders_3_io_output ? proc_5_io_next_header_41 : _GEN_2285; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2350 = 3'h5 == encoders_3_io_output ? proc_5_io_next_header_42 : _GEN_2286; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2351 = 3'h5 == encoders_3_io_output ? proc_5_io_next_header_43 : _GEN_2287; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2352 = 3'h5 == encoders_3_io_output ? proc_5_io_next_header_44 : _GEN_2288; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2353 = 3'h5 == encoders_3_io_output ? proc_5_io_next_header_45 : _GEN_2289; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2354 = 3'h5 == encoders_3_io_output ? proc_5_io_next_header_46 : _GEN_2290; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2355 = 3'h5 == encoders_3_io_output ? proc_5_io_next_header_47 : _GEN_2291; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2356 = 3'h5 == encoders_3_io_output ? proc_5_io_next_header_48 : _GEN_2292; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2357 = 3'h5 == encoders_3_io_output ? proc_5_io_next_header_49 : _GEN_2293; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2358 = 3'h5 == encoders_3_io_output ? proc_5_io_next_header_50 : _GEN_2294; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2359 = 3'h5 == encoders_3_io_output ? proc_5_io_next_header_51 : _GEN_2295; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2360 = 3'h5 == encoders_3_io_output ? proc_5_io_next_header_52 : _GEN_2296; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2361 = 3'h5 == encoders_3_io_output ? proc_5_io_next_header_53 : _GEN_2297; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2362 = 3'h5 == encoders_3_io_output ? proc_5_io_next_header_54 : _GEN_2298; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2363 = 3'h5 == encoders_3_io_output ? proc_5_io_next_header_55 : _GEN_2299; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2364 = 3'h5 == encoders_3_io_output ? proc_5_io_next_header_56 : _GEN_2300; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2365 = 3'h5 == encoders_3_io_output ? proc_5_io_next_header_57 : _GEN_2301; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2366 = 3'h5 == encoders_3_io_output ? proc_5_io_next_header_58 : _GEN_2302; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2367 = 3'h5 == encoders_3_io_output ? proc_5_io_next_header_59 : _GEN_2303; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2368 = 3'h5 == encoders_3_io_output ? proc_5_io_next_header_60 : _GEN_2304; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2369 = 3'h5 == encoders_3_io_output ? proc_5_io_next_header_61 : _GEN_2305; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2370 = 3'h5 == encoders_3_io_output ? proc_5_io_next_header_62 : _GEN_2306; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2371 = 3'h5 == encoders_3_io_output ? proc_5_io_next_header_63 : _GEN_2307; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2372 = 3'h6 == encoders_3_io_output ? proc_6_io_next_header_0 : _GEN_2308; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2373 = 3'h6 == encoders_3_io_output ? proc_6_io_next_header_1 : _GEN_2309; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2374 = 3'h6 == encoders_3_io_output ? proc_6_io_next_header_2 : _GEN_2310; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2375 = 3'h6 == encoders_3_io_output ? proc_6_io_next_header_3 : _GEN_2311; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2376 = 3'h6 == encoders_3_io_output ? proc_6_io_next_header_4 : _GEN_2312; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2377 = 3'h6 == encoders_3_io_output ? proc_6_io_next_header_5 : _GEN_2313; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2378 = 3'h6 == encoders_3_io_output ? proc_6_io_next_header_6 : _GEN_2314; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2379 = 3'h6 == encoders_3_io_output ? proc_6_io_next_header_7 : _GEN_2315; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2380 = 3'h6 == encoders_3_io_output ? proc_6_io_next_header_8 : _GEN_2316; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2381 = 3'h6 == encoders_3_io_output ? proc_6_io_next_header_9 : _GEN_2317; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2382 = 3'h6 == encoders_3_io_output ? proc_6_io_next_header_10 : _GEN_2318; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2383 = 3'h6 == encoders_3_io_output ? proc_6_io_next_header_11 : _GEN_2319; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2384 = 3'h6 == encoders_3_io_output ? proc_6_io_next_header_12 : _GEN_2320; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2385 = 3'h6 == encoders_3_io_output ? proc_6_io_next_header_13 : _GEN_2321; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2386 = 3'h6 == encoders_3_io_output ? proc_6_io_next_header_14 : _GEN_2322; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2387 = 3'h6 == encoders_3_io_output ? proc_6_io_next_header_15 : _GEN_2323; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2388 = 3'h6 == encoders_3_io_output ? proc_6_io_next_header_16 : _GEN_2324; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2389 = 3'h6 == encoders_3_io_output ? proc_6_io_next_header_17 : _GEN_2325; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2390 = 3'h6 == encoders_3_io_output ? proc_6_io_next_header_18 : _GEN_2326; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2391 = 3'h6 == encoders_3_io_output ? proc_6_io_next_header_19 : _GEN_2327; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2392 = 3'h6 == encoders_3_io_output ? proc_6_io_next_header_20 : _GEN_2328; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2393 = 3'h6 == encoders_3_io_output ? proc_6_io_next_header_21 : _GEN_2329; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2394 = 3'h6 == encoders_3_io_output ? proc_6_io_next_header_22 : _GEN_2330; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2395 = 3'h6 == encoders_3_io_output ? proc_6_io_next_header_23 : _GEN_2331; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2396 = 3'h6 == encoders_3_io_output ? proc_6_io_next_header_24 : _GEN_2332; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2397 = 3'h6 == encoders_3_io_output ? proc_6_io_next_header_25 : _GEN_2333; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2398 = 3'h6 == encoders_3_io_output ? proc_6_io_next_header_26 : _GEN_2334; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2399 = 3'h6 == encoders_3_io_output ? proc_6_io_next_header_27 : _GEN_2335; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2400 = 3'h6 == encoders_3_io_output ? proc_6_io_next_header_28 : _GEN_2336; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2401 = 3'h6 == encoders_3_io_output ? proc_6_io_next_header_29 : _GEN_2337; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2402 = 3'h6 == encoders_3_io_output ? proc_6_io_next_header_30 : _GEN_2338; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2403 = 3'h6 == encoders_3_io_output ? proc_6_io_next_header_31 : _GEN_2339; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2404 = 3'h6 == encoders_3_io_output ? proc_6_io_next_header_32 : _GEN_2340; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2405 = 3'h6 == encoders_3_io_output ? proc_6_io_next_header_33 : _GEN_2341; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2406 = 3'h6 == encoders_3_io_output ? proc_6_io_next_header_34 : _GEN_2342; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2407 = 3'h6 == encoders_3_io_output ? proc_6_io_next_header_35 : _GEN_2343; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2408 = 3'h6 == encoders_3_io_output ? proc_6_io_next_header_36 : _GEN_2344; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2409 = 3'h6 == encoders_3_io_output ? proc_6_io_next_header_37 : _GEN_2345; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2410 = 3'h6 == encoders_3_io_output ? proc_6_io_next_header_38 : _GEN_2346; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2411 = 3'h6 == encoders_3_io_output ? proc_6_io_next_header_39 : _GEN_2347; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2412 = 3'h6 == encoders_3_io_output ? proc_6_io_next_header_40 : _GEN_2348; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2413 = 3'h6 == encoders_3_io_output ? proc_6_io_next_header_41 : _GEN_2349; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2414 = 3'h6 == encoders_3_io_output ? proc_6_io_next_header_42 : _GEN_2350; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2415 = 3'h6 == encoders_3_io_output ? proc_6_io_next_header_43 : _GEN_2351; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2416 = 3'h6 == encoders_3_io_output ? proc_6_io_next_header_44 : _GEN_2352; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2417 = 3'h6 == encoders_3_io_output ? proc_6_io_next_header_45 : _GEN_2353; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2418 = 3'h6 == encoders_3_io_output ? proc_6_io_next_header_46 : _GEN_2354; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2419 = 3'h6 == encoders_3_io_output ? proc_6_io_next_header_47 : _GEN_2355; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2420 = 3'h6 == encoders_3_io_output ? proc_6_io_next_header_48 : _GEN_2356; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2421 = 3'h6 == encoders_3_io_output ? proc_6_io_next_header_49 : _GEN_2357; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2422 = 3'h6 == encoders_3_io_output ? proc_6_io_next_header_50 : _GEN_2358; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2423 = 3'h6 == encoders_3_io_output ? proc_6_io_next_header_51 : _GEN_2359; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2424 = 3'h6 == encoders_3_io_output ? proc_6_io_next_header_52 : _GEN_2360; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2425 = 3'h6 == encoders_3_io_output ? proc_6_io_next_header_53 : _GEN_2361; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2426 = 3'h6 == encoders_3_io_output ? proc_6_io_next_header_54 : _GEN_2362; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2427 = 3'h6 == encoders_3_io_output ? proc_6_io_next_header_55 : _GEN_2363; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2428 = 3'h6 == encoders_3_io_output ? proc_6_io_next_header_56 : _GEN_2364; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2429 = 3'h6 == encoders_3_io_output ? proc_6_io_next_header_57 : _GEN_2365; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2430 = 3'h6 == encoders_3_io_output ? proc_6_io_next_header_58 : _GEN_2366; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2431 = 3'h6 == encoders_3_io_output ? proc_6_io_next_header_59 : _GEN_2367; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2432 = 3'h6 == encoders_3_io_output ? proc_6_io_next_header_60 : _GEN_2368; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2433 = 3'h6 == encoders_3_io_output ? proc_6_io_next_header_61 : _GEN_2369; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2434 = 3'h6 == encoders_3_io_output ? proc_6_io_next_header_62 : _GEN_2370; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2435 = 3'h6 == encoders_3_io_output ? proc_6_io_next_header_63 : _GEN_2371; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2436 = 3'h7 == encoders_3_io_output ? proc_7_io_next_header_0 : _GEN_2372; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2437 = 3'h7 == encoders_3_io_output ? proc_7_io_next_header_1 : _GEN_2373; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2438 = 3'h7 == encoders_3_io_output ? proc_7_io_next_header_2 : _GEN_2374; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2439 = 3'h7 == encoders_3_io_output ? proc_7_io_next_header_3 : _GEN_2375; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2440 = 3'h7 == encoders_3_io_output ? proc_7_io_next_header_4 : _GEN_2376; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2441 = 3'h7 == encoders_3_io_output ? proc_7_io_next_header_5 : _GEN_2377; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2442 = 3'h7 == encoders_3_io_output ? proc_7_io_next_header_6 : _GEN_2378; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2443 = 3'h7 == encoders_3_io_output ? proc_7_io_next_header_7 : _GEN_2379; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2444 = 3'h7 == encoders_3_io_output ? proc_7_io_next_header_8 : _GEN_2380; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2445 = 3'h7 == encoders_3_io_output ? proc_7_io_next_header_9 : _GEN_2381; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2446 = 3'h7 == encoders_3_io_output ? proc_7_io_next_header_10 : _GEN_2382; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2447 = 3'h7 == encoders_3_io_output ? proc_7_io_next_header_11 : _GEN_2383; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2448 = 3'h7 == encoders_3_io_output ? proc_7_io_next_header_12 : _GEN_2384; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2449 = 3'h7 == encoders_3_io_output ? proc_7_io_next_header_13 : _GEN_2385; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2450 = 3'h7 == encoders_3_io_output ? proc_7_io_next_header_14 : _GEN_2386; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2451 = 3'h7 == encoders_3_io_output ? proc_7_io_next_header_15 : _GEN_2387; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2452 = 3'h7 == encoders_3_io_output ? proc_7_io_next_header_16 : _GEN_2388; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2453 = 3'h7 == encoders_3_io_output ? proc_7_io_next_header_17 : _GEN_2389; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2454 = 3'h7 == encoders_3_io_output ? proc_7_io_next_header_18 : _GEN_2390; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2455 = 3'h7 == encoders_3_io_output ? proc_7_io_next_header_19 : _GEN_2391; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2456 = 3'h7 == encoders_3_io_output ? proc_7_io_next_header_20 : _GEN_2392; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2457 = 3'h7 == encoders_3_io_output ? proc_7_io_next_header_21 : _GEN_2393; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2458 = 3'h7 == encoders_3_io_output ? proc_7_io_next_header_22 : _GEN_2394; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2459 = 3'h7 == encoders_3_io_output ? proc_7_io_next_header_23 : _GEN_2395; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2460 = 3'h7 == encoders_3_io_output ? proc_7_io_next_header_24 : _GEN_2396; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2461 = 3'h7 == encoders_3_io_output ? proc_7_io_next_header_25 : _GEN_2397; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2462 = 3'h7 == encoders_3_io_output ? proc_7_io_next_header_26 : _GEN_2398; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2463 = 3'h7 == encoders_3_io_output ? proc_7_io_next_header_27 : _GEN_2399; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2464 = 3'h7 == encoders_3_io_output ? proc_7_io_next_header_28 : _GEN_2400; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2465 = 3'h7 == encoders_3_io_output ? proc_7_io_next_header_29 : _GEN_2401; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2466 = 3'h7 == encoders_3_io_output ? proc_7_io_next_header_30 : _GEN_2402; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2467 = 3'h7 == encoders_3_io_output ? proc_7_io_next_header_31 : _GEN_2403; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2468 = 3'h7 == encoders_3_io_output ? proc_7_io_next_header_32 : _GEN_2404; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2469 = 3'h7 == encoders_3_io_output ? proc_7_io_next_header_33 : _GEN_2405; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2470 = 3'h7 == encoders_3_io_output ? proc_7_io_next_header_34 : _GEN_2406; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2471 = 3'h7 == encoders_3_io_output ? proc_7_io_next_header_35 : _GEN_2407; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2472 = 3'h7 == encoders_3_io_output ? proc_7_io_next_header_36 : _GEN_2408; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2473 = 3'h7 == encoders_3_io_output ? proc_7_io_next_header_37 : _GEN_2409; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2474 = 3'h7 == encoders_3_io_output ? proc_7_io_next_header_38 : _GEN_2410; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2475 = 3'h7 == encoders_3_io_output ? proc_7_io_next_header_39 : _GEN_2411; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2476 = 3'h7 == encoders_3_io_output ? proc_7_io_next_header_40 : _GEN_2412; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2477 = 3'h7 == encoders_3_io_output ? proc_7_io_next_header_41 : _GEN_2413; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2478 = 3'h7 == encoders_3_io_output ? proc_7_io_next_header_42 : _GEN_2414; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2479 = 3'h7 == encoders_3_io_output ? proc_7_io_next_header_43 : _GEN_2415; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2480 = 3'h7 == encoders_3_io_output ? proc_7_io_next_header_44 : _GEN_2416; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2481 = 3'h7 == encoders_3_io_output ? proc_7_io_next_header_45 : _GEN_2417; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2482 = 3'h7 == encoders_3_io_output ? proc_7_io_next_header_46 : _GEN_2418; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2483 = 3'h7 == encoders_3_io_output ? proc_7_io_next_header_47 : _GEN_2419; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2484 = 3'h7 == encoders_3_io_output ? proc_7_io_next_header_48 : _GEN_2420; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2485 = 3'h7 == encoders_3_io_output ? proc_7_io_next_header_49 : _GEN_2421; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2486 = 3'h7 == encoders_3_io_output ? proc_7_io_next_header_50 : _GEN_2422; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2487 = 3'h7 == encoders_3_io_output ? proc_7_io_next_header_51 : _GEN_2423; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2488 = 3'h7 == encoders_3_io_output ? proc_7_io_next_header_52 : _GEN_2424; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2489 = 3'h7 == encoders_3_io_output ? proc_7_io_next_header_53 : _GEN_2425; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2490 = 3'h7 == encoders_3_io_output ? proc_7_io_next_header_54 : _GEN_2426; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2491 = 3'h7 == encoders_3_io_output ? proc_7_io_next_header_55 : _GEN_2427; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2492 = 3'h7 == encoders_3_io_output ? proc_7_io_next_header_56 : _GEN_2428; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2493 = 3'h7 == encoders_3_io_output ? proc_7_io_next_header_57 : _GEN_2429; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2494 = 3'h7 == encoders_3_io_output ? proc_7_io_next_header_58 : _GEN_2430; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2495 = 3'h7 == encoders_3_io_output ? proc_7_io_next_header_59 : _GEN_2431; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2496 = 3'h7 == encoders_3_io_output ? proc_7_io_next_header_60 : _GEN_2432; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2497 = 3'h7 == encoders_3_io_output ? proc_7_io_next_header_61 : _GEN_2433; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2498 = 3'h7 == encoders_3_io_output ? proc_7_io_next_header_62 : _GEN_2434; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2499 = 3'h7 == encoders_3_io_output ? proc_7_io_next_header_63 : _GEN_2435; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2565 = 3'h0 == encoders_4_io_output ? proc_0_io_next_header_0 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2566 = 3'h0 == encoders_4_io_output ? proc_0_io_next_header_1 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2567 = 3'h0 == encoders_4_io_output ? proc_0_io_next_header_2 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2568 = 3'h0 == encoders_4_io_output ? proc_0_io_next_header_3 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2569 = 3'h0 == encoders_4_io_output ? proc_0_io_next_header_4 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2570 = 3'h0 == encoders_4_io_output ? proc_0_io_next_header_5 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2571 = 3'h0 == encoders_4_io_output ? proc_0_io_next_header_6 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2572 = 3'h0 == encoders_4_io_output ? proc_0_io_next_header_7 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2573 = 3'h0 == encoders_4_io_output ? proc_0_io_next_header_8 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2574 = 3'h0 == encoders_4_io_output ? proc_0_io_next_header_9 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2575 = 3'h0 == encoders_4_io_output ? proc_0_io_next_header_10 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2576 = 3'h0 == encoders_4_io_output ? proc_0_io_next_header_11 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2577 = 3'h0 == encoders_4_io_output ? proc_0_io_next_header_12 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2578 = 3'h0 == encoders_4_io_output ? proc_0_io_next_header_13 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2579 = 3'h0 == encoders_4_io_output ? proc_0_io_next_header_14 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2580 = 3'h0 == encoders_4_io_output ? proc_0_io_next_header_15 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2581 = 3'h0 == encoders_4_io_output ? proc_0_io_next_header_16 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2582 = 3'h0 == encoders_4_io_output ? proc_0_io_next_header_17 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2583 = 3'h0 == encoders_4_io_output ? proc_0_io_next_header_18 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2584 = 3'h0 == encoders_4_io_output ? proc_0_io_next_header_19 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2585 = 3'h0 == encoders_4_io_output ? proc_0_io_next_header_20 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2586 = 3'h0 == encoders_4_io_output ? proc_0_io_next_header_21 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2587 = 3'h0 == encoders_4_io_output ? proc_0_io_next_header_22 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2588 = 3'h0 == encoders_4_io_output ? proc_0_io_next_header_23 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2589 = 3'h0 == encoders_4_io_output ? proc_0_io_next_header_24 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2590 = 3'h0 == encoders_4_io_output ? proc_0_io_next_header_25 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2591 = 3'h0 == encoders_4_io_output ? proc_0_io_next_header_26 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2592 = 3'h0 == encoders_4_io_output ? proc_0_io_next_header_27 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2593 = 3'h0 == encoders_4_io_output ? proc_0_io_next_header_28 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2594 = 3'h0 == encoders_4_io_output ? proc_0_io_next_header_29 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2595 = 3'h0 == encoders_4_io_output ? proc_0_io_next_header_30 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2596 = 3'h0 == encoders_4_io_output ? proc_0_io_next_header_31 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2597 = 3'h0 == encoders_4_io_output ? proc_0_io_next_header_32 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2598 = 3'h0 == encoders_4_io_output ? proc_0_io_next_header_33 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2599 = 3'h0 == encoders_4_io_output ? proc_0_io_next_header_34 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2600 = 3'h0 == encoders_4_io_output ? proc_0_io_next_header_35 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2601 = 3'h0 == encoders_4_io_output ? proc_0_io_next_header_36 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2602 = 3'h0 == encoders_4_io_output ? proc_0_io_next_header_37 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2603 = 3'h0 == encoders_4_io_output ? proc_0_io_next_header_38 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2604 = 3'h0 == encoders_4_io_output ? proc_0_io_next_header_39 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2605 = 3'h0 == encoders_4_io_output ? proc_0_io_next_header_40 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2606 = 3'h0 == encoders_4_io_output ? proc_0_io_next_header_41 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2607 = 3'h0 == encoders_4_io_output ? proc_0_io_next_header_42 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2608 = 3'h0 == encoders_4_io_output ? proc_0_io_next_header_43 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2609 = 3'h0 == encoders_4_io_output ? proc_0_io_next_header_44 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2610 = 3'h0 == encoders_4_io_output ? proc_0_io_next_header_45 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2611 = 3'h0 == encoders_4_io_output ? proc_0_io_next_header_46 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2612 = 3'h0 == encoders_4_io_output ? proc_0_io_next_header_47 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2613 = 3'h0 == encoders_4_io_output ? proc_0_io_next_header_48 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2614 = 3'h0 == encoders_4_io_output ? proc_0_io_next_header_49 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2615 = 3'h0 == encoders_4_io_output ? proc_0_io_next_header_50 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2616 = 3'h0 == encoders_4_io_output ? proc_0_io_next_header_51 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2617 = 3'h0 == encoders_4_io_output ? proc_0_io_next_header_52 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2618 = 3'h0 == encoders_4_io_output ? proc_0_io_next_header_53 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2619 = 3'h0 == encoders_4_io_output ? proc_0_io_next_header_54 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2620 = 3'h0 == encoders_4_io_output ? proc_0_io_next_header_55 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2621 = 3'h0 == encoders_4_io_output ? proc_0_io_next_header_56 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2622 = 3'h0 == encoders_4_io_output ? proc_0_io_next_header_57 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2623 = 3'h0 == encoders_4_io_output ? proc_0_io_next_header_58 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2624 = 3'h0 == encoders_4_io_output ? proc_0_io_next_header_59 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2625 = 3'h0 == encoders_4_io_output ? proc_0_io_next_header_60 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2626 = 3'h0 == encoders_4_io_output ? proc_0_io_next_header_61 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2627 = 3'h0 == encoders_4_io_output ? proc_0_io_next_header_62 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2628 = 3'h0 == encoders_4_io_output ? proc_0_io_next_header_63 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_2629 = 3'h1 == encoders_4_io_output ? proc_1_io_next_header_0 : _GEN_2565; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2630 = 3'h1 == encoders_4_io_output ? proc_1_io_next_header_1 : _GEN_2566; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2631 = 3'h1 == encoders_4_io_output ? proc_1_io_next_header_2 : _GEN_2567; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2632 = 3'h1 == encoders_4_io_output ? proc_1_io_next_header_3 : _GEN_2568; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2633 = 3'h1 == encoders_4_io_output ? proc_1_io_next_header_4 : _GEN_2569; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2634 = 3'h1 == encoders_4_io_output ? proc_1_io_next_header_5 : _GEN_2570; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2635 = 3'h1 == encoders_4_io_output ? proc_1_io_next_header_6 : _GEN_2571; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2636 = 3'h1 == encoders_4_io_output ? proc_1_io_next_header_7 : _GEN_2572; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2637 = 3'h1 == encoders_4_io_output ? proc_1_io_next_header_8 : _GEN_2573; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2638 = 3'h1 == encoders_4_io_output ? proc_1_io_next_header_9 : _GEN_2574; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2639 = 3'h1 == encoders_4_io_output ? proc_1_io_next_header_10 : _GEN_2575; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2640 = 3'h1 == encoders_4_io_output ? proc_1_io_next_header_11 : _GEN_2576; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2641 = 3'h1 == encoders_4_io_output ? proc_1_io_next_header_12 : _GEN_2577; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2642 = 3'h1 == encoders_4_io_output ? proc_1_io_next_header_13 : _GEN_2578; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2643 = 3'h1 == encoders_4_io_output ? proc_1_io_next_header_14 : _GEN_2579; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2644 = 3'h1 == encoders_4_io_output ? proc_1_io_next_header_15 : _GEN_2580; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2645 = 3'h1 == encoders_4_io_output ? proc_1_io_next_header_16 : _GEN_2581; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2646 = 3'h1 == encoders_4_io_output ? proc_1_io_next_header_17 : _GEN_2582; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2647 = 3'h1 == encoders_4_io_output ? proc_1_io_next_header_18 : _GEN_2583; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2648 = 3'h1 == encoders_4_io_output ? proc_1_io_next_header_19 : _GEN_2584; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2649 = 3'h1 == encoders_4_io_output ? proc_1_io_next_header_20 : _GEN_2585; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2650 = 3'h1 == encoders_4_io_output ? proc_1_io_next_header_21 : _GEN_2586; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2651 = 3'h1 == encoders_4_io_output ? proc_1_io_next_header_22 : _GEN_2587; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2652 = 3'h1 == encoders_4_io_output ? proc_1_io_next_header_23 : _GEN_2588; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2653 = 3'h1 == encoders_4_io_output ? proc_1_io_next_header_24 : _GEN_2589; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2654 = 3'h1 == encoders_4_io_output ? proc_1_io_next_header_25 : _GEN_2590; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2655 = 3'h1 == encoders_4_io_output ? proc_1_io_next_header_26 : _GEN_2591; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2656 = 3'h1 == encoders_4_io_output ? proc_1_io_next_header_27 : _GEN_2592; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2657 = 3'h1 == encoders_4_io_output ? proc_1_io_next_header_28 : _GEN_2593; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2658 = 3'h1 == encoders_4_io_output ? proc_1_io_next_header_29 : _GEN_2594; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2659 = 3'h1 == encoders_4_io_output ? proc_1_io_next_header_30 : _GEN_2595; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2660 = 3'h1 == encoders_4_io_output ? proc_1_io_next_header_31 : _GEN_2596; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2661 = 3'h1 == encoders_4_io_output ? proc_1_io_next_header_32 : _GEN_2597; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2662 = 3'h1 == encoders_4_io_output ? proc_1_io_next_header_33 : _GEN_2598; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2663 = 3'h1 == encoders_4_io_output ? proc_1_io_next_header_34 : _GEN_2599; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2664 = 3'h1 == encoders_4_io_output ? proc_1_io_next_header_35 : _GEN_2600; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2665 = 3'h1 == encoders_4_io_output ? proc_1_io_next_header_36 : _GEN_2601; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2666 = 3'h1 == encoders_4_io_output ? proc_1_io_next_header_37 : _GEN_2602; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2667 = 3'h1 == encoders_4_io_output ? proc_1_io_next_header_38 : _GEN_2603; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2668 = 3'h1 == encoders_4_io_output ? proc_1_io_next_header_39 : _GEN_2604; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2669 = 3'h1 == encoders_4_io_output ? proc_1_io_next_header_40 : _GEN_2605; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2670 = 3'h1 == encoders_4_io_output ? proc_1_io_next_header_41 : _GEN_2606; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2671 = 3'h1 == encoders_4_io_output ? proc_1_io_next_header_42 : _GEN_2607; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2672 = 3'h1 == encoders_4_io_output ? proc_1_io_next_header_43 : _GEN_2608; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2673 = 3'h1 == encoders_4_io_output ? proc_1_io_next_header_44 : _GEN_2609; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2674 = 3'h1 == encoders_4_io_output ? proc_1_io_next_header_45 : _GEN_2610; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2675 = 3'h1 == encoders_4_io_output ? proc_1_io_next_header_46 : _GEN_2611; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2676 = 3'h1 == encoders_4_io_output ? proc_1_io_next_header_47 : _GEN_2612; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2677 = 3'h1 == encoders_4_io_output ? proc_1_io_next_header_48 : _GEN_2613; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2678 = 3'h1 == encoders_4_io_output ? proc_1_io_next_header_49 : _GEN_2614; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2679 = 3'h1 == encoders_4_io_output ? proc_1_io_next_header_50 : _GEN_2615; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2680 = 3'h1 == encoders_4_io_output ? proc_1_io_next_header_51 : _GEN_2616; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2681 = 3'h1 == encoders_4_io_output ? proc_1_io_next_header_52 : _GEN_2617; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2682 = 3'h1 == encoders_4_io_output ? proc_1_io_next_header_53 : _GEN_2618; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2683 = 3'h1 == encoders_4_io_output ? proc_1_io_next_header_54 : _GEN_2619; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2684 = 3'h1 == encoders_4_io_output ? proc_1_io_next_header_55 : _GEN_2620; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2685 = 3'h1 == encoders_4_io_output ? proc_1_io_next_header_56 : _GEN_2621; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2686 = 3'h1 == encoders_4_io_output ? proc_1_io_next_header_57 : _GEN_2622; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2687 = 3'h1 == encoders_4_io_output ? proc_1_io_next_header_58 : _GEN_2623; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2688 = 3'h1 == encoders_4_io_output ? proc_1_io_next_header_59 : _GEN_2624; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2689 = 3'h1 == encoders_4_io_output ? proc_1_io_next_header_60 : _GEN_2625; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2690 = 3'h1 == encoders_4_io_output ? proc_1_io_next_header_61 : _GEN_2626; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2691 = 3'h1 == encoders_4_io_output ? proc_1_io_next_header_62 : _GEN_2627; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2692 = 3'h1 == encoders_4_io_output ? proc_1_io_next_header_63 : _GEN_2628; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2693 = 3'h2 == encoders_4_io_output ? proc_2_io_next_header_0 : _GEN_2629; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2694 = 3'h2 == encoders_4_io_output ? proc_2_io_next_header_1 : _GEN_2630; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2695 = 3'h2 == encoders_4_io_output ? proc_2_io_next_header_2 : _GEN_2631; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2696 = 3'h2 == encoders_4_io_output ? proc_2_io_next_header_3 : _GEN_2632; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2697 = 3'h2 == encoders_4_io_output ? proc_2_io_next_header_4 : _GEN_2633; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2698 = 3'h2 == encoders_4_io_output ? proc_2_io_next_header_5 : _GEN_2634; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2699 = 3'h2 == encoders_4_io_output ? proc_2_io_next_header_6 : _GEN_2635; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2700 = 3'h2 == encoders_4_io_output ? proc_2_io_next_header_7 : _GEN_2636; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2701 = 3'h2 == encoders_4_io_output ? proc_2_io_next_header_8 : _GEN_2637; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2702 = 3'h2 == encoders_4_io_output ? proc_2_io_next_header_9 : _GEN_2638; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2703 = 3'h2 == encoders_4_io_output ? proc_2_io_next_header_10 : _GEN_2639; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2704 = 3'h2 == encoders_4_io_output ? proc_2_io_next_header_11 : _GEN_2640; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2705 = 3'h2 == encoders_4_io_output ? proc_2_io_next_header_12 : _GEN_2641; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2706 = 3'h2 == encoders_4_io_output ? proc_2_io_next_header_13 : _GEN_2642; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2707 = 3'h2 == encoders_4_io_output ? proc_2_io_next_header_14 : _GEN_2643; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2708 = 3'h2 == encoders_4_io_output ? proc_2_io_next_header_15 : _GEN_2644; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2709 = 3'h2 == encoders_4_io_output ? proc_2_io_next_header_16 : _GEN_2645; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2710 = 3'h2 == encoders_4_io_output ? proc_2_io_next_header_17 : _GEN_2646; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2711 = 3'h2 == encoders_4_io_output ? proc_2_io_next_header_18 : _GEN_2647; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2712 = 3'h2 == encoders_4_io_output ? proc_2_io_next_header_19 : _GEN_2648; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2713 = 3'h2 == encoders_4_io_output ? proc_2_io_next_header_20 : _GEN_2649; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2714 = 3'h2 == encoders_4_io_output ? proc_2_io_next_header_21 : _GEN_2650; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2715 = 3'h2 == encoders_4_io_output ? proc_2_io_next_header_22 : _GEN_2651; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2716 = 3'h2 == encoders_4_io_output ? proc_2_io_next_header_23 : _GEN_2652; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2717 = 3'h2 == encoders_4_io_output ? proc_2_io_next_header_24 : _GEN_2653; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2718 = 3'h2 == encoders_4_io_output ? proc_2_io_next_header_25 : _GEN_2654; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2719 = 3'h2 == encoders_4_io_output ? proc_2_io_next_header_26 : _GEN_2655; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2720 = 3'h2 == encoders_4_io_output ? proc_2_io_next_header_27 : _GEN_2656; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2721 = 3'h2 == encoders_4_io_output ? proc_2_io_next_header_28 : _GEN_2657; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2722 = 3'h2 == encoders_4_io_output ? proc_2_io_next_header_29 : _GEN_2658; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2723 = 3'h2 == encoders_4_io_output ? proc_2_io_next_header_30 : _GEN_2659; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2724 = 3'h2 == encoders_4_io_output ? proc_2_io_next_header_31 : _GEN_2660; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2725 = 3'h2 == encoders_4_io_output ? proc_2_io_next_header_32 : _GEN_2661; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2726 = 3'h2 == encoders_4_io_output ? proc_2_io_next_header_33 : _GEN_2662; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2727 = 3'h2 == encoders_4_io_output ? proc_2_io_next_header_34 : _GEN_2663; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2728 = 3'h2 == encoders_4_io_output ? proc_2_io_next_header_35 : _GEN_2664; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2729 = 3'h2 == encoders_4_io_output ? proc_2_io_next_header_36 : _GEN_2665; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2730 = 3'h2 == encoders_4_io_output ? proc_2_io_next_header_37 : _GEN_2666; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2731 = 3'h2 == encoders_4_io_output ? proc_2_io_next_header_38 : _GEN_2667; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2732 = 3'h2 == encoders_4_io_output ? proc_2_io_next_header_39 : _GEN_2668; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2733 = 3'h2 == encoders_4_io_output ? proc_2_io_next_header_40 : _GEN_2669; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2734 = 3'h2 == encoders_4_io_output ? proc_2_io_next_header_41 : _GEN_2670; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2735 = 3'h2 == encoders_4_io_output ? proc_2_io_next_header_42 : _GEN_2671; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2736 = 3'h2 == encoders_4_io_output ? proc_2_io_next_header_43 : _GEN_2672; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2737 = 3'h2 == encoders_4_io_output ? proc_2_io_next_header_44 : _GEN_2673; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2738 = 3'h2 == encoders_4_io_output ? proc_2_io_next_header_45 : _GEN_2674; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2739 = 3'h2 == encoders_4_io_output ? proc_2_io_next_header_46 : _GEN_2675; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2740 = 3'h2 == encoders_4_io_output ? proc_2_io_next_header_47 : _GEN_2676; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2741 = 3'h2 == encoders_4_io_output ? proc_2_io_next_header_48 : _GEN_2677; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2742 = 3'h2 == encoders_4_io_output ? proc_2_io_next_header_49 : _GEN_2678; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2743 = 3'h2 == encoders_4_io_output ? proc_2_io_next_header_50 : _GEN_2679; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2744 = 3'h2 == encoders_4_io_output ? proc_2_io_next_header_51 : _GEN_2680; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2745 = 3'h2 == encoders_4_io_output ? proc_2_io_next_header_52 : _GEN_2681; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2746 = 3'h2 == encoders_4_io_output ? proc_2_io_next_header_53 : _GEN_2682; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2747 = 3'h2 == encoders_4_io_output ? proc_2_io_next_header_54 : _GEN_2683; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2748 = 3'h2 == encoders_4_io_output ? proc_2_io_next_header_55 : _GEN_2684; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2749 = 3'h2 == encoders_4_io_output ? proc_2_io_next_header_56 : _GEN_2685; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2750 = 3'h2 == encoders_4_io_output ? proc_2_io_next_header_57 : _GEN_2686; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2751 = 3'h2 == encoders_4_io_output ? proc_2_io_next_header_58 : _GEN_2687; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2752 = 3'h2 == encoders_4_io_output ? proc_2_io_next_header_59 : _GEN_2688; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2753 = 3'h2 == encoders_4_io_output ? proc_2_io_next_header_60 : _GEN_2689; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2754 = 3'h2 == encoders_4_io_output ? proc_2_io_next_header_61 : _GEN_2690; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2755 = 3'h2 == encoders_4_io_output ? proc_2_io_next_header_62 : _GEN_2691; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2756 = 3'h2 == encoders_4_io_output ? proc_2_io_next_header_63 : _GEN_2692; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2757 = 3'h3 == encoders_4_io_output ? proc_3_io_next_header_0 : _GEN_2693; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2758 = 3'h3 == encoders_4_io_output ? proc_3_io_next_header_1 : _GEN_2694; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2759 = 3'h3 == encoders_4_io_output ? proc_3_io_next_header_2 : _GEN_2695; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2760 = 3'h3 == encoders_4_io_output ? proc_3_io_next_header_3 : _GEN_2696; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2761 = 3'h3 == encoders_4_io_output ? proc_3_io_next_header_4 : _GEN_2697; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2762 = 3'h3 == encoders_4_io_output ? proc_3_io_next_header_5 : _GEN_2698; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2763 = 3'h3 == encoders_4_io_output ? proc_3_io_next_header_6 : _GEN_2699; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2764 = 3'h3 == encoders_4_io_output ? proc_3_io_next_header_7 : _GEN_2700; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2765 = 3'h3 == encoders_4_io_output ? proc_3_io_next_header_8 : _GEN_2701; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2766 = 3'h3 == encoders_4_io_output ? proc_3_io_next_header_9 : _GEN_2702; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2767 = 3'h3 == encoders_4_io_output ? proc_3_io_next_header_10 : _GEN_2703; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2768 = 3'h3 == encoders_4_io_output ? proc_3_io_next_header_11 : _GEN_2704; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2769 = 3'h3 == encoders_4_io_output ? proc_3_io_next_header_12 : _GEN_2705; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2770 = 3'h3 == encoders_4_io_output ? proc_3_io_next_header_13 : _GEN_2706; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2771 = 3'h3 == encoders_4_io_output ? proc_3_io_next_header_14 : _GEN_2707; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2772 = 3'h3 == encoders_4_io_output ? proc_3_io_next_header_15 : _GEN_2708; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2773 = 3'h3 == encoders_4_io_output ? proc_3_io_next_header_16 : _GEN_2709; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2774 = 3'h3 == encoders_4_io_output ? proc_3_io_next_header_17 : _GEN_2710; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2775 = 3'h3 == encoders_4_io_output ? proc_3_io_next_header_18 : _GEN_2711; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2776 = 3'h3 == encoders_4_io_output ? proc_3_io_next_header_19 : _GEN_2712; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2777 = 3'h3 == encoders_4_io_output ? proc_3_io_next_header_20 : _GEN_2713; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2778 = 3'h3 == encoders_4_io_output ? proc_3_io_next_header_21 : _GEN_2714; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2779 = 3'h3 == encoders_4_io_output ? proc_3_io_next_header_22 : _GEN_2715; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2780 = 3'h3 == encoders_4_io_output ? proc_3_io_next_header_23 : _GEN_2716; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2781 = 3'h3 == encoders_4_io_output ? proc_3_io_next_header_24 : _GEN_2717; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2782 = 3'h3 == encoders_4_io_output ? proc_3_io_next_header_25 : _GEN_2718; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2783 = 3'h3 == encoders_4_io_output ? proc_3_io_next_header_26 : _GEN_2719; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2784 = 3'h3 == encoders_4_io_output ? proc_3_io_next_header_27 : _GEN_2720; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2785 = 3'h3 == encoders_4_io_output ? proc_3_io_next_header_28 : _GEN_2721; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2786 = 3'h3 == encoders_4_io_output ? proc_3_io_next_header_29 : _GEN_2722; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2787 = 3'h3 == encoders_4_io_output ? proc_3_io_next_header_30 : _GEN_2723; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2788 = 3'h3 == encoders_4_io_output ? proc_3_io_next_header_31 : _GEN_2724; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2789 = 3'h3 == encoders_4_io_output ? proc_3_io_next_header_32 : _GEN_2725; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2790 = 3'h3 == encoders_4_io_output ? proc_3_io_next_header_33 : _GEN_2726; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2791 = 3'h3 == encoders_4_io_output ? proc_3_io_next_header_34 : _GEN_2727; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2792 = 3'h3 == encoders_4_io_output ? proc_3_io_next_header_35 : _GEN_2728; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2793 = 3'h3 == encoders_4_io_output ? proc_3_io_next_header_36 : _GEN_2729; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2794 = 3'h3 == encoders_4_io_output ? proc_3_io_next_header_37 : _GEN_2730; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2795 = 3'h3 == encoders_4_io_output ? proc_3_io_next_header_38 : _GEN_2731; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2796 = 3'h3 == encoders_4_io_output ? proc_3_io_next_header_39 : _GEN_2732; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2797 = 3'h3 == encoders_4_io_output ? proc_3_io_next_header_40 : _GEN_2733; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2798 = 3'h3 == encoders_4_io_output ? proc_3_io_next_header_41 : _GEN_2734; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2799 = 3'h3 == encoders_4_io_output ? proc_3_io_next_header_42 : _GEN_2735; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2800 = 3'h3 == encoders_4_io_output ? proc_3_io_next_header_43 : _GEN_2736; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2801 = 3'h3 == encoders_4_io_output ? proc_3_io_next_header_44 : _GEN_2737; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2802 = 3'h3 == encoders_4_io_output ? proc_3_io_next_header_45 : _GEN_2738; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2803 = 3'h3 == encoders_4_io_output ? proc_3_io_next_header_46 : _GEN_2739; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2804 = 3'h3 == encoders_4_io_output ? proc_3_io_next_header_47 : _GEN_2740; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2805 = 3'h3 == encoders_4_io_output ? proc_3_io_next_header_48 : _GEN_2741; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2806 = 3'h3 == encoders_4_io_output ? proc_3_io_next_header_49 : _GEN_2742; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2807 = 3'h3 == encoders_4_io_output ? proc_3_io_next_header_50 : _GEN_2743; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2808 = 3'h3 == encoders_4_io_output ? proc_3_io_next_header_51 : _GEN_2744; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2809 = 3'h3 == encoders_4_io_output ? proc_3_io_next_header_52 : _GEN_2745; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2810 = 3'h3 == encoders_4_io_output ? proc_3_io_next_header_53 : _GEN_2746; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2811 = 3'h3 == encoders_4_io_output ? proc_3_io_next_header_54 : _GEN_2747; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2812 = 3'h3 == encoders_4_io_output ? proc_3_io_next_header_55 : _GEN_2748; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2813 = 3'h3 == encoders_4_io_output ? proc_3_io_next_header_56 : _GEN_2749; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2814 = 3'h3 == encoders_4_io_output ? proc_3_io_next_header_57 : _GEN_2750; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2815 = 3'h3 == encoders_4_io_output ? proc_3_io_next_header_58 : _GEN_2751; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2816 = 3'h3 == encoders_4_io_output ? proc_3_io_next_header_59 : _GEN_2752; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2817 = 3'h3 == encoders_4_io_output ? proc_3_io_next_header_60 : _GEN_2753; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2818 = 3'h3 == encoders_4_io_output ? proc_3_io_next_header_61 : _GEN_2754; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2819 = 3'h3 == encoders_4_io_output ? proc_3_io_next_header_62 : _GEN_2755; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2820 = 3'h3 == encoders_4_io_output ? proc_3_io_next_header_63 : _GEN_2756; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2821 = 3'h4 == encoders_4_io_output ? proc_4_io_next_header_0 : _GEN_2757; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2822 = 3'h4 == encoders_4_io_output ? proc_4_io_next_header_1 : _GEN_2758; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2823 = 3'h4 == encoders_4_io_output ? proc_4_io_next_header_2 : _GEN_2759; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2824 = 3'h4 == encoders_4_io_output ? proc_4_io_next_header_3 : _GEN_2760; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2825 = 3'h4 == encoders_4_io_output ? proc_4_io_next_header_4 : _GEN_2761; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2826 = 3'h4 == encoders_4_io_output ? proc_4_io_next_header_5 : _GEN_2762; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2827 = 3'h4 == encoders_4_io_output ? proc_4_io_next_header_6 : _GEN_2763; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2828 = 3'h4 == encoders_4_io_output ? proc_4_io_next_header_7 : _GEN_2764; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2829 = 3'h4 == encoders_4_io_output ? proc_4_io_next_header_8 : _GEN_2765; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2830 = 3'h4 == encoders_4_io_output ? proc_4_io_next_header_9 : _GEN_2766; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2831 = 3'h4 == encoders_4_io_output ? proc_4_io_next_header_10 : _GEN_2767; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2832 = 3'h4 == encoders_4_io_output ? proc_4_io_next_header_11 : _GEN_2768; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2833 = 3'h4 == encoders_4_io_output ? proc_4_io_next_header_12 : _GEN_2769; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2834 = 3'h4 == encoders_4_io_output ? proc_4_io_next_header_13 : _GEN_2770; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2835 = 3'h4 == encoders_4_io_output ? proc_4_io_next_header_14 : _GEN_2771; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2836 = 3'h4 == encoders_4_io_output ? proc_4_io_next_header_15 : _GEN_2772; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2837 = 3'h4 == encoders_4_io_output ? proc_4_io_next_header_16 : _GEN_2773; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2838 = 3'h4 == encoders_4_io_output ? proc_4_io_next_header_17 : _GEN_2774; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2839 = 3'h4 == encoders_4_io_output ? proc_4_io_next_header_18 : _GEN_2775; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2840 = 3'h4 == encoders_4_io_output ? proc_4_io_next_header_19 : _GEN_2776; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2841 = 3'h4 == encoders_4_io_output ? proc_4_io_next_header_20 : _GEN_2777; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2842 = 3'h4 == encoders_4_io_output ? proc_4_io_next_header_21 : _GEN_2778; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2843 = 3'h4 == encoders_4_io_output ? proc_4_io_next_header_22 : _GEN_2779; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2844 = 3'h4 == encoders_4_io_output ? proc_4_io_next_header_23 : _GEN_2780; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2845 = 3'h4 == encoders_4_io_output ? proc_4_io_next_header_24 : _GEN_2781; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2846 = 3'h4 == encoders_4_io_output ? proc_4_io_next_header_25 : _GEN_2782; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2847 = 3'h4 == encoders_4_io_output ? proc_4_io_next_header_26 : _GEN_2783; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2848 = 3'h4 == encoders_4_io_output ? proc_4_io_next_header_27 : _GEN_2784; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2849 = 3'h4 == encoders_4_io_output ? proc_4_io_next_header_28 : _GEN_2785; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2850 = 3'h4 == encoders_4_io_output ? proc_4_io_next_header_29 : _GEN_2786; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2851 = 3'h4 == encoders_4_io_output ? proc_4_io_next_header_30 : _GEN_2787; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2852 = 3'h4 == encoders_4_io_output ? proc_4_io_next_header_31 : _GEN_2788; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2853 = 3'h4 == encoders_4_io_output ? proc_4_io_next_header_32 : _GEN_2789; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2854 = 3'h4 == encoders_4_io_output ? proc_4_io_next_header_33 : _GEN_2790; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2855 = 3'h4 == encoders_4_io_output ? proc_4_io_next_header_34 : _GEN_2791; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2856 = 3'h4 == encoders_4_io_output ? proc_4_io_next_header_35 : _GEN_2792; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2857 = 3'h4 == encoders_4_io_output ? proc_4_io_next_header_36 : _GEN_2793; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2858 = 3'h4 == encoders_4_io_output ? proc_4_io_next_header_37 : _GEN_2794; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2859 = 3'h4 == encoders_4_io_output ? proc_4_io_next_header_38 : _GEN_2795; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2860 = 3'h4 == encoders_4_io_output ? proc_4_io_next_header_39 : _GEN_2796; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2861 = 3'h4 == encoders_4_io_output ? proc_4_io_next_header_40 : _GEN_2797; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2862 = 3'h4 == encoders_4_io_output ? proc_4_io_next_header_41 : _GEN_2798; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2863 = 3'h4 == encoders_4_io_output ? proc_4_io_next_header_42 : _GEN_2799; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2864 = 3'h4 == encoders_4_io_output ? proc_4_io_next_header_43 : _GEN_2800; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2865 = 3'h4 == encoders_4_io_output ? proc_4_io_next_header_44 : _GEN_2801; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2866 = 3'h4 == encoders_4_io_output ? proc_4_io_next_header_45 : _GEN_2802; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2867 = 3'h4 == encoders_4_io_output ? proc_4_io_next_header_46 : _GEN_2803; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2868 = 3'h4 == encoders_4_io_output ? proc_4_io_next_header_47 : _GEN_2804; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2869 = 3'h4 == encoders_4_io_output ? proc_4_io_next_header_48 : _GEN_2805; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2870 = 3'h4 == encoders_4_io_output ? proc_4_io_next_header_49 : _GEN_2806; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2871 = 3'h4 == encoders_4_io_output ? proc_4_io_next_header_50 : _GEN_2807; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2872 = 3'h4 == encoders_4_io_output ? proc_4_io_next_header_51 : _GEN_2808; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2873 = 3'h4 == encoders_4_io_output ? proc_4_io_next_header_52 : _GEN_2809; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2874 = 3'h4 == encoders_4_io_output ? proc_4_io_next_header_53 : _GEN_2810; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2875 = 3'h4 == encoders_4_io_output ? proc_4_io_next_header_54 : _GEN_2811; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2876 = 3'h4 == encoders_4_io_output ? proc_4_io_next_header_55 : _GEN_2812; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2877 = 3'h4 == encoders_4_io_output ? proc_4_io_next_header_56 : _GEN_2813; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2878 = 3'h4 == encoders_4_io_output ? proc_4_io_next_header_57 : _GEN_2814; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2879 = 3'h4 == encoders_4_io_output ? proc_4_io_next_header_58 : _GEN_2815; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2880 = 3'h4 == encoders_4_io_output ? proc_4_io_next_header_59 : _GEN_2816; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2881 = 3'h4 == encoders_4_io_output ? proc_4_io_next_header_60 : _GEN_2817; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2882 = 3'h4 == encoders_4_io_output ? proc_4_io_next_header_61 : _GEN_2818; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2883 = 3'h4 == encoders_4_io_output ? proc_4_io_next_header_62 : _GEN_2819; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2884 = 3'h4 == encoders_4_io_output ? proc_4_io_next_header_63 : _GEN_2820; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2885 = 3'h5 == encoders_4_io_output ? proc_5_io_next_header_0 : _GEN_2821; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2886 = 3'h5 == encoders_4_io_output ? proc_5_io_next_header_1 : _GEN_2822; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2887 = 3'h5 == encoders_4_io_output ? proc_5_io_next_header_2 : _GEN_2823; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2888 = 3'h5 == encoders_4_io_output ? proc_5_io_next_header_3 : _GEN_2824; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2889 = 3'h5 == encoders_4_io_output ? proc_5_io_next_header_4 : _GEN_2825; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2890 = 3'h5 == encoders_4_io_output ? proc_5_io_next_header_5 : _GEN_2826; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2891 = 3'h5 == encoders_4_io_output ? proc_5_io_next_header_6 : _GEN_2827; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2892 = 3'h5 == encoders_4_io_output ? proc_5_io_next_header_7 : _GEN_2828; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2893 = 3'h5 == encoders_4_io_output ? proc_5_io_next_header_8 : _GEN_2829; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2894 = 3'h5 == encoders_4_io_output ? proc_5_io_next_header_9 : _GEN_2830; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2895 = 3'h5 == encoders_4_io_output ? proc_5_io_next_header_10 : _GEN_2831; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2896 = 3'h5 == encoders_4_io_output ? proc_5_io_next_header_11 : _GEN_2832; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2897 = 3'h5 == encoders_4_io_output ? proc_5_io_next_header_12 : _GEN_2833; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2898 = 3'h5 == encoders_4_io_output ? proc_5_io_next_header_13 : _GEN_2834; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2899 = 3'h5 == encoders_4_io_output ? proc_5_io_next_header_14 : _GEN_2835; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2900 = 3'h5 == encoders_4_io_output ? proc_5_io_next_header_15 : _GEN_2836; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2901 = 3'h5 == encoders_4_io_output ? proc_5_io_next_header_16 : _GEN_2837; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2902 = 3'h5 == encoders_4_io_output ? proc_5_io_next_header_17 : _GEN_2838; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2903 = 3'h5 == encoders_4_io_output ? proc_5_io_next_header_18 : _GEN_2839; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2904 = 3'h5 == encoders_4_io_output ? proc_5_io_next_header_19 : _GEN_2840; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2905 = 3'h5 == encoders_4_io_output ? proc_5_io_next_header_20 : _GEN_2841; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2906 = 3'h5 == encoders_4_io_output ? proc_5_io_next_header_21 : _GEN_2842; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2907 = 3'h5 == encoders_4_io_output ? proc_5_io_next_header_22 : _GEN_2843; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2908 = 3'h5 == encoders_4_io_output ? proc_5_io_next_header_23 : _GEN_2844; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2909 = 3'h5 == encoders_4_io_output ? proc_5_io_next_header_24 : _GEN_2845; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2910 = 3'h5 == encoders_4_io_output ? proc_5_io_next_header_25 : _GEN_2846; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2911 = 3'h5 == encoders_4_io_output ? proc_5_io_next_header_26 : _GEN_2847; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2912 = 3'h5 == encoders_4_io_output ? proc_5_io_next_header_27 : _GEN_2848; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2913 = 3'h5 == encoders_4_io_output ? proc_5_io_next_header_28 : _GEN_2849; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2914 = 3'h5 == encoders_4_io_output ? proc_5_io_next_header_29 : _GEN_2850; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2915 = 3'h5 == encoders_4_io_output ? proc_5_io_next_header_30 : _GEN_2851; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2916 = 3'h5 == encoders_4_io_output ? proc_5_io_next_header_31 : _GEN_2852; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2917 = 3'h5 == encoders_4_io_output ? proc_5_io_next_header_32 : _GEN_2853; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2918 = 3'h5 == encoders_4_io_output ? proc_5_io_next_header_33 : _GEN_2854; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2919 = 3'h5 == encoders_4_io_output ? proc_5_io_next_header_34 : _GEN_2855; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2920 = 3'h5 == encoders_4_io_output ? proc_5_io_next_header_35 : _GEN_2856; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2921 = 3'h5 == encoders_4_io_output ? proc_5_io_next_header_36 : _GEN_2857; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2922 = 3'h5 == encoders_4_io_output ? proc_5_io_next_header_37 : _GEN_2858; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2923 = 3'h5 == encoders_4_io_output ? proc_5_io_next_header_38 : _GEN_2859; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2924 = 3'h5 == encoders_4_io_output ? proc_5_io_next_header_39 : _GEN_2860; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2925 = 3'h5 == encoders_4_io_output ? proc_5_io_next_header_40 : _GEN_2861; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2926 = 3'h5 == encoders_4_io_output ? proc_5_io_next_header_41 : _GEN_2862; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2927 = 3'h5 == encoders_4_io_output ? proc_5_io_next_header_42 : _GEN_2863; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2928 = 3'h5 == encoders_4_io_output ? proc_5_io_next_header_43 : _GEN_2864; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2929 = 3'h5 == encoders_4_io_output ? proc_5_io_next_header_44 : _GEN_2865; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2930 = 3'h5 == encoders_4_io_output ? proc_5_io_next_header_45 : _GEN_2866; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2931 = 3'h5 == encoders_4_io_output ? proc_5_io_next_header_46 : _GEN_2867; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2932 = 3'h5 == encoders_4_io_output ? proc_5_io_next_header_47 : _GEN_2868; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2933 = 3'h5 == encoders_4_io_output ? proc_5_io_next_header_48 : _GEN_2869; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2934 = 3'h5 == encoders_4_io_output ? proc_5_io_next_header_49 : _GEN_2870; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2935 = 3'h5 == encoders_4_io_output ? proc_5_io_next_header_50 : _GEN_2871; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2936 = 3'h5 == encoders_4_io_output ? proc_5_io_next_header_51 : _GEN_2872; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2937 = 3'h5 == encoders_4_io_output ? proc_5_io_next_header_52 : _GEN_2873; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2938 = 3'h5 == encoders_4_io_output ? proc_5_io_next_header_53 : _GEN_2874; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2939 = 3'h5 == encoders_4_io_output ? proc_5_io_next_header_54 : _GEN_2875; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2940 = 3'h5 == encoders_4_io_output ? proc_5_io_next_header_55 : _GEN_2876; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2941 = 3'h5 == encoders_4_io_output ? proc_5_io_next_header_56 : _GEN_2877; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2942 = 3'h5 == encoders_4_io_output ? proc_5_io_next_header_57 : _GEN_2878; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2943 = 3'h5 == encoders_4_io_output ? proc_5_io_next_header_58 : _GEN_2879; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2944 = 3'h5 == encoders_4_io_output ? proc_5_io_next_header_59 : _GEN_2880; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2945 = 3'h5 == encoders_4_io_output ? proc_5_io_next_header_60 : _GEN_2881; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2946 = 3'h5 == encoders_4_io_output ? proc_5_io_next_header_61 : _GEN_2882; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2947 = 3'h5 == encoders_4_io_output ? proc_5_io_next_header_62 : _GEN_2883; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2948 = 3'h5 == encoders_4_io_output ? proc_5_io_next_header_63 : _GEN_2884; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2949 = 3'h6 == encoders_4_io_output ? proc_6_io_next_header_0 : _GEN_2885; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2950 = 3'h6 == encoders_4_io_output ? proc_6_io_next_header_1 : _GEN_2886; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2951 = 3'h6 == encoders_4_io_output ? proc_6_io_next_header_2 : _GEN_2887; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2952 = 3'h6 == encoders_4_io_output ? proc_6_io_next_header_3 : _GEN_2888; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2953 = 3'h6 == encoders_4_io_output ? proc_6_io_next_header_4 : _GEN_2889; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2954 = 3'h6 == encoders_4_io_output ? proc_6_io_next_header_5 : _GEN_2890; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2955 = 3'h6 == encoders_4_io_output ? proc_6_io_next_header_6 : _GEN_2891; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2956 = 3'h6 == encoders_4_io_output ? proc_6_io_next_header_7 : _GEN_2892; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2957 = 3'h6 == encoders_4_io_output ? proc_6_io_next_header_8 : _GEN_2893; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2958 = 3'h6 == encoders_4_io_output ? proc_6_io_next_header_9 : _GEN_2894; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2959 = 3'h6 == encoders_4_io_output ? proc_6_io_next_header_10 : _GEN_2895; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2960 = 3'h6 == encoders_4_io_output ? proc_6_io_next_header_11 : _GEN_2896; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2961 = 3'h6 == encoders_4_io_output ? proc_6_io_next_header_12 : _GEN_2897; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2962 = 3'h6 == encoders_4_io_output ? proc_6_io_next_header_13 : _GEN_2898; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2963 = 3'h6 == encoders_4_io_output ? proc_6_io_next_header_14 : _GEN_2899; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2964 = 3'h6 == encoders_4_io_output ? proc_6_io_next_header_15 : _GEN_2900; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2965 = 3'h6 == encoders_4_io_output ? proc_6_io_next_header_16 : _GEN_2901; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2966 = 3'h6 == encoders_4_io_output ? proc_6_io_next_header_17 : _GEN_2902; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2967 = 3'h6 == encoders_4_io_output ? proc_6_io_next_header_18 : _GEN_2903; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2968 = 3'h6 == encoders_4_io_output ? proc_6_io_next_header_19 : _GEN_2904; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2969 = 3'h6 == encoders_4_io_output ? proc_6_io_next_header_20 : _GEN_2905; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2970 = 3'h6 == encoders_4_io_output ? proc_6_io_next_header_21 : _GEN_2906; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2971 = 3'h6 == encoders_4_io_output ? proc_6_io_next_header_22 : _GEN_2907; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2972 = 3'h6 == encoders_4_io_output ? proc_6_io_next_header_23 : _GEN_2908; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2973 = 3'h6 == encoders_4_io_output ? proc_6_io_next_header_24 : _GEN_2909; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2974 = 3'h6 == encoders_4_io_output ? proc_6_io_next_header_25 : _GEN_2910; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2975 = 3'h6 == encoders_4_io_output ? proc_6_io_next_header_26 : _GEN_2911; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2976 = 3'h6 == encoders_4_io_output ? proc_6_io_next_header_27 : _GEN_2912; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2977 = 3'h6 == encoders_4_io_output ? proc_6_io_next_header_28 : _GEN_2913; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2978 = 3'h6 == encoders_4_io_output ? proc_6_io_next_header_29 : _GEN_2914; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2979 = 3'h6 == encoders_4_io_output ? proc_6_io_next_header_30 : _GEN_2915; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2980 = 3'h6 == encoders_4_io_output ? proc_6_io_next_header_31 : _GEN_2916; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2981 = 3'h6 == encoders_4_io_output ? proc_6_io_next_header_32 : _GEN_2917; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2982 = 3'h6 == encoders_4_io_output ? proc_6_io_next_header_33 : _GEN_2918; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2983 = 3'h6 == encoders_4_io_output ? proc_6_io_next_header_34 : _GEN_2919; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2984 = 3'h6 == encoders_4_io_output ? proc_6_io_next_header_35 : _GEN_2920; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2985 = 3'h6 == encoders_4_io_output ? proc_6_io_next_header_36 : _GEN_2921; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2986 = 3'h6 == encoders_4_io_output ? proc_6_io_next_header_37 : _GEN_2922; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2987 = 3'h6 == encoders_4_io_output ? proc_6_io_next_header_38 : _GEN_2923; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2988 = 3'h6 == encoders_4_io_output ? proc_6_io_next_header_39 : _GEN_2924; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2989 = 3'h6 == encoders_4_io_output ? proc_6_io_next_header_40 : _GEN_2925; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2990 = 3'h6 == encoders_4_io_output ? proc_6_io_next_header_41 : _GEN_2926; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2991 = 3'h6 == encoders_4_io_output ? proc_6_io_next_header_42 : _GEN_2927; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2992 = 3'h6 == encoders_4_io_output ? proc_6_io_next_header_43 : _GEN_2928; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2993 = 3'h6 == encoders_4_io_output ? proc_6_io_next_header_44 : _GEN_2929; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2994 = 3'h6 == encoders_4_io_output ? proc_6_io_next_header_45 : _GEN_2930; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2995 = 3'h6 == encoders_4_io_output ? proc_6_io_next_header_46 : _GEN_2931; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2996 = 3'h6 == encoders_4_io_output ? proc_6_io_next_header_47 : _GEN_2932; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2997 = 3'h6 == encoders_4_io_output ? proc_6_io_next_header_48 : _GEN_2933; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2998 = 3'h6 == encoders_4_io_output ? proc_6_io_next_header_49 : _GEN_2934; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_2999 = 3'h6 == encoders_4_io_output ? proc_6_io_next_header_50 : _GEN_2935; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3000 = 3'h6 == encoders_4_io_output ? proc_6_io_next_header_51 : _GEN_2936; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3001 = 3'h6 == encoders_4_io_output ? proc_6_io_next_header_52 : _GEN_2937; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3002 = 3'h6 == encoders_4_io_output ? proc_6_io_next_header_53 : _GEN_2938; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3003 = 3'h6 == encoders_4_io_output ? proc_6_io_next_header_54 : _GEN_2939; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3004 = 3'h6 == encoders_4_io_output ? proc_6_io_next_header_55 : _GEN_2940; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3005 = 3'h6 == encoders_4_io_output ? proc_6_io_next_header_56 : _GEN_2941; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3006 = 3'h6 == encoders_4_io_output ? proc_6_io_next_header_57 : _GEN_2942; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3007 = 3'h6 == encoders_4_io_output ? proc_6_io_next_header_58 : _GEN_2943; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3008 = 3'h6 == encoders_4_io_output ? proc_6_io_next_header_59 : _GEN_2944; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3009 = 3'h6 == encoders_4_io_output ? proc_6_io_next_header_60 : _GEN_2945; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3010 = 3'h6 == encoders_4_io_output ? proc_6_io_next_header_61 : _GEN_2946; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3011 = 3'h6 == encoders_4_io_output ? proc_6_io_next_header_62 : _GEN_2947; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3012 = 3'h6 == encoders_4_io_output ? proc_6_io_next_header_63 : _GEN_2948; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3013 = 3'h7 == encoders_4_io_output ? proc_7_io_next_header_0 : _GEN_2949; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3014 = 3'h7 == encoders_4_io_output ? proc_7_io_next_header_1 : _GEN_2950; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3015 = 3'h7 == encoders_4_io_output ? proc_7_io_next_header_2 : _GEN_2951; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3016 = 3'h7 == encoders_4_io_output ? proc_7_io_next_header_3 : _GEN_2952; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3017 = 3'h7 == encoders_4_io_output ? proc_7_io_next_header_4 : _GEN_2953; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3018 = 3'h7 == encoders_4_io_output ? proc_7_io_next_header_5 : _GEN_2954; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3019 = 3'h7 == encoders_4_io_output ? proc_7_io_next_header_6 : _GEN_2955; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3020 = 3'h7 == encoders_4_io_output ? proc_7_io_next_header_7 : _GEN_2956; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3021 = 3'h7 == encoders_4_io_output ? proc_7_io_next_header_8 : _GEN_2957; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3022 = 3'h7 == encoders_4_io_output ? proc_7_io_next_header_9 : _GEN_2958; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3023 = 3'h7 == encoders_4_io_output ? proc_7_io_next_header_10 : _GEN_2959; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3024 = 3'h7 == encoders_4_io_output ? proc_7_io_next_header_11 : _GEN_2960; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3025 = 3'h7 == encoders_4_io_output ? proc_7_io_next_header_12 : _GEN_2961; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3026 = 3'h7 == encoders_4_io_output ? proc_7_io_next_header_13 : _GEN_2962; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3027 = 3'h7 == encoders_4_io_output ? proc_7_io_next_header_14 : _GEN_2963; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3028 = 3'h7 == encoders_4_io_output ? proc_7_io_next_header_15 : _GEN_2964; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3029 = 3'h7 == encoders_4_io_output ? proc_7_io_next_header_16 : _GEN_2965; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3030 = 3'h7 == encoders_4_io_output ? proc_7_io_next_header_17 : _GEN_2966; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3031 = 3'h7 == encoders_4_io_output ? proc_7_io_next_header_18 : _GEN_2967; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3032 = 3'h7 == encoders_4_io_output ? proc_7_io_next_header_19 : _GEN_2968; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3033 = 3'h7 == encoders_4_io_output ? proc_7_io_next_header_20 : _GEN_2969; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3034 = 3'h7 == encoders_4_io_output ? proc_7_io_next_header_21 : _GEN_2970; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3035 = 3'h7 == encoders_4_io_output ? proc_7_io_next_header_22 : _GEN_2971; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3036 = 3'h7 == encoders_4_io_output ? proc_7_io_next_header_23 : _GEN_2972; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3037 = 3'h7 == encoders_4_io_output ? proc_7_io_next_header_24 : _GEN_2973; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3038 = 3'h7 == encoders_4_io_output ? proc_7_io_next_header_25 : _GEN_2974; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3039 = 3'h7 == encoders_4_io_output ? proc_7_io_next_header_26 : _GEN_2975; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3040 = 3'h7 == encoders_4_io_output ? proc_7_io_next_header_27 : _GEN_2976; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3041 = 3'h7 == encoders_4_io_output ? proc_7_io_next_header_28 : _GEN_2977; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3042 = 3'h7 == encoders_4_io_output ? proc_7_io_next_header_29 : _GEN_2978; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3043 = 3'h7 == encoders_4_io_output ? proc_7_io_next_header_30 : _GEN_2979; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3044 = 3'h7 == encoders_4_io_output ? proc_7_io_next_header_31 : _GEN_2980; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3045 = 3'h7 == encoders_4_io_output ? proc_7_io_next_header_32 : _GEN_2981; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3046 = 3'h7 == encoders_4_io_output ? proc_7_io_next_header_33 : _GEN_2982; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3047 = 3'h7 == encoders_4_io_output ? proc_7_io_next_header_34 : _GEN_2983; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3048 = 3'h7 == encoders_4_io_output ? proc_7_io_next_header_35 : _GEN_2984; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3049 = 3'h7 == encoders_4_io_output ? proc_7_io_next_header_36 : _GEN_2985; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3050 = 3'h7 == encoders_4_io_output ? proc_7_io_next_header_37 : _GEN_2986; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3051 = 3'h7 == encoders_4_io_output ? proc_7_io_next_header_38 : _GEN_2987; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3052 = 3'h7 == encoders_4_io_output ? proc_7_io_next_header_39 : _GEN_2988; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3053 = 3'h7 == encoders_4_io_output ? proc_7_io_next_header_40 : _GEN_2989; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3054 = 3'h7 == encoders_4_io_output ? proc_7_io_next_header_41 : _GEN_2990; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3055 = 3'h7 == encoders_4_io_output ? proc_7_io_next_header_42 : _GEN_2991; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3056 = 3'h7 == encoders_4_io_output ? proc_7_io_next_header_43 : _GEN_2992; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3057 = 3'h7 == encoders_4_io_output ? proc_7_io_next_header_44 : _GEN_2993; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3058 = 3'h7 == encoders_4_io_output ? proc_7_io_next_header_45 : _GEN_2994; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3059 = 3'h7 == encoders_4_io_output ? proc_7_io_next_header_46 : _GEN_2995; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3060 = 3'h7 == encoders_4_io_output ? proc_7_io_next_header_47 : _GEN_2996; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3061 = 3'h7 == encoders_4_io_output ? proc_7_io_next_header_48 : _GEN_2997; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3062 = 3'h7 == encoders_4_io_output ? proc_7_io_next_header_49 : _GEN_2998; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3063 = 3'h7 == encoders_4_io_output ? proc_7_io_next_header_50 : _GEN_2999; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3064 = 3'h7 == encoders_4_io_output ? proc_7_io_next_header_51 : _GEN_3000; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3065 = 3'h7 == encoders_4_io_output ? proc_7_io_next_header_52 : _GEN_3001; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3066 = 3'h7 == encoders_4_io_output ? proc_7_io_next_header_53 : _GEN_3002; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3067 = 3'h7 == encoders_4_io_output ? proc_7_io_next_header_54 : _GEN_3003; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3068 = 3'h7 == encoders_4_io_output ? proc_7_io_next_header_55 : _GEN_3004; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3069 = 3'h7 == encoders_4_io_output ? proc_7_io_next_header_56 : _GEN_3005; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3070 = 3'h7 == encoders_4_io_output ? proc_7_io_next_header_57 : _GEN_3006; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3071 = 3'h7 == encoders_4_io_output ? proc_7_io_next_header_58 : _GEN_3007; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3072 = 3'h7 == encoders_4_io_output ? proc_7_io_next_header_59 : _GEN_3008; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3073 = 3'h7 == encoders_4_io_output ? proc_7_io_next_header_60 : _GEN_3009; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3074 = 3'h7 == encoders_4_io_output ? proc_7_io_next_header_61 : _GEN_3010; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3075 = 3'h7 == encoders_4_io_output ? proc_7_io_next_header_62 : _GEN_3011; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3076 = 3'h7 == encoders_4_io_output ? proc_7_io_next_header_63 : _GEN_3012; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3142 = 3'h0 == encoders_5_io_output ? proc_0_io_next_header_0 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3143 = 3'h0 == encoders_5_io_output ? proc_0_io_next_header_1 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3144 = 3'h0 == encoders_5_io_output ? proc_0_io_next_header_2 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3145 = 3'h0 == encoders_5_io_output ? proc_0_io_next_header_3 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3146 = 3'h0 == encoders_5_io_output ? proc_0_io_next_header_4 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3147 = 3'h0 == encoders_5_io_output ? proc_0_io_next_header_5 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3148 = 3'h0 == encoders_5_io_output ? proc_0_io_next_header_6 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3149 = 3'h0 == encoders_5_io_output ? proc_0_io_next_header_7 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3150 = 3'h0 == encoders_5_io_output ? proc_0_io_next_header_8 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3151 = 3'h0 == encoders_5_io_output ? proc_0_io_next_header_9 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3152 = 3'h0 == encoders_5_io_output ? proc_0_io_next_header_10 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3153 = 3'h0 == encoders_5_io_output ? proc_0_io_next_header_11 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3154 = 3'h0 == encoders_5_io_output ? proc_0_io_next_header_12 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3155 = 3'h0 == encoders_5_io_output ? proc_0_io_next_header_13 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3156 = 3'h0 == encoders_5_io_output ? proc_0_io_next_header_14 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3157 = 3'h0 == encoders_5_io_output ? proc_0_io_next_header_15 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3158 = 3'h0 == encoders_5_io_output ? proc_0_io_next_header_16 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3159 = 3'h0 == encoders_5_io_output ? proc_0_io_next_header_17 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3160 = 3'h0 == encoders_5_io_output ? proc_0_io_next_header_18 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3161 = 3'h0 == encoders_5_io_output ? proc_0_io_next_header_19 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3162 = 3'h0 == encoders_5_io_output ? proc_0_io_next_header_20 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3163 = 3'h0 == encoders_5_io_output ? proc_0_io_next_header_21 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3164 = 3'h0 == encoders_5_io_output ? proc_0_io_next_header_22 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3165 = 3'h0 == encoders_5_io_output ? proc_0_io_next_header_23 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3166 = 3'h0 == encoders_5_io_output ? proc_0_io_next_header_24 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3167 = 3'h0 == encoders_5_io_output ? proc_0_io_next_header_25 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3168 = 3'h0 == encoders_5_io_output ? proc_0_io_next_header_26 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3169 = 3'h0 == encoders_5_io_output ? proc_0_io_next_header_27 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3170 = 3'h0 == encoders_5_io_output ? proc_0_io_next_header_28 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3171 = 3'h0 == encoders_5_io_output ? proc_0_io_next_header_29 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3172 = 3'h0 == encoders_5_io_output ? proc_0_io_next_header_30 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3173 = 3'h0 == encoders_5_io_output ? proc_0_io_next_header_31 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3174 = 3'h0 == encoders_5_io_output ? proc_0_io_next_header_32 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3175 = 3'h0 == encoders_5_io_output ? proc_0_io_next_header_33 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3176 = 3'h0 == encoders_5_io_output ? proc_0_io_next_header_34 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3177 = 3'h0 == encoders_5_io_output ? proc_0_io_next_header_35 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3178 = 3'h0 == encoders_5_io_output ? proc_0_io_next_header_36 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3179 = 3'h0 == encoders_5_io_output ? proc_0_io_next_header_37 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3180 = 3'h0 == encoders_5_io_output ? proc_0_io_next_header_38 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3181 = 3'h0 == encoders_5_io_output ? proc_0_io_next_header_39 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3182 = 3'h0 == encoders_5_io_output ? proc_0_io_next_header_40 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3183 = 3'h0 == encoders_5_io_output ? proc_0_io_next_header_41 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3184 = 3'h0 == encoders_5_io_output ? proc_0_io_next_header_42 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3185 = 3'h0 == encoders_5_io_output ? proc_0_io_next_header_43 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3186 = 3'h0 == encoders_5_io_output ? proc_0_io_next_header_44 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3187 = 3'h0 == encoders_5_io_output ? proc_0_io_next_header_45 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3188 = 3'h0 == encoders_5_io_output ? proc_0_io_next_header_46 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3189 = 3'h0 == encoders_5_io_output ? proc_0_io_next_header_47 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3190 = 3'h0 == encoders_5_io_output ? proc_0_io_next_header_48 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3191 = 3'h0 == encoders_5_io_output ? proc_0_io_next_header_49 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3192 = 3'h0 == encoders_5_io_output ? proc_0_io_next_header_50 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3193 = 3'h0 == encoders_5_io_output ? proc_0_io_next_header_51 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3194 = 3'h0 == encoders_5_io_output ? proc_0_io_next_header_52 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3195 = 3'h0 == encoders_5_io_output ? proc_0_io_next_header_53 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3196 = 3'h0 == encoders_5_io_output ? proc_0_io_next_header_54 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3197 = 3'h0 == encoders_5_io_output ? proc_0_io_next_header_55 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3198 = 3'h0 == encoders_5_io_output ? proc_0_io_next_header_56 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3199 = 3'h0 == encoders_5_io_output ? proc_0_io_next_header_57 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3200 = 3'h0 == encoders_5_io_output ? proc_0_io_next_header_58 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3201 = 3'h0 == encoders_5_io_output ? proc_0_io_next_header_59 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3202 = 3'h0 == encoders_5_io_output ? proc_0_io_next_header_60 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3203 = 3'h0 == encoders_5_io_output ? proc_0_io_next_header_61 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3204 = 3'h0 == encoders_5_io_output ? proc_0_io_next_header_62 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3205 = 3'h0 == encoders_5_io_output ? proc_0_io_next_header_63 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3206 = 3'h1 == encoders_5_io_output ? proc_1_io_next_header_0 : _GEN_3142; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3207 = 3'h1 == encoders_5_io_output ? proc_1_io_next_header_1 : _GEN_3143; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3208 = 3'h1 == encoders_5_io_output ? proc_1_io_next_header_2 : _GEN_3144; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3209 = 3'h1 == encoders_5_io_output ? proc_1_io_next_header_3 : _GEN_3145; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3210 = 3'h1 == encoders_5_io_output ? proc_1_io_next_header_4 : _GEN_3146; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3211 = 3'h1 == encoders_5_io_output ? proc_1_io_next_header_5 : _GEN_3147; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3212 = 3'h1 == encoders_5_io_output ? proc_1_io_next_header_6 : _GEN_3148; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3213 = 3'h1 == encoders_5_io_output ? proc_1_io_next_header_7 : _GEN_3149; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3214 = 3'h1 == encoders_5_io_output ? proc_1_io_next_header_8 : _GEN_3150; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3215 = 3'h1 == encoders_5_io_output ? proc_1_io_next_header_9 : _GEN_3151; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3216 = 3'h1 == encoders_5_io_output ? proc_1_io_next_header_10 : _GEN_3152; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3217 = 3'h1 == encoders_5_io_output ? proc_1_io_next_header_11 : _GEN_3153; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3218 = 3'h1 == encoders_5_io_output ? proc_1_io_next_header_12 : _GEN_3154; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3219 = 3'h1 == encoders_5_io_output ? proc_1_io_next_header_13 : _GEN_3155; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3220 = 3'h1 == encoders_5_io_output ? proc_1_io_next_header_14 : _GEN_3156; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3221 = 3'h1 == encoders_5_io_output ? proc_1_io_next_header_15 : _GEN_3157; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3222 = 3'h1 == encoders_5_io_output ? proc_1_io_next_header_16 : _GEN_3158; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3223 = 3'h1 == encoders_5_io_output ? proc_1_io_next_header_17 : _GEN_3159; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3224 = 3'h1 == encoders_5_io_output ? proc_1_io_next_header_18 : _GEN_3160; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3225 = 3'h1 == encoders_5_io_output ? proc_1_io_next_header_19 : _GEN_3161; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3226 = 3'h1 == encoders_5_io_output ? proc_1_io_next_header_20 : _GEN_3162; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3227 = 3'h1 == encoders_5_io_output ? proc_1_io_next_header_21 : _GEN_3163; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3228 = 3'h1 == encoders_5_io_output ? proc_1_io_next_header_22 : _GEN_3164; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3229 = 3'h1 == encoders_5_io_output ? proc_1_io_next_header_23 : _GEN_3165; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3230 = 3'h1 == encoders_5_io_output ? proc_1_io_next_header_24 : _GEN_3166; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3231 = 3'h1 == encoders_5_io_output ? proc_1_io_next_header_25 : _GEN_3167; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3232 = 3'h1 == encoders_5_io_output ? proc_1_io_next_header_26 : _GEN_3168; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3233 = 3'h1 == encoders_5_io_output ? proc_1_io_next_header_27 : _GEN_3169; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3234 = 3'h1 == encoders_5_io_output ? proc_1_io_next_header_28 : _GEN_3170; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3235 = 3'h1 == encoders_5_io_output ? proc_1_io_next_header_29 : _GEN_3171; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3236 = 3'h1 == encoders_5_io_output ? proc_1_io_next_header_30 : _GEN_3172; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3237 = 3'h1 == encoders_5_io_output ? proc_1_io_next_header_31 : _GEN_3173; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3238 = 3'h1 == encoders_5_io_output ? proc_1_io_next_header_32 : _GEN_3174; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3239 = 3'h1 == encoders_5_io_output ? proc_1_io_next_header_33 : _GEN_3175; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3240 = 3'h1 == encoders_5_io_output ? proc_1_io_next_header_34 : _GEN_3176; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3241 = 3'h1 == encoders_5_io_output ? proc_1_io_next_header_35 : _GEN_3177; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3242 = 3'h1 == encoders_5_io_output ? proc_1_io_next_header_36 : _GEN_3178; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3243 = 3'h1 == encoders_5_io_output ? proc_1_io_next_header_37 : _GEN_3179; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3244 = 3'h1 == encoders_5_io_output ? proc_1_io_next_header_38 : _GEN_3180; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3245 = 3'h1 == encoders_5_io_output ? proc_1_io_next_header_39 : _GEN_3181; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3246 = 3'h1 == encoders_5_io_output ? proc_1_io_next_header_40 : _GEN_3182; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3247 = 3'h1 == encoders_5_io_output ? proc_1_io_next_header_41 : _GEN_3183; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3248 = 3'h1 == encoders_5_io_output ? proc_1_io_next_header_42 : _GEN_3184; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3249 = 3'h1 == encoders_5_io_output ? proc_1_io_next_header_43 : _GEN_3185; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3250 = 3'h1 == encoders_5_io_output ? proc_1_io_next_header_44 : _GEN_3186; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3251 = 3'h1 == encoders_5_io_output ? proc_1_io_next_header_45 : _GEN_3187; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3252 = 3'h1 == encoders_5_io_output ? proc_1_io_next_header_46 : _GEN_3188; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3253 = 3'h1 == encoders_5_io_output ? proc_1_io_next_header_47 : _GEN_3189; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3254 = 3'h1 == encoders_5_io_output ? proc_1_io_next_header_48 : _GEN_3190; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3255 = 3'h1 == encoders_5_io_output ? proc_1_io_next_header_49 : _GEN_3191; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3256 = 3'h1 == encoders_5_io_output ? proc_1_io_next_header_50 : _GEN_3192; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3257 = 3'h1 == encoders_5_io_output ? proc_1_io_next_header_51 : _GEN_3193; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3258 = 3'h1 == encoders_5_io_output ? proc_1_io_next_header_52 : _GEN_3194; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3259 = 3'h1 == encoders_5_io_output ? proc_1_io_next_header_53 : _GEN_3195; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3260 = 3'h1 == encoders_5_io_output ? proc_1_io_next_header_54 : _GEN_3196; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3261 = 3'h1 == encoders_5_io_output ? proc_1_io_next_header_55 : _GEN_3197; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3262 = 3'h1 == encoders_5_io_output ? proc_1_io_next_header_56 : _GEN_3198; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3263 = 3'h1 == encoders_5_io_output ? proc_1_io_next_header_57 : _GEN_3199; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3264 = 3'h1 == encoders_5_io_output ? proc_1_io_next_header_58 : _GEN_3200; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3265 = 3'h1 == encoders_5_io_output ? proc_1_io_next_header_59 : _GEN_3201; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3266 = 3'h1 == encoders_5_io_output ? proc_1_io_next_header_60 : _GEN_3202; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3267 = 3'h1 == encoders_5_io_output ? proc_1_io_next_header_61 : _GEN_3203; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3268 = 3'h1 == encoders_5_io_output ? proc_1_io_next_header_62 : _GEN_3204; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3269 = 3'h1 == encoders_5_io_output ? proc_1_io_next_header_63 : _GEN_3205; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3270 = 3'h2 == encoders_5_io_output ? proc_2_io_next_header_0 : _GEN_3206; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3271 = 3'h2 == encoders_5_io_output ? proc_2_io_next_header_1 : _GEN_3207; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3272 = 3'h2 == encoders_5_io_output ? proc_2_io_next_header_2 : _GEN_3208; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3273 = 3'h2 == encoders_5_io_output ? proc_2_io_next_header_3 : _GEN_3209; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3274 = 3'h2 == encoders_5_io_output ? proc_2_io_next_header_4 : _GEN_3210; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3275 = 3'h2 == encoders_5_io_output ? proc_2_io_next_header_5 : _GEN_3211; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3276 = 3'h2 == encoders_5_io_output ? proc_2_io_next_header_6 : _GEN_3212; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3277 = 3'h2 == encoders_5_io_output ? proc_2_io_next_header_7 : _GEN_3213; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3278 = 3'h2 == encoders_5_io_output ? proc_2_io_next_header_8 : _GEN_3214; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3279 = 3'h2 == encoders_5_io_output ? proc_2_io_next_header_9 : _GEN_3215; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3280 = 3'h2 == encoders_5_io_output ? proc_2_io_next_header_10 : _GEN_3216; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3281 = 3'h2 == encoders_5_io_output ? proc_2_io_next_header_11 : _GEN_3217; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3282 = 3'h2 == encoders_5_io_output ? proc_2_io_next_header_12 : _GEN_3218; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3283 = 3'h2 == encoders_5_io_output ? proc_2_io_next_header_13 : _GEN_3219; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3284 = 3'h2 == encoders_5_io_output ? proc_2_io_next_header_14 : _GEN_3220; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3285 = 3'h2 == encoders_5_io_output ? proc_2_io_next_header_15 : _GEN_3221; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3286 = 3'h2 == encoders_5_io_output ? proc_2_io_next_header_16 : _GEN_3222; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3287 = 3'h2 == encoders_5_io_output ? proc_2_io_next_header_17 : _GEN_3223; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3288 = 3'h2 == encoders_5_io_output ? proc_2_io_next_header_18 : _GEN_3224; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3289 = 3'h2 == encoders_5_io_output ? proc_2_io_next_header_19 : _GEN_3225; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3290 = 3'h2 == encoders_5_io_output ? proc_2_io_next_header_20 : _GEN_3226; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3291 = 3'h2 == encoders_5_io_output ? proc_2_io_next_header_21 : _GEN_3227; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3292 = 3'h2 == encoders_5_io_output ? proc_2_io_next_header_22 : _GEN_3228; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3293 = 3'h2 == encoders_5_io_output ? proc_2_io_next_header_23 : _GEN_3229; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3294 = 3'h2 == encoders_5_io_output ? proc_2_io_next_header_24 : _GEN_3230; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3295 = 3'h2 == encoders_5_io_output ? proc_2_io_next_header_25 : _GEN_3231; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3296 = 3'h2 == encoders_5_io_output ? proc_2_io_next_header_26 : _GEN_3232; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3297 = 3'h2 == encoders_5_io_output ? proc_2_io_next_header_27 : _GEN_3233; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3298 = 3'h2 == encoders_5_io_output ? proc_2_io_next_header_28 : _GEN_3234; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3299 = 3'h2 == encoders_5_io_output ? proc_2_io_next_header_29 : _GEN_3235; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3300 = 3'h2 == encoders_5_io_output ? proc_2_io_next_header_30 : _GEN_3236; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3301 = 3'h2 == encoders_5_io_output ? proc_2_io_next_header_31 : _GEN_3237; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3302 = 3'h2 == encoders_5_io_output ? proc_2_io_next_header_32 : _GEN_3238; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3303 = 3'h2 == encoders_5_io_output ? proc_2_io_next_header_33 : _GEN_3239; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3304 = 3'h2 == encoders_5_io_output ? proc_2_io_next_header_34 : _GEN_3240; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3305 = 3'h2 == encoders_5_io_output ? proc_2_io_next_header_35 : _GEN_3241; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3306 = 3'h2 == encoders_5_io_output ? proc_2_io_next_header_36 : _GEN_3242; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3307 = 3'h2 == encoders_5_io_output ? proc_2_io_next_header_37 : _GEN_3243; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3308 = 3'h2 == encoders_5_io_output ? proc_2_io_next_header_38 : _GEN_3244; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3309 = 3'h2 == encoders_5_io_output ? proc_2_io_next_header_39 : _GEN_3245; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3310 = 3'h2 == encoders_5_io_output ? proc_2_io_next_header_40 : _GEN_3246; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3311 = 3'h2 == encoders_5_io_output ? proc_2_io_next_header_41 : _GEN_3247; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3312 = 3'h2 == encoders_5_io_output ? proc_2_io_next_header_42 : _GEN_3248; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3313 = 3'h2 == encoders_5_io_output ? proc_2_io_next_header_43 : _GEN_3249; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3314 = 3'h2 == encoders_5_io_output ? proc_2_io_next_header_44 : _GEN_3250; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3315 = 3'h2 == encoders_5_io_output ? proc_2_io_next_header_45 : _GEN_3251; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3316 = 3'h2 == encoders_5_io_output ? proc_2_io_next_header_46 : _GEN_3252; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3317 = 3'h2 == encoders_5_io_output ? proc_2_io_next_header_47 : _GEN_3253; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3318 = 3'h2 == encoders_5_io_output ? proc_2_io_next_header_48 : _GEN_3254; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3319 = 3'h2 == encoders_5_io_output ? proc_2_io_next_header_49 : _GEN_3255; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3320 = 3'h2 == encoders_5_io_output ? proc_2_io_next_header_50 : _GEN_3256; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3321 = 3'h2 == encoders_5_io_output ? proc_2_io_next_header_51 : _GEN_3257; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3322 = 3'h2 == encoders_5_io_output ? proc_2_io_next_header_52 : _GEN_3258; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3323 = 3'h2 == encoders_5_io_output ? proc_2_io_next_header_53 : _GEN_3259; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3324 = 3'h2 == encoders_5_io_output ? proc_2_io_next_header_54 : _GEN_3260; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3325 = 3'h2 == encoders_5_io_output ? proc_2_io_next_header_55 : _GEN_3261; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3326 = 3'h2 == encoders_5_io_output ? proc_2_io_next_header_56 : _GEN_3262; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3327 = 3'h2 == encoders_5_io_output ? proc_2_io_next_header_57 : _GEN_3263; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3328 = 3'h2 == encoders_5_io_output ? proc_2_io_next_header_58 : _GEN_3264; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3329 = 3'h2 == encoders_5_io_output ? proc_2_io_next_header_59 : _GEN_3265; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3330 = 3'h2 == encoders_5_io_output ? proc_2_io_next_header_60 : _GEN_3266; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3331 = 3'h2 == encoders_5_io_output ? proc_2_io_next_header_61 : _GEN_3267; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3332 = 3'h2 == encoders_5_io_output ? proc_2_io_next_header_62 : _GEN_3268; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3333 = 3'h2 == encoders_5_io_output ? proc_2_io_next_header_63 : _GEN_3269; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3334 = 3'h3 == encoders_5_io_output ? proc_3_io_next_header_0 : _GEN_3270; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3335 = 3'h3 == encoders_5_io_output ? proc_3_io_next_header_1 : _GEN_3271; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3336 = 3'h3 == encoders_5_io_output ? proc_3_io_next_header_2 : _GEN_3272; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3337 = 3'h3 == encoders_5_io_output ? proc_3_io_next_header_3 : _GEN_3273; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3338 = 3'h3 == encoders_5_io_output ? proc_3_io_next_header_4 : _GEN_3274; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3339 = 3'h3 == encoders_5_io_output ? proc_3_io_next_header_5 : _GEN_3275; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3340 = 3'h3 == encoders_5_io_output ? proc_3_io_next_header_6 : _GEN_3276; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3341 = 3'h3 == encoders_5_io_output ? proc_3_io_next_header_7 : _GEN_3277; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3342 = 3'h3 == encoders_5_io_output ? proc_3_io_next_header_8 : _GEN_3278; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3343 = 3'h3 == encoders_5_io_output ? proc_3_io_next_header_9 : _GEN_3279; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3344 = 3'h3 == encoders_5_io_output ? proc_3_io_next_header_10 : _GEN_3280; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3345 = 3'h3 == encoders_5_io_output ? proc_3_io_next_header_11 : _GEN_3281; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3346 = 3'h3 == encoders_5_io_output ? proc_3_io_next_header_12 : _GEN_3282; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3347 = 3'h3 == encoders_5_io_output ? proc_3_io_next_header_13 : _GEN_3283; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3348 = 3'h3 == encoders_5_io_output ? proc_3_io_next_header_14 : _GEN_3284; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3349 = 3'h3 == encoders_5_io_output ? proc_3_io_next_header_15 : _GEN_3285; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3350 = 3'h3 == encoders_5_io_output ? proc_3_io_next_header_16 : _GEN_3286; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3351 = 3'h3 == encoders_5_io_output ? proc_3_io_next_header_17 : _GEN_3287; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3352 = 3'h3 == encoders_5_io_output ? proc_3_io_next_header_18 : _GEN_3288; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3353 = 3'h3 == encoders_5_io_output ? proc_3_io_next_header_19 : _GEN_3289; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3354 = 3'h3 == encoders_5_io_output ? proc_3_io_next_header_20 : _GEN_3290; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3355 = 3'h3 == encoders_5_io_output ? proc_3_io_next_header_21 : _GEN_3291; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3356 = 3'h3 == encoders_5_io_output ? proc_3_io_next_header_22 : _GEN_3292; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3357 = 3'h3 == encoders_5_io_output ? proc_3_io_next_header_23 : _GEN_3293; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3358 = 3'h3 == encoders_5_io_output ? proc_3_io_next_header_24 : _GEN_3294; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3359 = 3'h3 == encoders_5_io_output ? proc_3_io_next_header_25 : _GEN_3295; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3360 = 3'h3 == encoders_5_io_output ? proc_3_io_next_header_26 : _GEN_3296; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3361 = 3'h3 == encoders_5_io_output ? proc_3_io_next_header_27 : _GEN_3297; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3362 = 3'h3 == encoders_5_io_output ? proc_3_io_next_header_28 : _GEN_3298; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3363 = 3'h3 == encoders_5_io_output ? proc_3_io_next_header_29 : _GEN_3299; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3364 = 3'h3 == encoders_5_io_output ? proc_3_io_next_header_30 : _GEN_3300; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3365 = 3'h3 == encoders_5_io_output ? proc_3_io_next_header_31 : _GEN_3301; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3366 = 3'h3 == encoders_5_io_output ? proc_3_io_next_header_32 : _GEN_3302; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3367 = 3'h3 == encoders_5_io_output ? proc_3_io_next_header_33 : _GEN_3303; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3368 = 3'h3 == encoders_5_io_output ? proc_3_io_next_header_34 : _GEN_3304; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3369 = 3'h3 == encoders_5_io_output ? proc_3_io_next_header_35 : _GEN_3305; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3370 = 3'h3 == encoders_5_io_output ? proc_3_io_next_header_36 : _GEN_3306; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3371 = 3'h3 == encoders_5_io_output ? proc_3_io_next_header_37 : _GEN_3307; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3372 = 3'h3 == encoders_5_io_output ? proc_3_io_next_header_38 : _GEN_3308; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3373 = 3'h3 == encoders_5_io_output ? proc_3_io_next_header_39 : _GEN_3309; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3374 = 3'h3 == encoders_5_io_output ? proc_3_io_next_header_40 : _GEN_3310; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3375 = 3'h3 == encoders_5_io_output ? proc_3_io_next_header_41 : _GEN_3311; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3376 = 3'h3 == encoders_5_io_output ? proc_3_io_next_header_42 : _GEN_3312; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3377 = 3'h3 == encoders_5_io_output ? proc_3_io_next_header_43 : _GEN_3313; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3378 = 3'h3 == encoders_5_io_output ? proc_3_io_next_header_44 : _GEN_3314; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3379 = 3'h3 == encoders_5_io_output ? proc_3_io_next_header_45 : _GEN_3315; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3380 = 3'h3 == encoders_5_io_output ? proc_3_io_next_header_46 : _GEN_3316; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3381 = 3'h3 == encoders_5_io_output ? proc_3_io_next_header_47 : _GEN_3317; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3382 = 3'h3 == encoders_5_io_output ? proc_3_io_next_header_48 : _GEN_3318; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3383 = 3'h3 == encoders_5_io_output ? proc_3_io_next_header_49 : _GEN_3319; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3384 = 3'h3 == encoders_5_io_output ? proc_3_io_next_header_50 : _GEN_3320; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3385 = 3'h3 == encoders_5_io_output ? proc_3_io_next_header_51 : _GEN_3321; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3386 = 3'h3 == encoders_5_io_output ? proc_3_io_next_header_52 : _GEN_3322; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3387 = 3'h3 == encoders_5_io_output ? proc_3_io_next_header_53 : _GEN_3323; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3388 = 3'h3 == encoders_5_io_output ? proc_3_io_next_header_54 : _GEN_3324; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3389 = 3'h3 == encoders_5_io_output ? proc_3_io_next_header_55 : _GEN_3325; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3390 = 3'h3 == encoders_5_io_output ? proc_3_io_next_header_56 : _GEN_3326; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3391 = 3'h3 == encoders_5_io_output ? proc_3_io_next_header_57 : _GEN_3327; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3392 = 3'h3 == encoders_5_io_output ? proc_3_io_next_header_58 : _GEN_3328; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3393 = 3'h3 == encoders_5_io_output ? proc_3_io_next_header_59 : _GEN_3329; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3394 = 3'h3 == encoders_5_io_output ? proc_3_io_next_header_60 : _GEN_3330; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3395 = 3'h3 == encoders_5_io_output ? proc_3_io_next_header_61 : _GEN_3331; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3396 = 3'h3 == encoders_5_io_output ? proc_3_io_next_header_62 : _GEN_3332; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3397 = 3'h3 == encoders_5_io_output ? proc_3_io_next_header_63 : _GEN_3333; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3398 = 3'h4 == encoders_5_io_output ? proc_4_io_next_header_0 : _GEN_3334; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3399 = 3'h4 == encoders_5_io_output ? proc_4_io_next_header_1 : _GEN_3335; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3400 = 3'h4 == encoders_5_io_output ? proc_4_io_next_header_2 : _GEN_3336; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3401 = 3'h4 == encoders_5_io_output ? proc_4_io_next_header_3 : _GEN_3337; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3402 = 3'h4 == encoders_5_io_output ? proc_4_io_next_header_4 : _GEN_3338; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3403 = 3'h4 == encoders_5_io_output ? proc_4_io_next_header_5 : _GEN_3339; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3404 = 3'h4 == encoders_5_io_output ? proc_4_io_next_header_6 : _GEN_3340; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3405 = 3'h4 == encoders_5_io_output ? proc_4_io_next_header_7 : _GEN_3341; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3406 = 3'h4 == encoders_5_io_output ? proc_4_io_next_header_8 : _GEN_3342; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3407 = 3'h4 == encoders_5_io_output ? proc_4_io_next_header_9 : _GEN_3343; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3408 = 3'h4 == encoders_5_io_output ? proc_4_io_next_header_10 : _GEN_3344; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3409 = 3'h4 == encoders_5_io_output ? proc_4_io_next_header_11 : _GEN_3345; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3410 = 3'h4 == encoders_5_io_output ? proc_4_io_next_header_12 : _GEN_3346; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3411 = 3'h4 == encoders_5_io_output ? proc_4_io_next_header_13 : _GEN_3347; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3412 = 3'h4 == encoders_5_io_output ? proc_4_io_next_header_14 : _GEN_3348; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3413 = 3'h4 == encoders_5_io_output ? proc_4_io_next_header_15 : _GEN_3349; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3414 = 3'h4 == encoders_5_io_output ? proc_4_io_next_header_16 : _GEN_3350; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3415 = 3'h4 == encoders_5_io_output ? proc_4_io_next_header_17 : _GEN_3351; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3416 = 3'h4 == encoders_5_io_output ? proc_4_io_next_header_18 : _GEN_3352; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3417 = 3'h4 == encoders_5_io_output ? proc_4_io_next_header_19 : _GEN_3353; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3418 = 3'h4 == encoders_5_io_output ? proc_4_io_next_header_20 : _GEN_3354; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3419 = 3'h4 == encoders_5_io_output ? proc_4_io_next_header_21 : _GEN_3355; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3420 = 3'h4 == encoders_5_io_output ? proc_4_io_next_header_22 : _GEN_3356; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3421 = 3'h4 == encoders_5_io_output ? proc_4_io_next_header_23 : _GEN_3357; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3422 = 3'h4 == encoders_5_io_output ? proc_4_io_next_header_24 : _GEN_3358; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3423 = 3'h4 == encoders_5_io_output ? proc_4_io_next_header_25 : _GEN_3359; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3424 = 3'h4 == encoders_5_io_output ? proc_4_io_next_header_26 : _GEN_3360; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3425 = 3'h4 == encoders_5_io_output ? proc_4_io_next_header_27 : _GEN_3361; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3426 = 3'h4 == encoders_5_io_output ? proc_4_io_next_header_28 : _GEN_3362; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3427 = 3'h4 == encoders_5_io_output ? proc_4_io_next_header_29 : _GEN_3363; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3428 = 3'h4 == encoders_5_io_output ? proc_4_io_next_header_30 : _GEN_3364; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3429 = 3'h4 == encoders_5_io_output ? proc_4_io_next_header_31 : _GEN_3365; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3430 = 3'h4 == encoders_5_io_output ? proc_4_io_next_header_32 : _GEN_3366; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3431 = 3'h4 == encoders_5_io_output ? proc_4_io_next_header_33 : _GEN_3367; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3432 = 3'h4 == encoders_5_io_output ? proc_4_io_next_header_34 : _GEN_3368; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3433 = 3'h4 == encoders_5_io_output ? proc_4_io_next_header_35 : _GEN_3369; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3434 = 3'h4 == encoders_5_io_output ? proc_4_io_next_header_36 : _GEN_3370; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3435 = 3'h4 == encoders_5_io_output ? proc_4_io_next_header_37 : _GEN_3371; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3436 = 3'h4 == encoders_5_io_output ? proc_4_io_next_header_38 : _GEN_3372; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3437 = 3'h4 == encoders_5_io_output ? proc_4_io_next_header_39 : _GEN_3373; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3438 = 3'h4 == encoders_5_io_output ? proc_4_io_next_header_40 : _GEN_3374; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3439 = 3'h4 == encoders_5_io_output ? proc_4_io_next_header_41 : _GEN_3375; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3440 = 3'h4 == encoders_5_io_output ? proc_4_io_next_header_42 : _GEN_3376; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3441 = 3'h4 == encoders_5_io_output ? proc_4_io_next_header_43 : _GEN_3377; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3442 = 3'h4 == encoders_5_io_output ? proc_4_io_next_header_44 : _GEN_3378; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3443 = 3'h4 == encoders_5_io_output ? proc_4_io_next_header_45 : _GEN_3379; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3444 = 3'h4 == encoders_5_io_output ? proc_4_io_next_header_46 : _GEN_3380; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3445 = 3'h4 == encoders_5_io_output ? proc_4_io_next_header_47 : _GEN_3381; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3446 = 3'h4 == encoders_5_io_output ? proc_4_io_next_header_48 : _GEN_3382; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3447 = 3'h4 == encoders_5_io_output ? proc_4_io_next_header_49 : _GEN_3383; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3448 = 3'h4 == encoders_5_io_output ? proc_4_io_next_header_50 : _GEN_3384; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3449 = 3'h4 == encoders_5_io_output ? proc_4_io_next_header_51 : _GEN_3385; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3450 = 3'h4 == encoders_5_io_output ? proc_4_io_next_header_52 : _GEN_3386; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3451 = 3'h4 == encoders_5_io_output ? proc_4_io_next_header_53 : _GEN_3387; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3452 = 3'h4 == encoders_5_io_output ? proc_4_io_next_header_54 : _GEN_3388; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3453 = 3'h4 == encoders_5_io_output ? proc_4_io_next_header_55 : _GEN_3389; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3454 = 3'h4 == encoders_5_io_output ? proc_4_io_next_header_56 : _GEN_3390; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3455 = 3'h4 == encoders_5_io_output ? proc_4_io_next_header_57 : _GEN_3391; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3456 = 3'h4 == encoders_5_io_output ? proc_4_io_next_header_58 : _GEN_3392; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3457 = 3'h4 == encoders_5_io_output ? proc_4_io_next_header_59 : _GEN_3393; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3458 = 3'h4 == encoders_5_io_output ? proc_4_io_next_header_60 : _GEN_3394; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3459 = 3'h4 == encoders_5_io_output ? proc_4_io_next_header_61 : _GEN_3395; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3460 = 3'h4 == encoders_5_io_output ? proc_4_io_next_header_62 : _GEN_3396; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3461 = 3'h4 == encoders_5_io_output ? proc_4_io_next_header_63 : _GEN_3397; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3462 = 3'h5 == encoders_5_io_output ? proc_5_io_next_header_0 : _GEN_3398; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3463 = 3'h5 == encoders_5_io_output ? proc_5_io_next_header_1 : _GEN_3399; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3464 = 3'h5 == encoders_5_io_output ? proc_5_io_next_header_2 : _GEN_3400; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3465 = 3'h5 == encoders_5_io_output ? proc_5_io_next_header_3 : _GEN_3401; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3466 = 3'h5 == encoders_5_io_output ? proc_5_io_next_header_4 : _GEN_3402; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3467 = 3'h5 == encoders_5_io_output ? proc_5_io_next_header_5 : _GEN_3403; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3468 = 3'h5 == encoders_5_io_output ? proc_5_io_next_header_6 : _GEN_3404; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3469 = 3'h5 == encoders_5_io_output ? proc_5_io_next_header_7 : _GEN_3405; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3470 = 3'h5 == encoders_5_io_output ? proc_5_io_next_header_8 : _GEN_3406; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3471 = 3'h5 == encoders_5_io_output ? proc_5_io_next_header_9 : _GEN_3407; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3472 = 3'h5 == encoders_5_io_output ? proc_5_io_next_header_10 : _GEN_3408; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3473 = 3'h5 == encoders_5_io_output ? proc_5_io_next_header_11 : _GEN_3409; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3474 = 3'h5 == encoders_5_io_output ? proc_5_io_next_header_12 : _GEN_3410; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3475 = 3'h5 == encoders_5_io_output ? proc_5_io_next_header_13 : _GEN_3411; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3476 = 3'h5 == encoders_5_io_output ? proc_5_io_next_header_14 : _GEN_3412; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3477 = 3'h5 == encoders_5_io_output ? proc_5_io_next_header_15 : _GEN_3413; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3478 = 3'h5 == encoders_5_io_output ? proc_5_io_next_header_16 : _GEN_3414; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3479 = 3'h5 == encoders_5_io_output ? proc_5_io_next_header_17 : _GEN_3415; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3480 = 3'h5 == encoders_5_io_output ? proc_5_io_next_header_18 : _GEN_3416; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3481 = 3'h5 == encoders_5_io_output ? proc_5_io_next_header_19 : _GEN_3417; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3482 = 3'h5 == encoders_5_io_output ? proc_5_io_next_header_20 : _GEN_3418; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3483 = 3'h5 == encoders_5_io_output ? proc_5_io_next_header_21 : _GEN_3419; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3484 = 3'h5 == encoders_5_io_output ? proc_5_io_next_header_22 : _GEN_3420; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3485 = 3'h5 == encoders_5_io_output ? proc_5_io_next_header_23 : _GEN_3421; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3486 = 3'h5 == encoders_5_io_output ? proc_5_io_next_header_24 : _GEN_3422; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3487 = 3'h5 == encoders_5_io_output ? proc_5_io_next_header_25 : _GEN_3423; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3488 = 3'h5 == encoders_5_io_output ? proc_5_io_next_header_26 : _GEN_3424; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3489 = 3'h5 == encoders_5_io_output ? proc_5_io_next_header_27 : _GEN_3425; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3490 = 3'h5 == encoders_5_io_output ? proc_5_io_next_header_28 : _GEN_3426; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3491 = 3'h5 == encoders_5_io_output ? proc_5_io_next_header_29 : _GEN_3427; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3492 = 3'h5 == encoders_5_io_output ? proc_5_io_next_header_30 : _GEN_3428; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3493 = 3'h5 == encoders_5_io_output ? proc_5_io_next_header_31 : _GEN_3429; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3494 = 3'h5 == encoders_5_io_output ? proc_5_io_next_header_32 : _GEN_3430; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3495 = 3'h5 == encoders_5_io_output ? proc_5_io_next_header_33 : _GEN_3431; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3496 = 3'h5 == encoders_5_io_output ? proc_5_io_next_header_34 : _GEN_3432; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3497 = 3'h5 == encoders_5_io_output ? proc_5_io_next_header_35 : _GEN_3433; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3498 = 3'h5 == encoders_5_io_output ? proc_5_io_next_header_36 : _GEN_3434; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3499 = 3'h5 == encoders_5_io_output ? proc_5_io_next_header_37 : _GEN_3435; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3500 = 3'h5 == encoders_5_io_output ? proc_5_io_next_header_38 : _GEN_3436; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3501 = 3'h5 == encoders_5_io_output ? proc_5_io_next_header_39 : _GEN_3437; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3502 = 3'h5 == encoders_5_io_output ? proc_5_io_next_header_40 : _GEN_3438; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3503 = 3'h5 == encoders_5_io_output ? proc_5_io_next_header_41 : _GEN_3439; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3504 = 3'h5 == encoders_5_io_output ? proc_5_io_next_header_42 : _GEN_3440; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3505 = 3'h5 == encoders_5_io_output ? proc_5_io_next_header_43 : _GEN_3441; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3506 = 3'h5 == encoders_5_io_output ? proc_5_io_next_header_44 : _GEN_3442; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3507 = 3'h5 == encoders_5_io_output ? proc_5_io_next_header_45 : _GEN_3443; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3508 = 3'h5 == encoders_5_io_output ? proc_5_io_next_header_46 : _GEN_3444; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3509 = 3'h5 == encoders_5_io_output ? proc_5_io_next_header_47 : _GEN_3445; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3510 = 3'h5 == encoders_5_io_output ? proc_5_io_next_header_48 : _GEN_3446; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3511 = 3'h5 == encoders_5_io_output ? proc_5_io_next_header_49 : _GEN_3447; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3512 = 3'h5 == encoders_5_io_output ? proc_5_io_next_header_50 : _GEN_3448; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3513 = 3'h5 == encoders_5_io_output ? proc_5_io_next_header_51 : _GEN_3449; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3514 = 3'h5 == encoders_5_io_output ? proc_5_io_next_header_52 : _GEN_3450; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3515 = 3'h5 == encoders_5_io_output ? proc_5_io_next_header_53 : _GEN_3451; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3516 = 3'h5 == encoders_5_io_output ? proc_5_io_next_header_54 : _GEN_3452; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3517 = 3'h5 == encoders_5_io_output ? proc_5_io_next_header_55 : _GEN_3453; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3518 = 3'h5 == encoders_5_io_output ? proc_5_io_next_header_56 : _GEN_3454; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3519 = 3'h5 == encoders_5_io_output ? proc_5_io_next_header_57 : _GEN_3455; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3520 = 3'h5 == encoders_5_io_output ? proc_5_io_next_header_58 : _GEN_3456; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3521 = 3'h5 == encoders_5_io_output ? proc_5_io_next_header_59 : _GEN_3457; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3522 = 3'h5 == encoders_5_io_output ? proc_5_io_next_header_60 : _GEN_3458; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3523 = 3'h5 == encoders_5_io_output ? proc_5_io_next_header_61 : _GEN_3459; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3524 = 3'h5 == encoders_5_io_output ? proc_5_io_next_header_62 : _GEN_3460; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3525 = 3'h5 == encoders_5_io_output ? proc_5_io_next_header_63 : _GEN_3461; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3526 = 3'h6 == encoders_5_io_output ? proc_6_io_next_header_0 : _GEN_3462; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3527 = 3'h6 == encoders_5_io_output ? proc_6_io_next_header_1 : _GEN_3463; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3528 = 3'h6 == encoders_5_io_output ? proc_6_io_next_header_2 : _GEN_3464; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3529 = 3'h6 == encoders_5_io_output ? proc_6_io_next_header_3 : _GEN_3465; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3530 = 3'h6 == encoders_5_io_output ? proc_6_io_next_header_4 : _GEN_3466; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3531 = 3'h6 == encoders_5_io_output ? proc_6_io_next_header_5 : _GEN_3467; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3532 = 3'h6 == encoders_5_io_output ? proc_6_io_next_header_6 : _GEN_3468; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3533 = 3'h6 == encoders_5_io_output ? proc_6_io_next_header_7 : _GEN_3469; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3534 = 3'h6 == encoders_5_io_output ? proc_6_io_next_header_8 : _GEN_3470; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3535 = 3'h6 == encoders_5_io_output ? proc_6_io_next_header_9 : _GEN_3471; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3536 = 3'h6 == encoders_5_io_output ? proc_6_io_next_header_10 : _GEN_3472; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3537 = 3'h6 == encoders_5_io_output ? proc_6_io_next_header_11 : _GEN_3473; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3538 = 3'h6 == encoders_5_io_output ? proc_6_io_next_header_12 : _GEN_3474; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3539 = 3'h6 == encoders_5_io_output ? proc_6_io_next_header_13 : _GEN_3475; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3540 = 3'h6 == encoders_5_io_output ? proc_6_io_next_header_14 : _GEN_3476; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3541 = 3'h6 == encoders_5_io_output ? proc_6_io_next_header_15 : _GEN_3477; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3542 = 3'h6 == encoders_5_io_output ? proc_6_io_next_header_16 : _GEN_3478; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3543 = 3'h6 == encoders_5_io_output ? proc_6_io_next_header_17 : _GEN_3479; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3544 = 3'h6 == encoders_5_io_output ? proc_6_io_next_header_18 : _GEN_3480; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3545 = 3'h6 == encoders_5_io_output ? proc_6_io_next_header_19 : _GEN_3481; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3546 = 3'h6 == encoders_5_io_output ? proc_6_io_next_header_20 : _GEN_3482; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3547 = 3'h6 == encoders_5_io_output ? proc_6_io_next_header_21 : _GEN_3483; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3548 = 3'h6 == encoders_5_io_output ? proc_6_io_next_header_22 : _GEN_3484; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3549 = 3'h6 == encoders_5_io_output ? proc_6_io_next_header_23 : _GEN_3485; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3550 = 3'h6 == encoders_5_io_output ? proc_6_io_next_header_24 : _GEN_3486; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3551 = 3'h6 == encoders_5_io_output ? proc_6_io_next_header_25 : _GEN_3487; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3552 = 3'h6 == encoders_5_io_output ? proc_6_io_next_header_26 : _GEN_3488; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3553 = 3'h6 == encoders_5_io_output ? proc_6_io_next_header_27 : _GEN_3489; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3554 = 3'h6 == encoders_5_io_output ? proc_6_io_next_header_28 : _GEN_3490; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3555 = 3'h6 == encoders_5_io_output ? proc_6_io_next_header_29 : _GEN_3491; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3556 = 3'h6 == encoders_5_io_output ? proc_6_io_next_header_30 : _GEN_3492; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3557 = 3'h6 == encoders_5_io_output ? proc_6_io_next_header_31 : _GEN_3493; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3558 = 3'h6 == encoders_5_io_output ? proc_6_io_next_header_32 : _GEN_3494; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3559 = 3'h6 == encoders_5_io_output ? proc_6_io_next_header_33 : _GEN_3495; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3560 = 3'h6 == encoders_5_io_output ? proc_6_io_next_header_34 : _GEN_3496; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3561 = 3'h6 == encoders_5_io_output ? proc_6_io_next_header_35 : _GEN_3497; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3562 = 3'h6 == encoders_5_io_output ? proc_6_io_next_header_36 : _GEN_3498; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3563 = 3'h6 == encoders_5_io_output ? proc_6_io_next_header_37 : _GEN_3499; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3564 = 3'h6 == encoders_5_io_output ? proc_6_io_next_header_38 : _GEN_3500; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3565 = 3'h6 == encoders_5_io_output ? proc_6_io_next_header_39 : _GEN_3501; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3566 = 3'h6 == encoders_5_io_output ? proc_6_io_next_header_40 : _GEN_3502; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3567 = 3'h6 == encoders_5_io_output ? proc_6_io_next_header_41 : _GEN_3503; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3568 = 3'h6 == encoders_5_io_output ? proc_6_io_next_header_42 : _GEN_3504; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3569 = 3'h6 == encoders_5_io_output ? proc_6_io_next_header_43 : _GEN_3505; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3570 = 3'h6 == encoders_5_io_output ? proc_6_io_next_header_44 : _GEN_3506; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3571 = 3'h6 == encoders_5_io_output ? proc_6_io_next_header_45 : _GEN_3507; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3572 = 3'h6 == encoders_5_io_output ? proc_6_io_next_header_46 : _GEN_3508; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3573 = 3'h6 == encoders_5_io_output ? proc_6_io_next_header_47 : _GEN_3509; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3574 = 3'h6 == encoders_5_io_output ? proc_6_io_next_header_48 : _GEN_3510; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3575 = 3'h6 == encoders_5_io_output ? proc_6_io_next_header_49 : _GEN_3511; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3576 = 3'h6 == encoders_5_io_output ? proc_6_io_next_header_50 : _GEN_3512; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3577 = 3'h6 == encoders_5_io_output ? proc_6_io_next_header_51 : _GEN_3513; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3578 = 3'h6 == encoders_5_io_output ? proc_6_io_next_header_52 : _GEN_3514; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3579 = 3'h6 == encoders_5_io_output ? proc_6_io_next_header_53 : _GEN_3515; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3580 = 3'h6 == encoders_5_io_output ? proc_6_io_next_header_54 : _GEN_3516; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3581 = 3'h6 == encoders_5_io_output ? proc_6_io_next_header_55 : _GEN_3517; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3582 = 3'h6 == encoders_5_io_output ? proc_6_io_next_header_56 : _GEN_3518; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3583 = 3'h6 == encoders_5_io_output ? proc_6_io_next_header_57 : _GEN_3519; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3584 = 3'h6 == encoders_5_io_output ? proc_6_io_next_header_58 : _GEN_3520; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3585 = 3'h6 == encoders_5_io_output ? proc_6_io_next_header_59 : _GEN_3521; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3586 = 3'h6 == encoders_5_io_output ? proc_6_io_next_header_60 : _GEN_3522; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3587 = 3'h6 == encoders_5_io_output ? proc_6_io_next_header_61 : _GEN_3523; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3588 = 3'h6 == encoders_5_io_output ? proc_6_io_next_header_62 : _GEN_3524; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3589 = 3'h6 == encoders_5_io_output ? proc_6_io_next_header_63 : _GEN_3525; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3590 = 3'h7 == encoders_5_io_output ? proc_7_io_next_header_0 : _GEN_3526; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3591 = 3'h7 == encoders_5_io_output ? proc_7_io_next_header_1 : _GEN_3527; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3592 = 3'h7 == encoders_5_io_output ? proc_7_io_next_header_2 : _GEN_3528; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3593 = 3'h7 == encoders_5_io_output ? proc_7_io_next_header_3 : _GEN_3529; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3594 = 3'h7 == encoders_5_io_output ? proc_7_io_next_header_4 : _GEN_3530; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3595 = 3'h7 == encoders_5_io_output ? proc_7_io_next_header_5 : _GEN_3531; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3596 = 3'h7 == encoders_5_io_output ? proc_7_io_next_header_6 : _GEN_3532; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3597 = 3'h7 == encoders_5_io_output ? proc_7_io_next_header_7 : _GEN_3533; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3598 = 3'h7 == encoders_5_io_output ? proc_7_io_next_header_8 : _GEN_3534; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3599 = 3'h7 == encoders_5_io_output ? proc_7_io_next_header_9 : _GEN_3535; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3600 = 3'h7 == encoders_5_io_output ? proc_7_io_next_header_10 : _GEN_3536; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3601 = 3'h7 == encoders_5_io_output ? proc_7_io_next_header_11 : _GEN_3537; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3602 = 3'h7 == encoders_5_io_output ? proc_7_io_next_header_12 : _GEN_3538; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3603 = 3'h7 == encoders_5_io_output ? proc_7_io_next_header_13 : _GEN_3539; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3604 = 3'h7 == encoders_5_io_output ? proc_7_io_next_header_14 : _GEN_3540; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3605 = 3'h7 == encoders_5_io_output ? proc_7_io_next_header_15 : _GEN_3541; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3606 = 3'h7 == encoders_5_io_output ? proc_7_io_next_header_16 : _GEN_3542; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3607 = 3'h7 == encoders_5_io_output ? proc_7_io_next_header_17 : _GEN_3543; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3608 = 3'h7 == encoders_5_io_output ? proc_7_io_next_header_18 : _GEN_3544; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3609 = 3'h7 == encoders_5_io_output ? proc_7_io_next_header_19 : _GEN_3545; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3610 = 3'h7 == encoders_5_io_output ? proc_7_io_next_header_20 : _GEN_3546; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3611 = 3'h7 == encoders_5_io_output ? proc_7_io_next_header_21 : _GEN_3547; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3612 = 3'h7 == encoders_5_io_output ? proc_7_io_next_header_22 : _GEN_3548; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3613 = 3'h7 == encoders_5_io_output ? proc_7_io_next_header_23 : _GEN_3549; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3614 = 3'h7 == encoders_5_io_output ? proc_7_io_next_header_24 : _GEN_3550; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3615 = 3'h7 == encoders_5_io_output ? proc_7_io_next_header_25 : _GEN_3551; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3616 = 3'h7 == encoders_5_io_output ? proc_7_io_next_header_26 : _GEN_3552; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3617 = 3'h7 == encoders_5_io_output ? proc_7_io_next_header_27 : _GEN_3553; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3618 = 3'h7 == encoders_5_io_output ? proc_7_io_next_header_28 : _GEN_3554; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3619 = 3'h7 == encoders_5_io_output ? proc_7_io_next_header_29 : _GEN_3555; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3620 = 3'h7 == encoders_5_io_output ? proc_7_io_next_header_30 : _GEN_3556; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3621 = 3'h7 == encoders_5_io_output ? proc_7_io_next_header_31 : _GEN_3557; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3622 = 3'h7 == encoders_5_io_output ? proc_7_io_next_header_32 : _GEN_3558; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3623 = 3'h7 == encoders_5_io_output ? proc_7_io_next_header_33 : _GEN_3559; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3624 = 3'h7 == encoders_5_io_output ? proc_7_io_next_header_34 : _GEN_3560; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3625 = 3'h7 == encoders_5_io_output ? proc_7_io_next_header_35 : _GEN_3561; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3626 = 3'h7 == encoders_5_io_output ? proc_7_io_next_header_36 : _GEN_3562; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3627 = 3'h7 == encoders_5_io_output ? proc_7_io_next_header_37 : _GEN_3563; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3628 = 3'h7 == encoders_5_io_output ? proc_7_io_next_header_38 : _GEN_3564; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3629 = 3'h7 == encoders_5_io_output ? proc_7_io_next_header_39 : _GEN_3565; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3630 = 3'h7 == encoders_5_io_output ? proc_7_io_next_header_40 : _GEN_3566; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3631 = 3'h7 == encoders_5_io_output ? proc_7_io_next_header_41 : _GEN_3567; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3632 = 3'h7 == encoders_5_io_output ? proc_7_io_next_header_42 : _GEN_3568; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3633 = 3'h7 == encoders_5_io_output ? proc_7_io_next_header_43 : _GEN_3569; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3634 = 3'h7 == encoders_5_io_output ? proc_7_io_next_header_44 : _GEN_3570; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3635 = 3'h7 == encoders_5_io_output ? proc_7_io_next_header_45 : _GEN_3571; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3636 = 3'h7 == encoders_5_io_output ? proc_7_io_next_header_46 : _GEN_3572; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3637 = 3'h7 == encoders_5_io_output ? proc_7_io_next_header_47 : _GEN_3573; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3638 = 3'h7 == encoders_5_io_output ? proc_7_io_next_header_48 : _GEN_3574; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3639 = 3'h7 == encoders_5_io_output ? proc_7_io_next_header_49 : _GEN_3575; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3640 = 3'h7 == encoders_5_io_output ? proc_7_io_next_header_50 : _GEN_3576; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3641 = 3'h7 == encoders_5_io_output ? proc_7_io_next_header_51 : _GEN_3577; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3642 = 3'h7 == encoders_5_io_output ? proc_7_io_next_header_52 : _GEN_3578; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3643 = 3'h7 == encoders_5_io_output ? proc_7_io_next_header_53 : _GEN_3579; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3644 = 3'h7 == encoders_5_io_output ? proc_7_io_next_header_54 : _GEN_3580; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3645 = 3'h7 == encoders_5_io_output ? proc_7_io_next_header_55 : _GEN_3581; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3646 = 3'h7 == encoders_5_io_output ? proc_7_io_next_header_56 : _GEN_3582; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3647 = 3'h7 == encoders_5_io_output ? proc_7_io_next_header_57 : _GEN_3583; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3648 = 3'h7 == encoders_5_io_output ? proc_7_io_next_header_58 : _GEN_3584; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3649 = 3'h7 == encoders_5_io_output ? proc_7_io_next_header_59 : _GEN_3585; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3650 = 3'h7 == encoders_5_io_output ? proc_7_io_next_header_60 : _GEN_3586; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3651 = 3'h7 == encoders_5_io_output ? proc_7_io_next_header_61 : _GEN_3587; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3652 = 3'h7 == encoders_5_io_output ? proc_7_io_next_header_62 : _GEN_3588; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3653 = 3'h7 == encoders_5_io_output ? proc_7_io_next_header_63 : _GEN_3589; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3719 = 3'h0 == encoders_6_io_output ? proc_0_io_next_header_0 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3720 = 3'h0 == encoders_6_io_output ? proc_0_io_next_header_1 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3721 = 3'h0 == encoders_6_io_output ? proc_0_io_next_header_2 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3722 = 3'h0 == encoders_6_io_output ? proc_0_io_next_header_3 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3723 = 3'h0 == encoders_6_io_output ? proc_0_io_next_header_4 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3724 = 3'h0 == encoders_6_io_output ? proc_0_io_next_header_5 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3725 = 3'h0 == encoders_6_io_output ? proc_0_io_next_header_6 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3726 = 3'h0 == encoders_6_io_output ? proc_0_io_next_header_7 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3727 = 3'h0 == encoders_6_io_output ? proc_0_io_next_header_8 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3728 = 3'h0 == encoders_6_io_output ? proc_0_io_next_header_9 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3729 = 3'h0 == encoders_6_io_output ? proc_0_io_next_header_10 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3730 = 3'h0 == encoders_6_io_output ? proc_0_io_next_header_11 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3731 = 3'h0 == encoders_6_io_output ? proc_0_io_next_header_12 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3732 = 3'h0 == encoders_6_io_output ? proc_0_io_next_header_13 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3733 = 3'h0 == encoders_6_io_output ? proc_0_io_next_header_14 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3734 = 3'h0 == encoders_6_io_output ? proc_0_io_next_header_15 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3735 = 3'h0 == encoders_6_io_output ? proc_0_io_next_header_16 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3736 = 3'h0 == encoders_6_io_output ? proc_0_io_next_header_17 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3737 = 3'h0 == encoders_6_io_output ? proc_0_io_next_header_18 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3738 = 3'h0 == encoders_6_io_output ? proc_0_io_next_header_19 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3739 = 3'h0 == encoders_6_io_output ? proc_0_io_next_header_20 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3740 = 3'h0 == encoders_6_io_output ? proc_0_io_next_header_21 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3741 = 3'h0 == encoders_6_io_output ? proc_0_io_next_header_22 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3742 = 3'h0 == encoders_6_io_output ? proc_0_io_next_header_23 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3743 = 3'h0 == encoders_6_io_output ? proc_0_io_next_header_24 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3744 = 3'h0 == encoders_6_io_output ? proc_0_io_next_header_25 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3745 = 3'h0 == encoders_6_io_output ? proc_0_io_next_header_26 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3746 = 3'h0 == encoders_6_io_output ? proc_0_io_next_header_27 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3747 = 3'h0 == encoders_6_io_output ? proc_0_io_next_header_28 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3748 = 3'h0 == encoders_6_io_output ? proc_0_io_next_header_29 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3749 = 3'h0 == encoders_6_io_output ? proc_0_io_next_header_30 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3750 = 3'h0 == encoders_6_io_output ? proc_0_io_next_header_31 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3751 = 3'h0 == encoders_6_io_output ? proc_0_io_next_header_32 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3752 = 3'h0 == encoders_6_io_output ? proc_0_io_next_header_33 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3753 = 3'h0 == encoders_6_io_output ? proc_0_io_next_header_34 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3754 = 3'h0 == encoders_6_io_output ? proc_0_io_next_header_35 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3755 = 3'h0 == encoders_6_io_output ? proc_0_io_next_header_36 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3756 = 3'h0 == encoders_6_io_output ? proc_0_io_next_header_37 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3757 = 3'h0 == encoders_6_io_output ? proc_0_io_next_header_38 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3758 = 3'h0 == encoders_6_io_output ? proc_0_io_next_header_39 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3759 = 3'h0 == encoders_6_io_output ? proc_0_io_next_header_40 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3760 = 3'h0 == encoders_6_io_output ? proc_0_io_next_header_41 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3761 = 3'h0 == encoders_6_io_output ? proc_0_io_next_header_42 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3762 = 3'h0 == encoders_6_io_output ? proc_0_io_next_header_43 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3763 = 3'h0 == encoders_6_io_output ? proc_0_io_next_header_44 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3764 = 3'h0 == encoders_6_io_output ? proc_0_io_next_header_45 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3765 = 3'h0 == encoders_6_io_output ? proc_0_io_next_header_46 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3766 = 3'h0 == encoders_6_io_output ? proc_0_io_next_header_47 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3767 = 3'h0 == encoders_6_io_output ? proc_0_io_next_header_48 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3768 = 3'h0 == encoders_6_io_output ? proc_0_io_next_header_49 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3769 = 3'h0 == encoders_6_io_output ? proc_0_io_next_header_50 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3770 = 3'h0 == encoders_6_io_output ? proc_0_io_next_header_51 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3771 = 3'h0 == encoders_6_io_output ? proc_0_io_next_header_52 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3772 = 3'h0 == encoders_6_io_output ? proc_0_io_next_header_53 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3773 = 3'h0 == encoders_6_io_output ? proc_0_io_next_header_54 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3774 = 3'h0 == encoders_6_io_output ? proc_0_io_next_header_55 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3775 = 3'h0 == encoders_6_io_output ? proc_0_io_next_header_56 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3776 = 3'h0 == encoders_6_io_output ? proc_0_io_next_header_57 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3777 = 3'h0 == encoders_6_io_output ? proc_0_io_next_header_58 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3778 = 3'h0 == encoders_6_io_output ? proc_0_io_next_header_59 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3779 = 3'h0 == encoders_6_io_output ? proc_0_io_next_header_60 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3780 = 3'h0 == encoders_6_io_output ? proc_0_io_next_header_61 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3781 = 3'h0 == encoders_6_io_output ? proc_0_io_next_header_62 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3782 = 3'h0 == encoders_6_io_output ? proc_0_io_next_header_63 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_3783 = 3'h1 == encoders_6_io_output ? proc_1_io_next_header_0 : _GEN_3719; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3784 = 3'h1 == encoders_6_io_output ? proc_1_io_next_header_1 : _GEN_3720; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3785 = 3'h1 == encoders_6_io_output ? proc_1_io_next_header_2 : _GEN_3721; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3786 = 3'h1 == encoders_6_io_output ? proc_1_io_next_header_3 : _GEN_3722; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3787 = 3'h1 == encoders_6_io_output ? proc_1_io_next_header_4 : _GEN_3723; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3788 = 3'h1 == encoders_6_io_output ? proc_1_io_next_header_5 : _GEN_3724; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3789 = 3'h1 == encoders_6_io_output ? proc_1_io_next_header_6 : _GEN_3725; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3790 = 3'h1 == encoders_6_io_output ? proc_1_io_next_header_7 : _GEN_3726; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3791 = 3'h1 == encoders_6_io_output ? proc_1_io_next_header_8 : _GEN_3727; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3792 = 3'h1 == encoders_6_io_output ? proc_1_io_next_header_9 : _GEN_3728; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3793 = 3'h1 == encoders_6_io_output ? proc_1_io_next_header_10 : _GEN_3729; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3794 = 3'h1 == encoders_6_io_output ? proc_1_io_next_header_11 : _GEN_3730; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3795 = 3'h1 == encoders_6_io_output ? proc_1_io_next_header_12 : _GEN_3731; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3796 = 3'h1 == encoders_6_io_output ? proc_1_io_next_header_13 : _GEN_3732; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3797 = 3'h1 == encoders_6_io_output ? proc_1_io_next_header_14 : _GEN_3733; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3798 = 3'h1 == encoders_6_io_output ? proc_1_io_next_header_15 : _GEN_3734; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3799 = 3'h1 == encoders_6_io_output ? proc_1_io_next_header_16 : _GEN_3735; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3800 = 3'h1 == encoders_6_io_output ? proc_1_io_next_header_17 : _GEN_3736; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3801 = 3'h1 == encoders_6_io_output ? proc_1_io_next_header_18 : _GEN_3737; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3802 = 3'h1 == encoders_6_io_output ? proc_1_io_next_header_19 : _GEN_3738; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3803 = 3'h1 == encoders_6_io_output ? proc_1_io_next_header_20 : _GEN_3739; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3804 = 3'h1 == encoders_6_io_output ? proc_1_io_next_header_21 : _GEN_3740; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3805 = 3'h1 == encoders_6_io_output ? proc_1_io_next_header_22 : _GEN_3741; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3806 = 3'h1 == encoders_6_io_output ? proc_1_io_next_header_23 : _GEN_3742; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3807 = 3'h1 == encoders_6_io_output ? proc_1_io_next_header_24 : _GEN_3743; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3808 = 3'h1 == encoders_6_io_output ? proc_1_io_next_header_25 : _GEN_3744; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3809 = 3'h1 == encoders_6_io_output ? proc_1_io_next_header_26 : _GEN_3745; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3810 = 3'h1 == encoders_6_io_output ? proc_1_io_next_header_27 : _GEN_3746; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3811 = 3'h1 == encoders_6_io_output ? proc_1_io_next_header_28 : _GEN_3747; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3812 = 3'h1 == encoders_6_io_output ? proc_1_io_next_header_29 : _GEN_3748; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3813 = 3'h1 == encoders_6_io_output ? proc_1_io_next_header_30 : _GEN_3749; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3814 = 3'h1 == encoders_6_io_output ? proc_1_io_next_header_31 : _GEN_3750; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3815 = 3'h1 == encoders_6_io_output ? proc_1_io_next_header_32 : _GEN_3751; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3816 = 3'h1 == encoders_6_io_output ? proc_1_io_next_header_33 : _GEN_3752; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3817 = 3'h1 == encoders_6_io_output ? proc_1_io_next_header_34 : _GEN_3753; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3818 = 3'h1 == encoders_6_io_output ? proc_1_io_next_header_35 : _GEN_3754; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3819 = 3'h1 == encoders_6_io_output ? proc_1_io_next_header_36 : _GEN_3755; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3820 = 3'h1 == encoders_6_io_output ? proc_1_io_next_header_37 : _GEN_3756; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3821 = 3'h1 == encoders_6_io_output ? proc_1_io_next_header_38 : _GEN_3757; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3822 = 3'h1 == encoders_6_io_output ? proc_1_io_next_header_39 : _GEN_3758; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3823 = 3'h1 == encoders_6_io_output ? proc_1_io_next_header_40 : _GEN_3759; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3824 = 3'h1 == encoders_6_io_output ? proc_1_io_next_header_41 : _GEN_3760; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3825 = 3'h1 == encoders_6_io_output ? proc_1_io_next_header_42 : _GEN_3761; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3826 = 3'h1 == encoders_6_io_output ? proc_1_io_next_header_43 : _GEN_3762; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3827 = 3'h1 == encoders_6_io_output ? proc_1_io_next_header_44 : _GEN_3763; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3828 = 3'h1 == encoders_6_io_output ? proc_1_io_next_header_45 : _GEN_3764; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3829 = 3'h1 == encoders_6_io_output ? proc_1_io_next_header_46 : _GEN_3765; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3830 = 3'h1 == encoders_6_io_output ? proc_1_io_next_header_47 : _GEN_3766; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3831 = 3'h1 == encoders_6_io_output ? proc_1_io_next_header_48 : _GEN_3767; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3832 = 3'h1 == encoders_6_io_output ? proc_1_io_next_header_49 : _GEN_3768; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3833 = 3'h1 == encoders_6_io_output ? proc_1_io_next_header_50 : _GEN_3769; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3834 = 3'h1 == encoders_6_io_output ? proc_1_io_next_header_51 : _GEN_3770; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3835 = 3'h1 == encoders_6_io_output ? proc_1_io_next_header_52 : _GEN_3771; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3836 = 3'h1 == encoders_6_io_output ? proc_1_io_next_header_53 : _GEN_3772; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3837 = 3'h1 == encoders_6_io_output ? proc_1_io_next_header_54 : _GEN_3773; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3838 = 3'h1 == encoders_6_io_output ? proc_1_io_next_header_55 : _GEN_3774; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3839 = 3'h1 == encoders_6_io_output ? proc_1_io_next_header_56 : _GEN_3775; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3840 = 3'h1 == encoders_6_io_output ? proc_1_io_next_header_57 : _GEN_3776; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3841 = 3'h1 == encoders_6_io_output ? proc_1_io_next_header_58 : _GEN_3777; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3842 = 3'h1 == encoders_6_io_output ? proc_1_io_next_header_59 : _GEN_3778; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3843 = 3'h1 == encoders_6_io_output ? proc_1_io_next_header_60 : _GEN_3779; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3844 = 3'h1 == encoders_6_io_output ? proc_1_io_next_header_61 : _GEN_3780; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3845 = 3'h1 == encoders_6_io_output ? proc_1_io_next_header_62 : _GEN_3781; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3846 = 3'h1 == encoders_6_io_output ? proc_1_io_next_header_63 : _GEN_3782; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3847 = 3'h2 == encoders_6_io_output ? proc_2_io_next_header_0 : _GEN_3783; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3848 = 3'h2 == encoders_6_io_output ? proc_2_io_next_header_1 : _GEN_3784; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3849 = 3'h2 == encoders_6_io_output ? proc_2_io_next_header_2 : _GEN_3785; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3850 = 3'h2 == encoders_6_io_output ? proc_2_io_next_header_3 : _GEN_3786; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3851 = 3'h2 == encoders_6_io_output ? proc_2_io_next_header_4 : _GEN_3787; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3852 = 3'h2 == encoders_6_io_output ? proc_2_io_next_header_5 : _GEN_3788; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3853 = 3'h2 == encoders_6_io_output ? proc_2_io_next_header_6 : _GEN_3789; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3854 = 3'h2 == encoders_6_io_output ? proc_2_io_next_header_7 : _GEN_3790; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3855 = 3'h2 == encoders_6_io_output ? proc_2_io_next_header_8 : _GEN_3791; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3856 = 3'h2 == encoders_6_io_output ? proc_2_io_next_header_9 : _GEN_3792; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3857 = 3'h2 == encoders_6_io_output ? proc_2_io_next_header_10 : _GEN_3793; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3858 = 3'h2 == encoders_6_io_output ? proc_2_io_next_header_11 : _GEN_3794; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3859 = 3'h2 == encoders_6_io_output ? proc_2_io_next_header_12 : _GEN_3795; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3860 = 3'h2 == encoders_6_io_output ? proc_2_io_next_header_13 : _GEN_3796; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3861 = 3'h2 == encoders_6_io_output ? proc_2_io_next_header_14 : _GEN_3797; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3862 = 3'h2 == encoders_6_io_output ? proc_2_io_next_header_15 : _GEN_3798; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3863 = 3'h2 == encoders_6_io_output ? proc_2_io_next_header_16 : _GEN_3799; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3864 = 3'h2 == encoders_6_io_output ? proc_2_io_next_header_17 : _GEN_3800; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3865 = 3'h2 == encoders_6_io_output ? proc_2_io_next_header_18 : _GEN_3801; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3866 = 3'h2 == encoders_6_io_output ? proc_2_io_next_header_19 : _GEN_3802; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3867 = 3'h2 == encoders_6_io_output ? proc_2_io_next_header_20 : _GEN_3803; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3868 = 3'h2 == encoders_6_io_output ? proc_2_io_next_header_21 : _GEN_3804; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3869 = 3'h2 == encoders_6_io_output ? proc_2_io_next_header_22 : _GEN_3805; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3870 = 3'h2 == encoders_6_io_output ? proc_2_io_next_header_23 : _GEN_3806; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3871 = 3'h2 == encoders_6_io_output ? proc_2_io_next_header_24 : _GEN_3807; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3872 = 3'h2 == encoders_6_io_output ? proc_2_io_next_header_25 : _GEN_3808; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3873 = 3'h2 == encoders_6_io_output ? proc_2_io_next_header_26 : _GEN_3809; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3874 = 3'h2 == encoders_6_io_output ? proc_2_io_next_header_27 : _GEN_3810; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3875 = 3'h2 == encoders_6_io_output ? proc_2_io_next_header_28 : _GEN_3811; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3876 = 3'h2 == encoders_6_io_output ? proc_2_io_next_header_29 : _GEN_3812; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3877 = 3'h2 == encoders_6_io_output ? proc_2_io_next_header_30 : _GEN_3813; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3878 = 3'h2 == encoders_6_io_output ? proc_2_io_next_header_31 : _GEN_3814; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3879 = 3'h2 == encoders_6_io_output ? proc_2_io_next_header_32 : _GEN_3815; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3880 = 3'h2 == encoders_6_io_output ? proc_2_io_next_header_33 : _GEN_3816; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3881 = 3'h2 == encoders_6_io_output ? proc_2_io_next_header_34 : _GEN_3817; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3882 = 3'h2 == encoders_6_io_output ? proc_2_io_next_header_35 : _GEN_3818; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3883 = 3'h2 == encoders_6_io_output ? proc_2_io_next_header_36 : _GEN_3819; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3884 = 3'h2 == encoders_6_io_output ? proc_2_io_next_header_37 : _GEN_3820; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3885 = 3'h2 == encoders_6_io_output ? proc_2_io_next_header_38 : _GEN_3821; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3886 = 3'h2 == encoders_6_io_output ? proc_2_io_next_header_39 : _GEN_3822; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3887 = 3'h2 == encoders_6_io_output ? proc_2_io_next_header_40 : _GEN_3823; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3888 = 3'h2 == encoders_6_io_output ? proc_2_io_next_header_41 : _GEN_3824; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3889 = 3'h2 == encoders_6_io_output ? proc_2_io_next_header_42 : _GEN_3825; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3890 = 3'h2 == encoders_6_io_output ? proc_2_io_next_header_43 : _GEN_3826; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3891 = 3'h2 == encoders_6_io_output ? proc_2_io_next_header_44 : _GEN_3827; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3892 = 3'h2 == encoders_6_io_output ? proc_2_io_next_header_45 : _GEN_3828; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3893 = 3'h2 == encoders_6_io_output ? proc_2_io_next_header_46 : _GEN_3829; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3894 = 3'h2 == encoders_6_io_output ? proc_2_io_next_header_47 : _GEN_3830; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3895 = 3'h2 == encoders_6_io_output ? proc_2_io_next_header_48 : _GEN_3831; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3896 = 3'h2 == encoders_6_io_output ? proc_2_io_next_header_49 : _GEN_3832; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3897 = 3'h2 == encoders_6_io_output ? proc_2_io_next_header_50 : _GEN_3833; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3898 = 3'h2 == encoders_6_io_output ? proc_2_io_next_header_51 : _GEN_3834; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3899 = 3'h2 == encoders_6_io_output ? proc_2_io_next_header_52 : _GEN_3835; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3900 = 3'h2 == encoders_6_io_output ? proc_2_io_next_header_53 : _GEN_3836; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3901 = 3'h2 == encoders_6_io_output ? proc_2_io_next_header_54 : _GEN_3837; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3902 = 3'h2 == encoders_6_io_output ? proc_2_io_next_header_55 : _GEN_3838; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3903 = 3'h2 == encoders_6_io_output ? proc_2_io_next_header_56 : _GEN_3839; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3904 = 3'h2 == encoders_6_io_output ? proc_2_io_next_header_57 : _GEN_3840; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3905 = 3'h2 == encoders_6_io_output ? proc_2_io_next_header_58 : _GEN_3841; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3906 = 3'h2 == encoders_6_io_output ? proc_2_io_next_header_59 : _GEN_3842; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3907 = 3'h2 == encoders_6_io_output ? proc_2_io_next_header_60 : _GEN_3843; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3908 = 3'h2 == encoders_6_io_output ? proc_2_io_next_header_61 : _GEN_3844; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3909 = 3'h2 == encoders_6_io_output ? proc_2_io_next_header_62 : _GEN_3845; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3910 = 3'h2 == encoders_6_io_output ? proc_2_io_next_header_63 : _GEN_3846; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3911 = 3'h3 == encoders_6_io_output ? proc_3_io_next_header_0 : _GEN_3847; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3912 = 3'h3 == encoders_6_io_output ? proc_3_io_next_header_1 : _GEN_3848; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3913 = 3'h3 == encoders_6_io_output ? proc_3_io_next_header_2 : _GEN_3849; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3914 = 3'h3 == encoders_6_io_output ? proc_3_io_next_header_3 : _GEN_3850; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3915 = 3'h3 == encoders_6_io_output ? proc_3_io_next_header_4 : _GEN_3851; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3916 = 3'h3 == encoders_6_io_output ? proc_3_io_next_header_5 : _GEN_3852; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3917 = 3'h3 == encoders_6_io_output ? proc_3_io_next_header_6 : _GEN_3853; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3918 = 3'h3 == encoders_6_io_output ? proc_3_io_next_header_7 : _GEN_3854; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3919 = 3'h3 == encoders_6_io_output ? proc_3_io_next_header_8 : _GEN_3855; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3920 = 3'h3 == encoders_6_io_output ? proc_3_io_next_header_9 : _GEN_3856; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3921 = 3'h3 == encoders_6_io_output ? proc_3_io_next_header_10 : _GEN_3857; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3922 = 3'h3 == encoders_6_io_output ? proc_3_io_next_header_11 : _GEN_3858; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3923 = 3'h3 == encoders_6_io_output ? proc_3_io_next_header_12 : _GEN_3859; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3924 = 3'h3 == encoders_6_io_output ? proc_3_io_next_header_13 : _GEN_3860; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3925 = 3'h3 == encoders_6_io_output ? proc_3_io_next_header_14 : _GEN_3861; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3926 = 3'h3 == encoders_6_io_output ? proc_3_io_next_header_15 : _GEN_3862; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3927 = 3'h3 == encoders_6_io_output ? proc_3_io_next_header_16 : _GEN_3863; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3928 = 3'h3 == encoders_6_io_output ? proc_3_io_next_header_17 : _GEN_3864; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3929 = 3'h3 == encoders_6_io_output ? proc_3_io_next_header_18 : _GEN_3865; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3930 = 3'h3 == encoders_6_io_output ? proc_3_io_next_header_19 : _GEN_3866; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3931 = 3'h3 == encoders_6_io_output ? proc_3_io_next_header_20 : _GEN_3867; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3932 = 3'h3 == encoders_6_io_output ? proc_3_io_next_header_21 : _GEN_3868; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3933 = 3'h3 == encoders_6_io_output ? proc_3_io_next_header_22 : _GEN_3869; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3934 = 3'h3 == encoders_6_io_output ? proc_3_io_next_header_23 : _GEN_3870; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3935 = 3'h3 == encoders_6_io_output ? proc_3_io_next_header_24 : _GEN_3871; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3936 = 3'h3 == encoders_6_io_output ? proc_3_io_next_header_25 : _GEN_3872; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3937 = 3'h3 == encoders_6_io_output ? proc_3_io_next_header_26 : _GEN_3873; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3938 = 3'h3 == encoders_6_io_output ? proc_3_io_next_header_27 : _GEN_3874; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3939 = 3'h3 == encoders_6_io_output ? proc_3_io_next_header_28 : _GEN_3875; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3940 = 3'h3 == encoders_6_io_output ? proc_3_io_next_header_29 : _GEN_3876; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3941 = 3'h3 == encoders_6_io_output ? proc_3_io_next_header_30 : _GEN_3877; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3942 = 3'h3 == encoders_6_io_output ? proc_3_io_next_header_31 : _GEN_3878; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3943 = 3'h3 == encoders_6_io_output ? proc_3_io_next_header_32 : _GEN_3879; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3944 = 3'h3 == encoders_6_io_output ? proc_3_io_next_header_33 : _GEN_3880; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3945 = 3'h3 == encoders_6_io_output ? proc_3_io_next_header_34 : _GEN_3881; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3946 = 3'h3 == encoders_6_io_output ? proc_3_io_next_header_35 : _GEN_3882; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3947 = 3'h3 == encoders_6_io_output ? proc_3_io_next_header_36 : _GEN_3883; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3948 = 3'h3 == encoders_6_io_output ? proc_3_io_next_header_37 : _GEN_3884; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3949 = 3'h3 == encoders_6_io_output ? proc_3_io_next_header_38 : _GEN_3885; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3950 = 3'h3 == encoders_6_io_output ? proc_3_io_next_header_39 : _GEN_3886; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3951 = 3'h3 == encoders_6_io_output ? proc_3_io_next_header_40 : _GEN_3887; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3952 = 3'h3 == encoders_6_io_output ? proc_3_io_next_header_41 : _GEN_3888; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3953 = 3'h3 == encoders_6_io_output ? proc_3_io_next_header_42 : _GEN_3889; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3954 = 3'h3 == encoders_6_io_output ? proc_3_io_next_header_43 : _GEN_3890; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3955 = 3'h3 == encoders_6_io_output ? proc_3_io_next_header_44 : _GEN_3891; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3956 = 3'h3 == encoders_6_io_output ? proc_3_io_next_header_45 : _GEN_3892; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3957 = 3'h3 == encoders_6_io_output ? proc_3_io_next_header_46 : _GEN_3893; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3958 = 3'h3 == encoders_6_io_output ? proc_3_io_next_header_47 : _GEN_3894; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3959 = 3'h3 == encoders_6_io_output ? proc_3_io_next_header_48 : _GEN_3895; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3960 = 3'h3 == encoders_6_io_output ? proc_3_io_next_header_49 : _GEN_3896; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3961 = 3'h3 == encoders_6_io_output ? proc_3_io_next_header_50 : _GEN_3897; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3962 = 3'h3 == encoders_6_io_output ? proc_3_io_next_header_51 : _GEN_3898; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3963 = 3'h3 == encoders_6_io_output ? proc_3_io_next_header_52 : _GEN_3899; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3964 = 3'h3 == encoders_6_io_output ? proc_3_io_next_header_53 : _GEN_3900; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3965 = 3'h3 == encoders_6_io_output ? proc_3_io_next_header_54 : _GEN_3901; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3966 = 3'h3 == encoders_6_io_output ? proc_3_io_next_header_55 : _GEN_3902; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3967 = 3'h3 == encoders_6_io_output ? proc_3_io_next_header_56 : _GEN_3903; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3968 = 3'h3 == encoders_6_io_output ? proc_3_io_next_header_57 : _GEN_3904; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3969 = 3'h3 == encoders_6_io_output ? proc_3_io_next_header_58 : _GEN_3905; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3970 = 3'h3 == encoders_6_io_output ? proc_3_io_next_header_59 : _GEN_3906; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3971 = 3'h3 == encoders_6_io_output ? proc_3_io_next_header_60 : _GEN_3907; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3972 = 3'h3 == encoders_6_io_output ? proc_3_io_next_header_61 : _GEN_3908; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3973 = 3'h3 == encoders_6_io_output ? proc_3_io_next_header_62 : _GEN_3909; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3974 = 3'h3 == encoders_6_io_output ? proc_3_io_next_header_63 : _GEN_3910; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3975 = 3'h4 == encoders_6_io_output ? proc_4_io_next_header_0 : _GEN_3911; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3976 = 3'h4 == encoders_6_io_output ? proc_4_io_next_header_1 : _GEN_3912; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3977 = 3'h4 == encoders_6_io_output ? proc_4_io_next_header_2 : _GEN_3913; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3978 = 3'h4 == encoders_6_io_output ? proc_4_io_next_header_3 : _GEN_3914; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3979 = 3'h4 == encoders_6_io_output ? proc_4_io_next_header_4 : _GEN_3915; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3980 = 3'h4 == encoders_6_io_output ? proc_4_io_next_header_5 : _GEN_3916; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3981 = 3'h4 == encoders_6_io_output ? proc_4_io_next_header_6 : _GEN_3917; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3982 = 3'h4 == encoders_6_io_output ? proc_4_io_next_header_7 : _GEN_3918; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3983 = 3'h4 == encoders_6_io_output ? proc_4_io_next_header_8 : _GEN_3919; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3984 = 3'h4 == encoders_6_io_output ? proc_4_io_next_header_9 : _GEN_3920; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3985 = 3'h4 == encoders_6_io_output ? proc_4_io_next_header_10 : _GEN_3921; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3986 = 3'h4 == encoders_6_io_output ? proc_4_io_next_header_11 : _GEN_3922; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3987 = 3'h4 == encoders_6_io_output ? proc_4_io_next_header_12 : _GEN_3923; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3988 = 3'h4 == encoders_6_io_output ? proc_4_io_next_header_13 : _GEN_3924; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3989 = 3'h4 == encoders_6_io_output ? proc_4_io_next_header_14 : _GEN_3925; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3990 = 3'h4 == encoders_6_io_output ? proc_4_io_next_header_15 : _GEN_3926; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3991 = 3'h4 == encoders_6_io_output ? proc_4_io_next_header_16 : _GEN_3927; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3992 = 3'h4 == encoders_6_io_output ? proc_4_io_next_header_17 : _GEN_3928; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3993 = 3'h4 == encoders_6_io_output ? proc_4_io_next_header_18 : _GEN_3929; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3994 = 3'h4 == encoders_6_io_output ? proc_4_io_next_header_19 : _GEN_3930; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3995 = 3'h4 == encoders_6_io_output ? proc_4_io_next_header_20 : _GEN_3931; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3996 = 3'h4 == encoders_6_io_output ? proc_4_io_next_header_21 : _GEN_3932; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3997 = 3'h4 == encoders_6_io_output ? proc_4_io_next_header_22 : _GEN_3933; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3998 = 3'h4 == encoders_6_io_output ? proc_4_io_next_header_23 : _GEN_3934; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_3999 = 3'h4 == encoders_6_io_output ? proc_4_io_next_header_24 : _GEN_3935; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4000 = 3'h4 == encoders_6_io_output ? proc_4_io_next_header_25 : _GEN_3936; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4001 = 3'h4 == encoders_6_io_output ? proc_4_io_next_header_26 : _GEN_3937; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4002 = 3'h4 == encoders_6_io_output ? proc_4_io_next_header_27 : _GEN_3938; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4003 = 3'h4 == encoders_6_io_output ? proc_4_io_next_header_28 : _GEN_3939; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4004 = 3'h4 == encoders_6_io_output ? proc_4_io_next_header_29 : _GEN_3940; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4005 = 3'h4 == encoders_6_io_output ? proc_4_io_next_header_30 : _GEN_3941; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4006 = 3'h4 == encoders_6_io_output ? proc_4_io_next_header_31 : _GEN_3942; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4007 = 3'h4 == encoders_6_io_output ? proc_4_io_next_header_32 : _GEN_3943; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4008 = 3'h4 == encoders_6_io_output ? proc_4_io_next_header_33 : _GEN_3944; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4009 = 3'h4 == encoders_6_io_output ? proc_4_io_next_header_34 : _GEN_3945; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4010 = 3'h4 == encoders_6_io_output ? proc_4_io_next_header_35 : _GEN_3946; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4011 = 3'h4 == encoders_6_io_output ? proc_4_io_next_header_36 : _GEN_3947; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4012 = 3'h4 == encoders_6_io_output ? proc_4_io_next_header_37 : _GEN_3948; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4013 = 3'h4 == encoders_6_io_output ? proc_4_io_next_header_38 : _GEN_3949; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4014 = 3'h4 == encoders_6_io_output ? proc_4_io_next_header_39 : _GEN_3950; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4015 = 3'h4 == encoders_6_io_output ? proc_4_io_next_header_40 : _GEN_3951; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4016 = 3'h4 == encoders_6_io_output ? proc_4_io_next_header_41 : _GEN_3952; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4017 = 3'h4 == encoders_6_io_output ? proc_4_io_next_header_42 : _GEN_3953; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4018 = 3'h4 == encoders_6_io_output ? proc_4_io_next_header_43 : _GEN_3954; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4019 = 3'h4 == encoders_6_io_output ? proc_4_io_next_header_44 : _GEN_3955; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4020 = 3'h4 == encoders_6_io_output ? proc_4_io_next_header_45 : _GEN_3956; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4021 = 3'h4 == encoders_6_io_output ? proc_4_io_next_header_46 : _GEN_3957; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4022 = 3'h4 == encoders_6_io_output ? proc_4_io_next_header_47 : _GEN_3958; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4023 = 3'h4 == encoders_6_io_output ? proc_4_io_next_header_48 : _GEN_3959; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4024 = 3'h4 == encoders_6_io_output ? proc_4_io_next_header_49 : _GEN_3960; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4025 = 3'h4 == encoders_6_io_output ? proc_4_io_next_header_50 : _GEN_3961; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4026 = 3'h4 == encoders_6_io_output ? proc_4_io_next_header_51 : _GEN_3962; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4027 = 3'h4 == encoders_6_io_output ? proc_4_io_next_header_52 : _GEN_3963; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4028 = 3'h4 == encoders_6_io_output ? proc_4_io_next_header_53 : _GEN_3964; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4029 = 3'h4 == encoders_6_io_output ? proc_4_io_next_header_54 : _GEN_3965; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4030 = 3'h4 == encoders_6_io_output ? proc_4_io_next_header_55 : _GEN_3966; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4031 = 3'h4 == encoders_6_io_output ? proc_4_io_next_header_56 : _GEN_3967; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4032 = 3'h4 == encoders_6_io_output ? proc_4_io_next_header_57 : _GEN_3968; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4033 = 3'h4 == encoders_6_io_output ? proc_4_io_next_header_58 : _GEN_3969; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4034 = 3'h4 == encoders_6_io_output ? proc_4_io_next_header_59 : _GEN_3970; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4035 = 3'h4 == encoders_6_io_output ? proc_4_io_next_header_60 : _GEN_3971; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4036 = 3'h4 == encoders_6_io_output ? proc_4_io_next_header_61 : _GEN_3972; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4037 = 3'h4 == encoders_6_io_output ? proc_4_io_next_header_62 : _GEN_3973; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4038 = 3'h4 == encoders_6_io_output ? proc_4_io_next_header_63 : _GEN_3974; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4039 = 3'h5 == encoders_6_io_output ? proc_5_io_next_header_0 : _GEN_3975; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4040 = 3'h5 == encoders_6_io_output ? proc_5_io_next_header_1 : _GEN_3976; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4041 = 3'h5 == encoders_6_io_output ? proc_5_io_next_header_2 : _GEN_3977; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4042 = 3'h5 == encoders_6_io_output ? proc_5_io_next_header_3 : _GEN_3978; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4043 = 3'h5 == encoders_6_io_output ? proc_5_io_next_header_4 : _GEN_3979; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4044 = 3'h5 == encoders_6_io_output ? proc_5_io_next_header_5 : _GEN_3980; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4045 = 3'h5 == encoders_6_io_output ? proc_5_io_next_header_6 : _GEN_3981; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4046 = 3'h5 == encoders_6_io_output ? proc_5_io_next_header_7 : _GEN_3982; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4047 = 3'h5 == encoders_6_io_output ? proc_5_io_next_header_8 : _GEN_3983; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4048 = 3'h5 == encoders_6_io_output ? proc_5_io_next_header_9 : _GEN_3984; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4049 = 3'h5 == encoders_6_io_output ? proc_5_io_next_header_10 : _GEN_3985; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4050 = 3'h5 == encoders_6_io_output ? proc_5_io_next_header_11 : _GEN_3986; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4051 = 3'h5 == encoders_6_io_output ? proc_5_io_next_header_12 : _GEN_3987; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4052 = 3'h5 == encoders_6_io_output ? proc_5_io_next_header_13 : _GEN_3988; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4053 = 3'h5 == encoders_6_io_output ? proc_5_io_next_header_14 : _GEN_3989; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4054 = 3'h5 == encoders_6_io_output ? proc_5_io_next_header_15 : _GEN_3990; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4055 = 3'h5 == encoders_6_io_output ? proc_5_io_next_header_16 : _GEN_3991; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4056 = 3'h5 == encoders_6_io_output ? proc_5_io_next_header_17 : _GEN_3992; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4057 = 3'h5 == encoders_6_io_output ? proc_5_io_next_header_18 : _GEN_3993; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4058 = 3'h5 == encoders_6_io_output ? proc_5_io_next_header_19 : _GEN_3994; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4059 = 3'h5 == encoders_6_io_output ? proc_5_io_next_header_20 : _GEN_3995; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4060 = 3'h5 == encoders_6_io_output ? proc_5_io_next_header_21 : _GEN_3996; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4061 = 3'h5 == encoders_6_io_output ? proc_5_io_next_header_22 : _GEN_3997; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4062 = 3'h5 == encoders_6_io_output ? proc_5_io_next_header_23 : _GEN_3998; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4063 = 3'h5 == encoders_6_io_output ? proc_5_io_next_header_24 : _GEN_3999; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4064 = 3'h5 == encoders_6_io_output ? proc_5_io_next_header_25 : _GEN_4000; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4065 = 3'h5 == encoders_6_io_output ? proc_5_io_next_header_26 : _GEN_4001; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4066 = 3'h5 == encoders_6_io_output ? proc_5_io_next_header_27 : _GEN_4002; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4067 = 3'h5 == encoders_6_io_output ? proc_5_io_next_header_28 : _GEN_4003; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4068 = 3'h5 == encoders_6_io_output ? proc_5_io_next_header_29 : _GEN_4004; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4069 = 3'h5 == encoders_6_io_output ? proc_5_io_next_header_30 : _GEN_4005; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4070 = 3'h5 == encoders_6_io_output ? proc_5_io_next_header_31 : _GEN_4006; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4071 = 3'h5 == encoders_6_io_output ? proc_5_io_next_header_32 : _GEN_4007; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4072 = 3'h5 == encoders_6_io_output ? proc_5_io_next_header_33 : _GEN_4008; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4073 = 3'h5 == encoders_6_io_output ? proc_5_io_next_header_34 : _GEN_4009; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4074 = 3'h5 == encoders_6_io_output ? proc_5_io_next_header_35 : _GEN_4010; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4075 = 3'h5 == encoders_6_io_output ? proc_5_io_next_header_36 : _GEN_4011; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4076 = 3'h5 == encoders_6_io_output ? proc_5_io_next_header_37 : _GEN_4012; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4077 = 3'h5 == encoders_6_io_output ? proc_5_io_next_header_38 : _GEN_4013; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4078 = 3'h5 == encoders_6_io_output ? proc_5_io_next_header_39 : _GEN_4014; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4079 = 3'h5 == encoders_6_io_output ? proc_5_io_next_header_40 : _GEN_4015; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4080 = 3'h5 == encoders_6_io_output ? proc_5_io_next_header_41 : _GEN_4016; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4081 = 3'h5 == encoders_6_io_output ? proc_5_io_next_header_42 : _GEN_4017; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4082 = 3'h5 == encoders_6_io_output ? proc_5_io_next_header_43 : _GEN_4018; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4083 = 3'h5 == encoders_6_io_output ? proc_5_io_next_header_44 : _GEN_4019; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4084 = 3'h5 == encoders_6_io_output ? proc_5_io_next_header_45 : _GEN_4020; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4085 = 3'h5 == encoders_6_io_output ? proc_5_io_next_header_46 : _GEN_4021; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4086 = 3'h5 == encoders_6_io_output ? proc_5_io_next_header_47 : _GEN_4022; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4087 = 3'h5 == encoders_6_io_output ? proc_5_io_next_header_48 : _GEN_4023; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4088 = 3'h5 == encoders_6_io_output ? proc_5_io_next_header_49 : _GEN_4024; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4089 = 3'h5 == encoders_6_io_output ? proc_5_io_next_header_50 : _GEN_4025; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4090 = 3'h5 == encoders_6_io_output ? proc_5_io_next_header_51 : _GEN_4026; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4091 = 3'h5 == encoders_6_io_output ? proc_5_io_next_header_52 : _GEN_4027; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4092 = 3'h5 == encoders_6_io_output ? proc_5_io_next_header_53 : _GEN_4028; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4093 = 3'h5 == encoders_6_io_output ? proc_5_io_next_header_54 : _GEN_4029; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4094 = 3'h5 == encoders_6_io_output ? proc_5_io_next_header_55 : _GEN_4030; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4095 = 3'h5 == encoders_6_io_output ? proc_5_io_next_header_56 : _GEN_4031; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4096 = 3'h5 == encoders_6_io_output ? proc_5_io_next_header_57 : _GEN_4032; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4097 = 3'h5 == encoders_6_io_output ? proc_5_io_next_header_58 : _GEN_4033; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4098 = 3'h5 == encoders_6_io_output ? proc_5_io_next_header_59 : _GEN_4034; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4099 = 3'h5 == encoders_6_io_output ? proc_5_io_next_header_60 : _GEN_4035; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4100 = 3'h5 == encoders_6_io_output ? proc_5_io_next_header_61 : _GEN_4036; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4101 = 3'h5 == encoders_6_io_output ? proc_5_io_next_header_62 : _GEN_4037; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4102 = 3'h5 == encoders_6_io_output ? proc_5_io_next_header_63 : _GEN_4038; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4103 = 3'h6 == encoders_6_io_output ? proc_6_io_next_header_0 : _GEN_4039; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4104 = 3'h6 == encoders_6_io_output ? proc_6_io_next_header_1 : _GEN_4040; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4105 = 3'h6 == encoders_6_io_output ? proc_6_io_next_header_2 : _GEN_4041; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4106 = 3'h6 == encoders_6_io_output ? proc_6_io_next_header_3 : _GEN_4042; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4107 = 3'h6 == encoders_6_io_output ? proc_6_io_next_header_4 : _GEN_4043; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4108 = 3'h6 == encoders_6_io_output ? proc_6_io_next_header_5 : _GEN_4044; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4109 = 3'h6 == encoders_6_io_output ? proc_6_io_next_header_6 : _GEN_4045; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4110 = 3'h6 == encoders_6_io_output ? proc_6_io_next_header_7 : _GEN_4046; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4111 = 3'h6 == encoders_6_io_output ? proc_6_io_next_header_8 : _GEN_4047; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4112 = 3'h6 == encoders_6_io_output ? proc_6_io_next_header_9 : _GEN_4048; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4113 = 3'h6 == encoders_6_io_output ? proc_6_io_next_header_10 : _GEN_4049; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4114 = 3'h6 == encoders_6_io_output ? proc_6_io_next_header_11 : _GEN_4050; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4115 = 3'h6 == encoders_6_io_output ? proc_6_io_next_header_12 : _GEN_4051; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4116 = 3'h6 == encoders_6_io_output ? proc_6_io_next_header_13 : _GEN_4052; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4117 = 3'h6 == encoders_6_io_output ? proc_6_io_next_header_14 : _GEN_4053; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4118 = 3'h6 == encoders_6_io_output ? proc_6_io_next_header_15 : _GEN_4054; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4119 = 3'h6 == encoders_6_io_output ? proc_6_io_next_header_16 : _GEN_4055; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4120 = 3'h6 == encoders_6_io_output ? proc_6_io_next_header_17 : _GEN_4056; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4121 = 3'h6 == encoders_6_io_output ? proc_6_io_next_header_18 : _GEN_4057; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4122 = 3'h6 == encoders_6_io_output ? proc_6_io_next_header_19 : _GEN_4058; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4123 = 3'h6 == encoders_6_io_output ? proc_6_io_next_header_20 : _GEN_4059; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4124 = 3'h6 == encoders_6_io_output ? proc_6_io_next_header_21 : _GEN_4060; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4125 = 3'h6 == encoders_6_io_output ? proc_6_io_next_header_22 : _GEN_4061; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4126 = 3'h6 == encoders_6_io_output ? proc_6_io_next_header_23 : _GEN_4062; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4127 = 3'h6 == encoders_6_io_output ? proc_6_io_next_header_24 : _GEN_4063; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4128 = 3'h6 == encoders_6_io_output ? proc_6_io_next_header_25 : _GEN_4064; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4129 = 3'h6 == encoders_6_io_output ? proc_6_io_next_header_26 : _GEN_4065; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4130 = 3'h6 == encoders_6_io_output ? proc_6_io_next_header_27 : _GEN_4066; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4131 = 3'h6 == encoders_6_io_output ? proc_6_io_next_header_28 : _GEN_4067; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4132 = 3'h6 == encoders_6_io_output ? proc_6_io_next_header_29 : _GEN_4068; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4133 = 3'h6 == encoders_6_io_output ? proc_6_io_next_header_30 : _GEN_4069; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4134 = 3'h6 == encoders_6_io_output ? proc_6_io_next_header_31 : _GEN_4070; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4135 = 3'h6 == encoders_6_io_output ? proc_6_io_next_header_32 : _GEN_4071; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4136 = 3'h6 == encoders_6_io_output ? proc_6_io_next_header_33 : _GEN_4072; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4137 = 3'h6 == encoders_6_io_output ? proc_6_io_next_header_34 : _GEN_4073; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4138 = 3'h6 == encoders_6_io_output ? proc_6_io_next_header_35 : _GEN_4074; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4139 = 3'h6 == encoders_6_io_output ? proc_6_io_next_header_36 : _GEN_4075; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4140 = 3'h6 == encoders_6_io_output ? proc_6_io_next_header_37 : _GEN_4076; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4141 = 3'h6 == encoders_6_io_output ? proc_6_io_next_header_38 : _GEN_4077; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4142 = 3'h6 == encoders_6_io_output ? proc_6_io_next_header_39 : _GEN_4078; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4143 = 3'h6 == encoders_6_io_output ? proc_6_io_next_header_40 : _GEN_4079; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4144 = 3'h6 == encoders_6_io_output ? proc_6_io_next_header_41 : _GEN_4080; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4145 = 3'h6 == encoders_6_io_output ? proc_6_io_next_header_42 : _GEN_4081; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4146 = 3'h6 == encoders_6_io_output ? proc_6_io_next_header_43 : _GEN_4082; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4147 = 3'h6 == encoders_6_io_output ? proc_6_io_next_header_44 : _GEN_4083; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4148 = 3'h6 == encoders_6_io_output ? proc_6_io_next_header_45 : _GEN_4084; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4149 = 3'h6 == encoders_6_io_output ? proc_6_io_next_header_46 : _GEN_4085; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4150 = 3'h6 == encoders_6_io_output ? proc_6_io_next_header_47 : _GEN_4086; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4151 = 3'h6 == encoders_6_io_output ? proc_6_io_next_header_48 : _GEN_4087; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4152 = 3'h6 == encoders_6_io_output ? proc_6_io_next_header_49 : _GEN_4088; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4153 = 3'h6 == encoders_6_io_output ? proc_6_io_next_header_50 : _GEN_4089; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4154 = 3'h6 == encoders_6_io_output ? proc_6_io_next_header_51 : _GEN_4090; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4155 = 3'h6 == encoders_6_io_output ? proc_6_io_next_header_52 : _GEN_4091; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4156 = 3'h6 == encoders_6_io_output ? proc_6_io_next_header_53 : _GEN_4092; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4157 = 3'h6 == encoders_6_io_output ? proc_6_io_next_header_54 : _GEN_4093; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4158 = 3'h6 == encoders_6_io_output ? proc_6_io_next_header_55 : _GEN_4094; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4159 = 3'h6 == encoders_6_io_output ? proc_6_io_next_header_56 : _GEN_4095; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4160 = 3'h6 == encoders_6_io_output ? proc_6_io_next_header_57 : _GEN_4096; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4161 = 3'h6 == encoders_6_io_output ? proc_6_io_next_header_58 : _GEN_4097; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4162 = 3'h6 == encoders_6_io_output ? proc_6_io_next_header_59 : _GEN_4098; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4163 = 3'h6 == encoders_6_io_output ? proc_6_io_next_header_60 : _GEN_4099; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4164 = 3'h6 == encoders_6_io_output ? proc_6_io_next_header_61 : _GEN_4100; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4165 = 3'h6 == encoders_6_io_output ? proc_6_io_next_header_62 : _GEN_4101; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4166 = 3'h6 == encoders_6_io_output ? proc_6_io_next_header_63 : _GEN_4102; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4167 = 3'h7 == encoders_6_io_output ? proc_7_io_next_header_0 : _GEN_4103; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4168 = 3'h7 == encoders_6_io_output ? proc_7_io_next_header_1 : _GEN_4104; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4169 = 3'h7 == encoders_6_io_output ? proc_7_io_next_header_2 : _GEN_4105; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4170 = 3'h7 == encoders_6_io_output ? proc_7_io_next_header_3 : _GEN_4106; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4171 = 3'h7 == encoders_6_io_output ? proc_7_io_next_header_4 : _GEN_4107; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4172 = 3'h7 == encoders_6_io_output ? proc_7_io_next_header_5 : _GEN_4108; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4173 = 3'h7 == encoders_6_io_output ? proc_7_io_next_header_6 : _GEN_4109; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4174 = 3'h7 == encoders_6_io_output ? proc_7_io_next_header_7 : _GEN_4110; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4175 = 3'h7 == encoders_6_io_output ? proc_7_io_next_header_8 : _GEN_4111; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4176 = 3'h7 == encoders_6_io_output ? proc_7_io_next_header_9 : _GEN_4112; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4177 = 3'h7 == encoders_6_io_output ? proc_7_io_next_header_10 : _GEN_4113; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4178 = 3'h7 == encoders_6_io_output ? proc_7_io_next_header_11 : _GEN_4114; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4179 = 3'h7 == encoders_6_io_output ? proc_7_io_next_header_12 : _GEN_4115; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4180 = 3'h7 == encoders_6_io_output ? proc_7_io_next_header_13 : _GEN_4116; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4181 = 3'h7 == encoders_6_io_output ? proc_7_io_next_header_14 : _GEN_4117; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4182 = 3'h7 == encoders_6_io_output ? proc_7_io_next_header_15 : _GEN_4118; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4183 = 3'h7 == encoders_6_io_output ? proc_7_io_next_header_16 : _GEN_4119; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4184 = 3'h7 == encoders_6_io_output ? proc_7_io_next_header_17 : _GEN_4120; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4185 = 3'h7 == encoders_6_io_output ? proc_7_io_next_header_18 : _GEN_4121; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4186 = 3'h7 == encoders_6_io_output ? proc_7_io_next_header_19 : _GEN_4122; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4187 = 3'h7 == encoders_6_io_output ? proc_7_io_next_header_20 : _GEN_4123; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4188 = 3'h7 == encoders_6_io_output ? proc_7_io_next_header_21 : _GEN_4124; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4189 = 3'h7 == encoders_6_io_output ? proc_7_io_next_header_22 : _GEN_4125; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4190 = 3'h7 == encoders_6_io_output ? proc_7_io_next_header_23 : _GEN_4126; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4191 = 3'h7 == encoders_6_io_output ? proc_7_io_next_header_24 : _GEN_4127; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4192 = 3'h7 == encoders_6_io_output ? proc_7_io_next_header_25 : _GEN_4128; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4193 = 3'h7 == encoders_6_io_output ? proc_7_io_next_header_26 : _GEN_4129; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4194 = 3'h7 == encoders_6_io_output ? proc_7_io_next_header_27 : _GEN_4130; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4195 = 3'h7 == encoders_6_io_output ? proc_7_io_next_header_28 : _GEN_4131; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4196 = 3'h7 == encoders_6_io_output ? proc_7_io_next_header_29 : _GEN_4132; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4197 = 3'h7 == encoders_6_io_output ? proc_7_io_next_header_30 : _GEN_4133; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4198 = 3'h7 == encoders_6_io_output ? proc_7_io_next_header_31 : _GEN_4134; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4199 = 3'h7 == encoders_6_io_output ? proc_7_io_next_header_32 : _GEN_4135; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4200 = 3'h7 == encoders_6_io_output ? proc_7_io_next_header_33 : _GEN_4136; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4201 = 3'h7 == encoders_6_io_output ? proc_7_io_next_header_34 : _GEN_4137; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4202 = 3'h7 == encoders_6_io_output ? proc_7_io_next_header_35 : _GEN_4138; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4203 = 3'h7 == encoders_6_io_output ? proc_7_io_next_header_36 : _GEN_4139; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4204 = 3'h7 == encoders_6_io_output ? proc_7_io_next_header_37 : _GEN_4140; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4205 = 3'h7 == encoders_6_io_output ? proc_7_io_next_header_38 : _GEN_4141; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4206 = 3'h7 == encoders_6_io_output ? proc_7_io_next_header_39 : _GEN_4142; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4207 = 3'h7 == encoders_6_io_output ? proc_7_io_next_header_40 : _GEN_4143; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4208 = 3'h7 == encoders_6_io_output ? proc_7_io_next_header_41 : _GEN_4144; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4209 = 3'h7 == encoders_6_io_output ? proc_7_io_next_header_42 : _GEN_4145; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4210 = 3'h7 == encoders_6_io_output ? proc_7_io_next_header_43 : _GEN_4146; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4211 = 3'h7 == encoders_6_io_output ? proc_7_io_next_header_44 : _GEN_4147; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4212 = 3'h7 == encoders_6_io_output ? proc_7_io_next_header_45 : _GEN_4148; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4213 = 3'h7 == encoders_6_io_output ? proc_7_io_next_header_46 : _GEN_4149; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4214 = 3'h7 == encoders_6_io_output ? proc_7_io_next_header_47 : _GEN_4150; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4215 = 3'h7 == encoders_6_io_output ? proc_7_io_next_header_48 : _GEN_4151; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4216 = 3'h7 == encoders_6_io_output ? proc_7_io_next_header_49 : _GEN_4152; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4217 = 3'h7 == encoders_6_io_output ? proc_7_io_next_header_50 : _GEN_4153; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4218 = 3'h7 == encoders_6_io_output ? proc_7_io_next_header_51 : _GEN_4154; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4219 = 3'h7 == encoders_6_io_output ? proc_7_io_next_header_52 : _GEN_4155; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4220 = 3'h7 == encoders_6_io_output ? proc_7_io_next_header_53 : _GEN_4156; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4221 = 3'h7 == encoders_6_io_output ? proc_7_io_next_header_54 : _GEN_4157; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4222 = 3'h7 == encoders_6_io_output ? proc_7_io_next_header_55 : _GEN_4158; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4223 = 3'h7 == encoders_6_io_output ? proc_7_io_next_header_56 : _GEN_4159; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4224 = 3'h7 == encoders_6_io_output ? proc_7_io_next_header_57 : _GEN_4160; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4225 = 3'h7 == encoders_6_io_output ? proc_7_io_next_header_58 : _GEN_4161; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4226 = 3'h7 == encoders_6_io_output ? proc_7_io_next_header_59 : _GEN_4162; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4227 = 3'h7 == encoders_6_io_output ? proc_7_io_next_header_60 : _GEN_4163; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4228 = 3'h7 == encoders_6_io_output ? proc_7_io_next_header_61 : _GEN_4164; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4229 = 3'h7 == encoders_6_io_output ? proc_7_io_next_header_62 : _GEN_4165; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4230 = 3'h7 == encoders_6_io_output ? proc_7_io_next_header_63 : _GEN_4166; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4296 = 3'h0 == encoders_7_io_output ? proc_0_io_next_header_0 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_4297 = 3'h0 == encoders_7_io_output ? proc_0_io_next_header_1 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_4298 = 3'h0 == encoders_7_io_output ? proc_0_io_next_header_2 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_4299 = 3'h0 == encoders_7_io_output ? proc_0_io_next_header_3 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_4300 = 3'h0 == encoders_7_io_output ? proc_0_io_next_header_4 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_4301 = 3'h0 == encoders_7_io_output ? proc_0_io_next_header_5 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_4302 = 3'h0 == encoders_7_io_output ? proc_0_io_next_header_6 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_4303 = 3'h0 == encoders_7_io_output ? proc_0_io_next_header_7 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_4304 = 3'h0 == encoders_7_io_output ? proc_0_io_next_header_8 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_4305 = 3'h0 == encoders_7_io_output ? proc_0_io_next_header_9 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_4306 = 3'h0 == encoders_7_io_output ? proc_0_io_next_header_10 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_4307 = 3'h0 == encoders_7_io_output ? proc_0_io_next_header_11 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_4308 = 3'h0 == encoders_7_io_output ? proc_0_io_next_header_12 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_4309 = 3'h0 == encoders_7_io_output ? proc_0_io_next_header_13 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_4310 = 3'h0 == encoders_7_io_output ? proc_0_io_next_header_14 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_4311 = 3'h0 == encoders_7_io_output ? proc_0_io_next_header_15 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_4312 = 3'h0 == encoders_7_io_output ? proc_0_io_next_header_16 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_4313 = 3'h0 == encoders_7_io_output ? proc_0_io_next_header_17 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_4314 = 3'h0 == encoders_7_io_output ? proc_0_io_next_header_18 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_4315 = 3'h0 == encoders_7_io_output ? proc_0_io_next_header_19 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_4316 = 3'h0 == encoders_7_io_output ? proc_0_io_next_header_20 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_4317 = 3'h0 == encoders_7_io_output ? proc_0_io_next_header_21 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_4318 = 3'h0 == encoders_7_io_output ? proc_0_io_next_header_22 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_4319 = 3'h0 == encoders_7_io_output ? proc_0_io_next_header_23 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_4320 = 3'h0 == encoders_7_io_output ? proc_0_io_next_header_24 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_4321 = 3'h0 == encoders_7_io_output ? proc_0_io_next_header_25 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_4322 = 3'h0 == encoders_7_io_output ? proc_0_io_next_header_26 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_4323 = 3'h0 == encoders_7_io_output ? proc_0_io_next_header_27 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_4324 = 3'h0 == encoders_7_io_output ? proc_0_io_next_header_28 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_4325 = 3'h0 == encoders_7_io_output ? proc_0_io_next_header_29 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_4326 = 3'h0 == encoders_7_io_output ? proc_0_io_next_header_30 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_4327 = 3'h0 == encoders_7_io_output ? proc_0_io_next_header_31 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_4328 = 3'h0 == encoders_7_io_output ? proc_0_io_next_header_32 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_4329 = 3'h0 == encoders_7_io_output ? proc_0_io_next_header_33 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_4330 = 3'h0 == encoders_7_io_output ? proc_0_io_next_header_34 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_4331 = 3'h0 == encoders_7_io_output ? proc_0_io_next_header_35 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_4332 = 3'h0 == encoders_7_io_output ? proc_0_io_next_header_36 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_4333 = 3'h0 == encoders_7_io_output ? proc_0_io_next_header_37 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_4334 = 3'h0 == encoders_7_io_output ? proc_0_io_next_header_38 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_4335 = 3'h0 == encoders_7_io_output ? proc_0_io_next_header_39 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_4336 = 3'h0 == encoders_7_io_output ? proc_0_io_next_header_40 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_4337 = 3'h0 == encoders_7_io_output ? proc_0_io_next_header_41 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_4338 = 3'h0 == encoders_7_io_output ? proc_0_io_next_header_42 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_4339 = 3'h0 == encoders_7_io_output ? proc_0_io_next_header_43 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_4340 = 3'h0 == encoders_7_io_output ? proc_0_io_next_header_44 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_4341 = 3'h0 == encoders_7_io_output ? proc_0_io_next_header_45 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_4342 = 3'h0 == encoders_7_io_output ? proc_0_io_next_header_46 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_4343 = 3'h0 == encoders_7_io_output ? proc_0_io_next_header_47 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_4344 = 3'h0 == encoders_7_io_output ? proc_0_io_next_header_48 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_4345 = 3'h0 == encoders_7_io_output ? proc_0_io_next_header_49 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_4346 = 3'h0 == encoders_7_io_output ? proc_0_io_next_header_50 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_4347 = 3'h0 == encoders_7_io_output ? proc_0_io_next_header_51 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_4348 = 3'h0 == encoders_7_io_output ? proc_0_io_next_header_52 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_4349 = 3'h0 == encoders_7_io_output ? proc_0_io_next_header_53 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_4350 = 3'h0 == encoders_7_io_output ? proc_0_io_next_header_54 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_4351 = 3'h0 == encoders_7_io_output ? proc_0_io_next_header_55 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_4352 = 3'h0 == encoders_7_io_output ? proc_0_io_next_header_56 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_4353 = 3'h0 == encoders_7_io_output ? proc_0_io_next_header_57 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_4354 = 3'h0 == encoders_7_io_output ? proc_0_io_next_header_58 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_4355 = 3'h0 == encoders_7_io_output ? proc_0_io_next_header_59 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_4356 = 3'h0 == encoders_7_io_output ? proc_0_io_next_header_60 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_4357 = 3'h0 == encoders_7_io_output ? proc_0_io_next_header_61 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_4358 = 3'h0 == encoders_7_io_output ? proc_0_io_next_header_62 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_4359 = 3'h0 == encoders_7_io_output ? proc_0_io_next_header_63 : 8'h0; // @[controller.scala 94:46 controller.scala 95:46 controller.scala 42:41]
  wire [7:0] _GEN_4360 = 3'h1 == encoders_7_io_output ? proc_1_io_next_header_0 : _GEN_4296; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4361 = 3'h1 == encoders_7_io_output ? proc_1_io_next_header_1 : _GEN_4297; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4362 = 3'h1 == encoders_7_io_output ? proc_1_io_next_header_2 : _GEN_4298; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4363 = 3'h1 == encoders_7_io_output ? proc_1_io_next_header_3 : _GEN_4299; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4364 = 3'h1 == encoders_7_io_output ? proc_1_io_next_header_4 : _GEN_4300; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4365 = 3'h1 == encoders_7_io_output ? proc_1_io_next_header_5 : _GEN_4301; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4366 = 3'h1 == encoders_7_io_output ? proc_1_io_next_header_6 : _GEN_4302; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4367 = 3'h1 == encoders_7_io_output ? proc_1_io_next_header_7 : _GEN_4303; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4368 = 3'h1 == encoders_7_io_output ? proc_1_io_next_header_8 : _GEN_4304; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4369 = 3'h1 == encoders_7_io_output ? proc_1_io_next_header_9 : _GEN_4305; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4370 = 3'h1 == encoders_7_io_output ? proc_1_io_next_header_10 : _GEN_4306; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4371 = 3'h1 == encoders_7_io_output ? proc_1_io_next_header_11 : _GEN_4307; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4372 = 3'h1 == encoders_7_io_output ? proc_1_io_next_header_12 : _GEN_4308; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4373 = 3'h1 == encoders_7_io_output ? proc_1_io_next_header_13 : _GEN_4309; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4374 = 3'h1 == encoders_7_io_output ? proc_1_io_next_header_14 : _GEN_4310; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4375 = 3'h1 == encoders_7_io_output ? proc_1_io_next_header_15 : _GEN_4311; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4376 = 3'h1 == encoders_7_io_output ? proc_1_io_next_header_16 : _GEN_4312; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4377 = 3'h1 == encoders_7_io_output ? proc_1_io_next_header_17 : _GEN_4313; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4378 = 3'h1 == encoders_7_io_output ? proc_1_io_next_header_18 : _GEN_4314; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4379 = 3'h1 == encoders_7_io_output ? proc_1_io_next_header_19 : _GEN_4315; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4380 = 3'h1 == encoders_7_io_output ? proc_1_io_next_header_20 : _GEN_4316; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4381 = 3'h1 == encoders_7_io_output ? proc_1_io_next_header_21 : _GEN_4317; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4382 = 3'h1 == encoders_7_io_output ? proc_1_io_next_header_22 : _GEN_4318; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4383 = 3'h1 == encoders_7_io_output ? proc_1_io_next_header_23 : _GEN_4319; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4384 = 3'h1 == encoders_7_io_output ? proc_1_io_next_header_24 : _GEN_4320; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4385 = 3'h1 == encoders_7_io_output ? proc_1_io_next_header_25 : _GEN_4321; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4386 = 3'h1 == encoders_7_io_output ? proc_1_io_next_header_26 : _GEN_4322; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4387 = 3'h1 == encoders_7_io_output ? proc_1_io_next_header_27 : _GEN_4323; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4388 = 3'h1 == encoders_7_io_output ? proc_1_io_next_header_28 : _GEN_4324; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4389 = 3'h1 == encoders_7_io_output ? proc_1_io_next_header_29 : _GEN_4325; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4390 = 3'h1 == encoders_7_io_output ? proc_1_io_next_header_30 : _GEN_4326; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4391 = 3'h1 == encoders_7_io_output ? proc_1_io_next_header_31 : _GEN_4327; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4392 = 3'h1 == encoders_7_io_output ? proc_1_io_next_header_32 : _GEN_4328; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4393 = 3'h1 == encoders_7_io_output ? proc_1_io_next_header_33 : _GEN_4329; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4394 = 3'h1 == encoders_7_io_output ? proc_1_io_next_header_34 : _GEN_4330; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4395 = 3'h1 == encoders_7_io_output ? proc_1_io_next_header_35 : _GEN_4331; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4396 = 3'h1 == encoders_7_io_output ? proc_1_io_next_header_36 : _GEN_4332; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4397 = 3'h1 == encoders_7_io_output ? proc_1_io_next_header_37 : _GEN_4333; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4398 = 3'h1 == encoders_7_io_output ? proc_1_io_next_header_38 : _GEN_4334; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4399 = 3'h1 == encoders_7_io_output ? proc_1_io_next_header_39 : _GEN_4335; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4400 = 3'h1 == encoders_7_io_output ? proc_1_io_next_header_40 : _GEN_4336; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4401 = 3'h1 == encoders_7_io_output ? proc_1_io_next_header_41 : _GEN_4337; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4402 = 3'h1 == encoders_7_io_output ? proc_1_io_next_header_42 : _GEN_4338; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4403 = 3'h1 == encoders_7_io_output ? proc_1_io_next_header_43 : _GEN_4339; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4404 = 3'h1 == encoders_7_io_output ? proc_1_io_next_header_44 : _GEN_4340; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4405 = 3'h1 == encoders_7_io_output ? proc_1_io_next_header_45 : _GEN_4341; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4406 = 3'h1 == encoders_7_io_output ? proc_1_io_next_header_46 : _GEN_4342; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4407 = 3'h1 == encoders_7_io_output ? proc_1_io_next_header_47 : _GEN_4343; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4408 = 3'h1 == encoders_7_io_output ? proc_1_io_next_header_48 : _GEN_4344; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4409 = 3'h1 == encoders_7_io_output ? proc_1_io_next_header_49 : _GEN_4345; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4410 = 3'h1 == encoders_7_io_output ? proc_1_io_next_header_50 : _GEN_4346; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4411 = 3'h1 == encoders_7_io_output ? proc_1_io_next_header_51 : _GEN_4347; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4412 = 3'h1 == encoders_7_io_output ? proc_1_io_next_header_52 : _GEN_4348; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4413 = 3'h1 == encoders_7_io_output ? proc_1_io_next_header_53 : _GEN_4349; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4414 = 3'h1 == encoders_7_io_output ? proc_1_io_next_header_54 : _GEN_4350; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4415 = 3'h1 == encoders_7_io_output ? proc_1_io_next_header_55 : _GEN_4351; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4416 = 3'h1 == encoders_7_io_output ? proc_1_io_next_header_56 : _GEN_4352; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4417 = 3'h1 == encoders_7_io_output ? proc_1_io_next_header_57 : _GEN_4353; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4418 = 3'h1 == encoders_7_io_output ? proc_1_io_next_header_58 : _GEN_4354; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4419 = 3'h1 == encoders_7_io_output ? proc_1_io_next_header_59 : _GEN_4355; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4420 = 3'h1 == encoders_7_io_output ? proc_1_io_next_header_60 : _GEN_4356; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4421 = 3'h1 == encoders_7_io_output ? proc_1_io_next_header_61 : _GEN_4357; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4422 = 3'h1 == encoders_7_io_output ? proc_1_io_next_header_62 : _GEN_4358; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4423 = 3'h1 == encoders_7_io_output ? proc_1_io_next_header_63 : _GEN_4359; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4424 = 3'h2 == encoders_7_io_output ? proc_2_io_next_header_0 : _GEN_4360; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4425 = 3'h2 == encoders_7_io_output ? proc_2_io_next_header_1 : _GEN_4361; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4426 = 3'h2 == encoders_7_io_output ? proc_2_io_next_header_2 : _GEN_4362; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4427 = 3'h2 == encoders_7_io_output ? proc_2_io_next_header_3 : _GEN_4363; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4428 = 3'h2 == encoders_7_io_output ? proc_2_io_next_header_4 : _GEN_4364; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4429 = 3'h2 == encoders_7_io_output ? proc_2_io_next_header_5 : _GEN_4365; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4430 = 3'h2 == encoders_7_io_output ? proc_2_io_next_header_6 : _GEN_4366; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4431 = 3'h2 == encoders_7_io_output ? proc_2_io_next_header_7 : _GEN_4367; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4432 = 3'h2 == encoders_7_io_output ? proc_2_io_next_header_8 : _GEN_4368; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4433 = 3'h2 == encoders_7_io_output ? proc_2_io_next_header_9 : _GEN_4369; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4434 = 3'h2 == encoders_7_io_output ? proc_2_io_next_header_10 : _GEN_4370; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4435 = 3'h2 == encoders_7_io_output ? proc_2_io_next_header_11 : _GEN_4371; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4436 = 3'h2 == encoders_7_io_output ? proc_2_io_next_header_12 : _GEN_4372; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4437 = 3'h2 == encoders_7_io_output ? proc_2_io_next_header_13 : _GEN_4373; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4438 = 3'h2 == encoders_7_io_output ? proc_2_io_next_header_14 : _GEN_4374; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4439 = 3'h2 == encoders_7_io_output ? proc_2_io_next_header_15 : _GEN_4375; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4440 = 3'h2 == encoders_7_io_output ? proc_2_io_next_header_16 : _GEN_4376; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4441 = 3'h2 == encoders_7_io_output ? proc_2_io_next_header_17 : _GEN_4377; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4442 = 3'h2 == encoders_7_io_output ? proc_2_io_next_header_18 : _GEN_4378; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4443 = 3'h2 == encoders_7_io_output ? proc_2_io_next_header_19 : _GEN_4379; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4444 = 3'h2 == encoders_7_io_output ? proc_2_io_next_header_20 : _GEN_4380; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4445 = 3'h2 == encoders_7_io_output ? proc_2_io_next_header_21 : _GEN_4381; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4446 = 3'h2 == encoders_7_io_output ? proc_2_io_next_header_22 : _GEN_4382; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4447 = 3'h2 == encoders_7_io_output ? proc_2_io_next_header_23 : _GEN_4383; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4448 = 3'h2 == encoders_7_io_output ? proc_2_io_next_header_24 : _GEN_4384; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4449 = 3'h2 == encoders_7_io_output ? proc_2_io_next_header_25 : _GEN_4385; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4450 = 3'h2 == encoders_7_io_output ? proc_2_io_next_header_26 : _GEN_4386; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4451 = 3'h2 == encoders_7_io_output ? proc_2_io_next_header_27 : _GEN_4387; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4452 = 3'h2 == encoders_7_io_output ? proc_2_io_next_header_28 : _GEN_4388; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4453 = 3'h2 == encoders_7_io_output ? proc_2_io_next_header_29 : _GEN_4389; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4454 = 3'h2 == encoders_7_io_output ? proc_2_io_next_header_30 : _GEN_4390; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4455 = 3'h2 == encoders_7_io_output ? proc_2_io_next_header_31 : _GEN_4391; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4456 = 3'h2 == encoders_7_io_output ? proc_2_io_next_header_32 : _GEN_4392; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4457 = 3'h2 == encoders_7_io_output ? proc_2_io_next_header_33 : _GEN_4393; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4458 = 3'h2 == encoders_7_io_output ? proc_2_io_next_header_34 : _GEN_4394; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4459 = 3'h2 == encoders_7_io_output ? proc_2_io_next_header_35 : _GEN_4395; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4460 = 3'h2 == encoders_7_io_output ? proc_2_io_next_header_36 : _GEN_4396; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4461 = 3'h2 == encoders_7_io_output ? proc_2_io_next_header_37 : _GEN_4397; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4462 = 3'h2 == encoders_7_io_output ? proc_2_io_next_header_38 : _GEN_4398; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4463 = 3'h2 == encoders_7_io_output ? proc_2_io_next_header_39 : _GEN_4399; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4464 = 3'h2 == encoders_7_io_output ? proc_2_io_next_header_40 : _GEN_4400; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4465 = 3'h2 == encoders_7_io_output ? proc_2_io_next_header_41 : _GEN_4401; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4466 = 3'h2 == encoders_7_io_output ? proc_2_io_next_header_42 : _GEN_4402; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4467 = 3'h2 == encoders_7_io_output ? proc_2_io_next_header_43 : _GEN_4403; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4468 = 3'h2 == encoders_7_io_output ? proc_2_io_next_header_44 : _GEN_4404; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4469 = 3'h2 == encoders_7_io_output ? proc_2_io_next_header_45 : _GEN_4405; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4470 = 3'h2 == encoders_7_io_output ? proc_2_io_next_header_46 : _GEN_4406; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4471 = 3'h2 == encoders_7_io_output ? proc_2_io_next_header_47 : _GEN_4407; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4472 = 3'h2 == encoders_7_io_output ? proc_2_io_next_header_48 : _GEN_4408; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4473 = 3'h2 == encoders_7_io_output ? proc_2_io_next_header_49 : _GEN_4409; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4474 = 3'h2 == encoders_7_io_output ? proc_2_io_next_header_50 : _GEN_4410; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4475 = 3'h2 == encoders_7_io_output ? proc_2_io_next_header_51 : _GEN_4411; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4476 = 3'h2 == encoders_7_io_output ? proc_2_io_next_header_52 : _GEN_4412; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4477 = 3'h2 == encoders_7_io_output ? proc_2_io_next_header_53 : _GEN_4413; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4478 = 3'h2 == encoders_7_io_output ? proc_2_io_next_header_54 : _GEN_4414; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4479 = 3'h2 == encoders_7_io_output ? proc_2_io_next_header_55 : _GEN_4415; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4480 = 3'h2 == encoders_7_io_output ? proc_2_io_next_header_56 : _GEN_4416; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4481 = 3'h2 == encoders_7_io_output ? proc_2_io_next_header_57 : _GEN_4417; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4482 = 3'h2 == encoders_7_io_output ? proc_2_io_next_header_58 : _GEN_4418; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4483 = 3'h2 == encoders_7_io_output ? proc_2_io_next_header_59 : _GEN_4419; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4484 = 3'h2 == encoders_7_io_output ? proc_2_io_next_header_60 : _GEN_4420; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4485 = 3'h2 == encoders_7_io_output ? proc_2_io_next_header_61 : _GEN_4421; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4486 = 3'h2 == encoders_7_io_output ? proc_2_io_next_header_62 : _GEN_4422; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4487 = 3'h2 == encoders_7_io_output ? proc_2_io_next_header_63 : _GEN_4423; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4488 = 3'h3 == encoders_7_io_output ? proc_3_io_next_header_0 : _GEN_4424; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4489 = 3'h3 == encoders_7_io_output ? proc_3_io_next_header_1 : _GEN_4425; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4490 = 3'h3 == encoders_7_io_output ? proc_3_io_next_header_2 : _GEN_4426; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4491 = 3'h3 == encoders_7_io_output ? proc_3_io_next_header_3 : _GEN_4427; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4492 = 3'h3 == encoders_7_io_output ? proc_3_io_next_header_4 : _GEN_4428; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4493 = 3'h3 == encoders_7_io_output ? proc_3_io_next_header_5 : _GEN_4429; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4494 = 3'h3 == encoders_7_io_output ? proc_3_io_next_header_6 : _GEN_4430; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4495 = 3'h3 == encoders_7_io_output ? proc_3_io_next_header_7 : _GEN_4431; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4496 = 3'h3 == encoders_7_io_output ? proc_3_io_next_header_8 : _GEN_4432; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4497 = 3'h3 == encoders_7_io_output ? proc_3_io_next_header_9 : _GEN_4433; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4498 = 3'h3 == encoders_7_io_output ? proc_3_io_next_header_10 : _GEN_4434; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4499 = 3'h3 == encoders_7_io_output ? proc_3_io_next_header_11 : _GEN_4435; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4500 = 3'h3 == encoders_7_io_output ? proc_3_io_next_header_12 : _GEN_4436; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4501 = 3'h3 == encoders_7_io_output ? proc_3_io_next_header_13 : _GEN_4437; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4502 = 3'h3 == encoders_7_io_output ? proc_3_io_next_header_14 : _GEN_4438; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4503 = 3'h3 == encoders_7_io_output ? proc_3_io_next_header_15 : _GEN_4439; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4504 = 3'h3 == encoders_7_io_output ? proc_3_io_next_header_16 : _GEN_4440; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4505 = 3'h3 == encoders_7_io_output ? proc_3_io_next_header_17 : _GEN_4441; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4506 = 3'h3 == encoders_7_io_output ? proc_3_io_next_header_18 : _GEN_4442; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4507 = 3'h3 == encoders_7_io_output ? proc_3_io_next_header_19 : _GEN_4443; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4508 = 3'h3 == encoders_7_io_output ? proc_3_io_next_header_20 : _GEN_4444; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4509 = 3'h3 == encoders_7_io_output ? proc_3_io_next_header_21 : _GEN_4445; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4510 = 3'h3 == encoders_7_io_output ? proc_3_io_next_header_22 : _GEN_4446; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4511 = 3'h3 == encoders_7_io_output ? proc_3_io_next_header_23 : _GEN_4447; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4512 = 3'h3 == encoders_7_io_output ? proc_3_io_next_header_24 : _GEN_4448; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4513 = 3'h3 == encoders_7_io_output ? proc_3_io_next_header_25 : _GEN_4449; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4514 = 3'h3 == encoders_7_io_output ? proc_3_io_next_header_26 : _GEN_4450; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4515 = 3'h3 == encoders_7_io_output ? proc_3_io_next_header_27 : _GEN_4451; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4516 = 3'h3 == encoders_7_io_output ? proc_3_io_next_header_28 : _GEN_4452; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4517 = 3'h3 == encoders_7_io_output ? proc_3_io_next_header_29 : _GEN_4453; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4518 = 3'h3 == encoders_7_io_output ? proc_3_io_next_header_30 : _GEN_4454; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4519 = 3'h3 == encoders_7_io_output ? proc_3_io_next_header_31 : _GEN_4455; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4520 = 3'h3 == encoders_7_io_output ? proc_3_io_next_header_32 : _GEN_4456; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4521 = 3'h3 == encoders_7_io_output ? proc_3_io_next_header_33 : _GEN_4457; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4522 = 3'h3 == encoders_7_io_output ? proc_3_io_next_header_34 : _GEN_4458; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4523 = 3'h3 == encoders_7_io_output ? proc_3_io_next_header_35 : _GEN_4459; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4524 = 3'h3 == encoders_7_io_output ? proc_3_io_next_header_36 : _GEN_4460; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4525 = 3'h3 == encoders_7_io_output ? proc_3_io_next_header_37 : _GEN_4461; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4526 = 3'h3 == encoders_7_io_output ? proc_3_io_next_header_38 : _GEN_4462; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4527 = 3'h3 == encoders_7_io_output ? proc_3_io_next_header_39 : _GEN_4463; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4528 = 3'h3 == encoders_7_io_output ? proc_3_io_next_header_40 : _GEN_4464; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4529 = 3'h3 == encoders_7_io_output ? proc_3_io_next_header_41 : _GEN_4465; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4530 = 3'h3 == encoders_7_io_output ? proc_3_io_next_header_42 : _GEN_4466; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4531 = 3'h3 == encoders_7_io_output ? proc_3_io_next_header_43 : _GEN_4467; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4532 = 3'h3 == encoders_7_io_output ? proc_3_io_next_header_44 : _GEN_4468; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4533 = 3'h3 == encoders_7_io_output ? proc_3_io_next_header_45 : _GEN_4469; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4534 = 3'h3 == encoders_7_io_output ? proc_3_io_next_header_46 : _GEN_4470; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4535 = 3'h3 == encoders_7_io_output ? proc_3_io_next_header_47 : _GEN_4471; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4536 = 3'h3 == encoders_7_io_output ? proc_3_io_next_header_48 : _GEN_4472; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4537 = 3'h3 == encoders_7_io_output ? proc_3_io_next_header_49 : _GEN_4473; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4538 = 3'h3 == encoders_7_io_output ? proc_3_io_next_header_50 : _GEN_4474; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4539 = 3'h3 == encoders_7_io_output ? proc_3_io_next_header_51 : _GEN_4475; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4540 = 3'h3 == encoders_7_io_output ? proc_3_io_next_header_52 : _GEN_4476; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4541 = 3'h3 == encoders_7_io_output ? proc_3_io_next_header_53 : _GEN_4477; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4542 = 3'h3 == encoders_7_io_output ? proc_3_io_next_header_54 : _GEN_4478; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4543 = 3'h3 == encoders_7_io_output ? proc_3_io_next_header_55 : _GEN_4479; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4544 = 3'h3 == encoders_7_io_output ? proc_3_io_next_header_56 : _GEN_4480; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4545 = 3'h3 == encoders_7_io_output ? proc_3_io_next_header_57 : _GEN_4481; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4546 = 3'h3 == encoders_7_io_output ? proc_3_io_next_header_58 : _GEN_4482; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4547 = 3'h3 == encoders_7_io_output ? proc_3_io_next_header_59 : _GEN_4483; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4548 = 3'h3 == encoders_7_io_output ? proc_3_io_next_header_60 : _GEN_4484; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4549 = 3'h3 == encoders_7_io_output ? proc_3_io_next_header_61 : _GEN_4485; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4550 = 3'h3 == encoders_7_io_output ? proc_3_io_next_header_62 : _GEN_4486; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4551 = 3'h3 == encoders_7_io_output ? proc_3_io_next_header_63 : _GEN_4487; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4552 = 3'h4 == encoders_7_io_output ? proc_4_io_next_header_0 : _GEN_4488; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4553 = 3'h4 == encoders_7_io_output ? proc_4_io_next_header_1 : _GEN_4489; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4554 = 3'h4 == encoders_7_io_output ? proc_4_io_next_header_2 : _GEN_4490; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4555 = 3'h4 == encoders_7_io_output ? proc_4_io_next_header_3 : _GEN_4491; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4556 = 3'h4 == encoders_7_io_output ? proc_4_io_next_header_4 : _GEN_4492; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4557 = 3'h4 == encoders_7_io_output ? proc_4_io_next_header_5 : _GEN_4493; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4558 = 3'h4 == encoders_7_io_output ? proc_4_io_next_header_6 : _GEN_4494; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4559 = 3'h4 == encoders_7_io_output ? proc_4_io_next_header_7 : _GEN_4495; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4560 = 3'h4 == encoders_7_io_output ? proc_4_io_next_header_8 : _GEN_4496; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4561 = 3'h4 == encoders_7_io_output ? proc_4_io_next_header_9 : _GEN_4497; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4562 = 3'h4 == encoders_7_io_output ? proc_4_io_next_header_10 : _GEN_4498; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4563 = 3'h4 == encoders_7_io_output ? proc_4_io_next_header_11 : _GEN_4499; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4564 = 3'h4 == encoders_7_io_output ? proc_4_io_next_header_12 : _GEN_4500; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4565 = 3'h4 == encoders_7_io_output ? proc_4_io_next_header_13 : _GEN_4501; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4566 = 3'h4 == encoders_7_io_output ? proc_4_io_next_header_14 : _GEN_4502; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4567 = 3'h4 == encoders_7_io_output ? proc_4_io_next_header_15 : _GEN_4503; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4568 = 3'h4 == encoders_7_io_output ? proc_4_io_next_header_16 : _GEN_4504; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4569 = 3'h4 == encoders_7_io_output ? proc_4_io_next_header_17 : _GEN_4505; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4570 = 3'h4 == encoders_7_io_output ? proc_4_io_next_header_18 : _GEN_4506; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4571 = 3'h4 == encoders_7_io_output ? proc_4_io_next_header_19 : _GEN_4507; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4572 = 3'h4 == encoders_7_io_output ? proc_4_io_next_header_20 : _GEN_4508; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4573 = 3'h4 == encoders_7_io_output ? proc_4_io_next_header_21 : _GEN_4509; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4574 = 3'h4 == encoders_7_io_output ? proc_4_io_next_header_22 : _GEN_4510; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4575 = 3'h4 == encoders_7_io_output ? proc_4_io_next_header_23 : _GEN_4511; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4576 = 3'h4 == encoders_7_io_output ? proc_4_io_next_header_24 : _GEN_4512; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4577 = 3'h4 == encoders_7_io_output ? proc_4_io_next_header_25 : _GEN_4513; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4578 = 3'h4 == encoders_7_io_output ? proc_4_io_next_header_26 : _GEN_4514; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4579 = 3'h4 == encoders_7_io_output ? proc_4_io_next_header_27 : _GEN_4515; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4580 = 3'h4 == encoders_7_io_output ? proc_4_io_next_header_28 : _GEN_4516; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4581 = 3'h4 == encoders_7_io_output ? proc_4_io_next_header_29 : _GEN_4517; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4582 = 3'h4 == encoders_7_io_output ? proc_4_io_next_header_30 : _GEN_4518; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4583 = 3'h4 == encoders_7_io_output ? proc_4_io_next_header_31 : _GEN_4519; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4584 = 3'h4 == encoders_7_io_output ? proc_4_io_next_header_32 : _GEN_4520; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4585 = 3'h4 == encoders_7_io_output ? proc_4_io_next_header_33 : _GEN_4521; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4586 = 3'h4 == encoders_7_io_output ? proc_4_io_next_header_34 : _GEN_4522; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4587 = 3'h4 == encoders_7_io_output ? proc_4_io_next_header_35 : _GEN_4523; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4588 = 3'h4 == encoders_7_io_output ? proc_4_io_next_header_36 : _GEN_4524; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4589 = 3'h4 == encoders_7_io_output ? proc_4_io_next_header_37 : _GEN_4525; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4590 = 3'h4 == encoders_7_io_output ? proc_4_io_next_header_38 : _GEN_4526; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4591 = 3'h4 == encoders_7_io_output ? proc_4_io_next_header_39 : _GEN_4527; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4592 = 3'h4 == encoders_7_io_output ? proc_4_io_next_header_40 : _GEN_4528; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4593 = 3'h4 == encoders_7_io_output ? proc_4_io_next_header_41 : _GEN_4529; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4594 = 3'h4 == encoders_7_io_output ? proc_4_io_next_header_42 : _GEN_4530; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4595 = 3'h4 == encoders_7_io_output ? proc_4_io_next_header_43 : _GEN_4531; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4596 = 3'h4 == encoders_7_io_output ? proc_4_io_next_header_44 : _GEN_4532; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4597 = 3'h4 == encoders_7_io_output ? proc_4_io_next_header_45 : _GEN_4533; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4598 = 3'h4 == encoders_7_io_output ? proc_4_io_next_header_46 : _GEN_4534; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4599 = 3'h4 == encoders_7_io_output ? proc_4_io_next_header_47 : _GEN_4535; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4600 = 3'h4 == encoders_7_io_output ? proc_4_io_next_header_48 : _GEN_4536; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4601 = 3'h4 == encoders_7_io_output ? proc_4_io_next_header_49 : _GEN_4537; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4602 = 3'h4 == encoders_7_io_output ? proc_4_io_next_header_50 : _GEN_4538; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4603 = 3'h4 == encoders_7_io_output ? proc_4_io_next_header_51 : _GEN_4539; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4604 = 3'h4 == encoders_7_io_output ? proc_4_io_next_header_52 : _GEN_4540; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4605 = 3'h4 == encoders_7_io_output ? proc_4_io_next_header_53 : _GEN_4541; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4606 = 3'h4 == encoders_7_io_output ? proc_4_io_next_header_54 : _GEN_4542; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4607 = 3'h4 == encoders_7_io_output ? proc_4_io_next_header_55 : _GEN_4543; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4608 = 3'h4 == encoders_7_io_output ? proc_4_io_next_header_56 : _GEN_4544; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4609 = 3'h4 == encoders_7_io_output ? proc_4_io_next_header_57 : _GEN_4545; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4610 = 3'h4 == encoders_7_io_output ? proc_4_io_next_header_58 : _GEN_4546; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4611 = 3'h4 == encoders_7_io_output ? proc_4_io_next_header_59 : _GEN_4547; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4612 = 3'h4 == encoders_7_io_output ? proc_4_io_next_header_60 : _GEN_4548; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4613 = 3'h4 == encoders_7_io_output ? proc_4_io_next_header_61 : _GEN_4549; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4614 = 3'h4 == encoders_7_io_output ? proc_4_io_next_header_62 : _GEN_4550; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4615 = 3'h4 == encoders_7_io_output ? proc_4_io_next_header_63 : _GEN_4551; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4616 = 3'h5 == encoders_7_io_output ? proc_5_io_next_header_0 : _GEN_4552; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4617 = 3'h5 == encoders_7_io_output ? proc_5_io_next_header_1 : _GEN_4553; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4618 = 3'h5 == encoders_7_io_output ? proc_5_io_next_header_2 : _GEN_4554; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4619 = 3'h5 == encoders_7_io_output ? proc_5_io_next_header_3 : _GEN_4555; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4620 = 3'h5 == encoders_7_io_output ? proc_5_io_next_header_4 : _GEN_4556; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4621 = 3'h5 == encoders_7_io_output ? proc_5_io_next_header_5 : _GEN_4557; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4622 = 3'h5 == encoders_7_io_output ? proc_5_io_next_header_6 : _GEN_4558; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4623 = 3'h5 == encoders_7_io_output ? proc_5_io_next_header_7 : _GEN_4559; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4624 = 3'h5 == encoders_7_io_output ? proc_5_io_next_header_8 : _GEN_4560; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4625 = 3'h5 == encoders_7_io_output ? proc_5_io_next_header_9 : _GEN_4561; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4626 = 3'h5 == encoders_7_io_output ? proc_5_io_next_header_10 : _GEN_4562; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4627 = 3'h5 == encoders_7_io_output ? proc_5_io_next_header_11 : _GEN_4563; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4628 = 3'h5 == encoders_7_io_output ? proc_5_io_next_header_12 : _GEN_4564; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4629 = 3'h5 == encoders_7_io_output ? proc_5_io_next_header_13 : _GEN_4565; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4630 = 3'h5 == encoders_7_io_output ? proc_5_io_next_header_14 : _GEN_4566; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4631 = 3'h5 == encoders_7_io_output ? proc_5_io_next_header_15 : _GEN_4567; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4632 = 3'h5 == encoders_7_io_output ? proc_5_io_next_header_16 : _GEN_4568; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4633 = 3'h5 == encoders_7_io_output ? proc_5_io_next_header_17 : _GEN_4569; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4634 = 3'h5 == encoders_7_io_output ? proc_5_io_next_header_18 : _GEN_4570; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4635 = 3'h5 == encoders_7_io_output ? proc_5_io_next_header_19 : _GEN_4571; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4636 = 3'h5 == encoders_7_io_output ? proc_5_io_next_header_20 : _GEN_4572; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4637 = 3'h5 == encoders_7_io_output ? proc_5_io_next_header_21 : _GEN_4573; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4638 = 3'h5 == encoders_7_io_output ? proc_5_io_next_header_22 : _GEN_4574; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4639 = 3'h5 == encoders_7_io_output ? proc_5_io_next_header_23 : _GEN_4575; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4640 = 3'h5 == encoders_7_io_output ? proc_5_io_next_header_24 : _GEN_4576; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4641 = 3'h5 == encoders_7_io_output ? proc_5_io_next_header_25 : _GEN_4577; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4642 = 3'h5 == encoders_7_io_output ? proc_5_io_next_header_26 : _GEN_4578; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4643 = 3'h5 == encoders_7_io_output ? proc_5_io_next_header_27 : _GEN_4579; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4644 = 3'h5 == encoders_7_io_output ? proc_5_io_next_header_28 : _GEN_4580; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4645 = 3'h5 == encoders_7_io_output ? proc_5_io_next_header_29 : _GEN_4581; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4646 = 3'h5 == encoders_7_io_output ? proc_5_io_next_header_30 : _GEN_4582; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4647 = 3'h5 == encoders_7_io_output ? proc_5_io_next_header_31 : _GEN_4583; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4648 = 3'h5 == encoders_7_io_output ? proc_5_io_next_header_32 : _GEN_4584; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4649 = 3'h5 == encoders_7_io_output ? proc_5_io_next_header_33 : _GEN_4585; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4650 = 3'h5 == encoders_7_io_output ? proc_5_io_next_header_34 : _GEN_4586; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4651 = 3'h5 == encoders_7_io_output ? proc_5_io_next_header_35 : _GEN_4587; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4652 = 3'h5 == encoders_7_io_output ? proc_5_io_next_header_36 : _GEN_4588; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4653 = 3'h5 == encoders_7_io_output ? proc_5_io_next_header_37 : _GEN_4589; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4654 = 3'h5 == encoders_7_io_output ? proc_5_io_next_header_38 : _GEN_4590; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4655 = 3'h5 == encoders_7_io_output ? proc_5_io_next_header_39 : _GEN_4591; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4656 = 3'h5 == encoders_7_io_output ? proc_5_io_next_header_40 : _GEN_4592; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4657 = 3'h5 == encoders_7_io_output ? proc_5_io_next_header_41 : _GEN_4593; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4658 = 3'h5 == encoders_7_io_output ? proc_5_io_next_header_42 : _GEN_4594; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4659 = 3'h5 == encoders_7_io_output ? proc_5_io_next_header_43 : _GEN_4595; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4660 = 3'h5 == encoders_7_io_output ? proc_5_io_next_header_44 : _GEN_4596; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4661 = 3'h5 == encoders_7_io_output ? proc_5_io_next_header_45 : _GEN_4597; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4662 = 3'h5 == encoders_7_io_output ? proc_5_io_next_header_46 : _GEN_4598; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4663 = 3'h5 == encoders_7_io_output ? proc_5_io_next_header_47 : _GEN_4599; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4664 = 3'h5 == encoders_7_io_output ? proc_5_io_next_header_48 : _GEN_4600; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4665 = 3'h5 == encoders_7_io_output ? proc_5_io_next_header_49 : _GEN_4601; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4666 = 3'h5 == encoders_7_io_output ? proc_5_io_next_header_50 : _GEN_4602; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4667 = 3'h5 == encoders_7_io_output ? proc_5_io_next_header_51 : _GEN_4603; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4668 = 3'h5 == encoders_7_io_output ? proc_5_io_next_header_52 : _GEN_4604; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4669 = 3'h5 == encoders_7_io_output ? proc_5_io_next_header_53 : _GEN_4605; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4670 = 3'h5 == encoders_7_io_output ? proc_5_io_next_header_54 : _GEN_4606; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4671 = 3'h5 == encoders_7_io_output ? proc_5_io_next_header_55 : _GEN_4607; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4672 = 3'h5 == encoders_7_io_output ? proc_5_io_next_header_56 : _GEN_4608; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4673 = 3'h5 == encoders_7_io_output ? proc_5_io_next_header_57 : _GEN_4609; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4674 = 3'h5 == encoders_7_io_output ? proc_5_io_next_header_58 : _GEN_4610; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4675 = 3'h5 == encoders_7_io_output ? proc_5_io_next_header_59 : _GEN_4611; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4676 = 3'h5 == encoders_7_io_output ? proc_5_io_next_header_60 : _GEN_4612; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4677 = 3'h5 == encoders_7_io_output ? proc_5_io_next_header_61 : _GEN_4613; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4678 = 3'h5 == encoders_7_io_output ? proc_5_io_next_header_62 : _GEN_4614; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4679 = 3'h5 == encoders_7_io_output ? proc_5_io_next_header_63 : _GEN_4615; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4680 = 3'h6 == encoders_7_io_output ? proc_6_io_next_header_0 : _GEN_4616; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4681 = 3'h6 == encoders_7_io_output ? proc_6_io_next_header_1 : _GEN_4617; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4682 = 3'h6 == encoders_7_io_output ? proc_6_io_next_header_2 : _GEN_4618; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4683 = 3'h6 == encoders_7_io_output ? proc_6_io_next_header_3 : _GEN_4619; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4684 = 3'h6 == encoders_7_io_output ? proc_6_io_next_header_4 : _GEN_4620; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4685 = 3'h6 == encoders_7_io_output ? proc_6_io_next_header_5 : _GEN_4621; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4686 = 3'h6 == encoders_7_io_output ? proc_6_io_next_header_6 : _GEN_4622; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4687 = 3'h6 == encoders_7_io_output ? proc_6_io_next_header_7 : _GEN_4623; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4688 = 3'h6 == encoders_7_io_output ? proc_6_io_next_header_8 : _GEN_4624; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4689 = 3'h6 == encoders_7_io_output ? proc_6_io_next_header_9 : _GEN_4625; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4690 = 3'h6 == encoders_7_io_output ? proc_6_io_next_header_10 : _GEN_4626; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4691 = 3'h6 == encoders_7_io_output ? proc_6_io_next_header_11 : _GEN_4627; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4692 = 3'h6 == encoders_7_io_output ? proc_6_io_next_header_12 : _GEN_4628; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4693 = 3'h6 == encoders_7_io_output ? proc_6_io_next_header_13 : _GEN_4629; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4694 = 3'h6 == encoders_7_io_output ? proc_6_io_next_header_14 : _GEN_4630; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4695 = 3'h6 == encoders_7_io_output ? proc_6_io_next_header_15 : _GEN_4631; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4696 = 3'h6 == encoders_7_io_output ? proc_6_io_next_header_16 : _GEN_4632; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4697 = 3'h6 == encoders_7_io_output ? proc_6_io_next_header_17 : _GEN_4633; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4698 = 3'h6 == encoders_7_io_output ? proc_6_io_next_header_18 : _GEN_4634; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4699 = 3'h6 == encoders_7_io_output ? proc_6_io_next_header_19 : _GEN_4635; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4700 = 3'h6 == encoders_7_io_output ? proc_6_io_next_header_20 : _GEN_4636; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4701 = 3'h6 == encoders_7_io_output ? proc_6_io_next_header_21 : _GEN_4637; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4702 = 3'h6 == encoders_7_io_output ? proc_6_io_next_header_22 : _GEN_4638; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4703 = 3'h6 == encoders_7_io_output ? proc_6_io_next_header_23 : _GEN_4639; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4704 = 3'h6 == encoders_7_io_output ? proc_6_io_next_header_24 : _GEN_4640; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4705 = 3'h6 == encoders_7_io_output ? proc_6_io_next_header_25 : _GEN_4641; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4706 = 3'h6 == encoders_7_io_output ? proc_6_io_next_header_26 : _GEN_4642; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4707 = 3'h6 == encoders_7_io_output ? proc_6_io_next_header_27 : _GEN_4643; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4708 = 3'h6 == encoders_7_io_output ? proc_6_io_next_header_28 : _GEN_4644; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4709 = 3'h6 == encoders_7_io_output ? proc_6_io_next_header_29 : _GEN_4645; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4710 = 3'h6 == encoders_7_io_output ? proc_6_io_next_header_30 : _GEN_4646; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4711 = 3'h6 == encoders_7_io_output ? proc_6_io_next_header_31 : _GEN_4647; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4712 = 3'h6 == encoders_7_io_output ? proc_6_io_next_header_32 : _GEN_4648; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4713 = 3'h6 == encoders_7_io_output ? proc_6_io_next_header_33 : _GEN_4649; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4714 = 3'h6 == encoders_7_io_output ? proc_6_io_next_header_34 : _GEN_4650; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4715 = 3'h6 == encoders_7_io_output ? proc_6_io_next_header_35 : _GEN_4651; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4716 = 3'h6 == encoders_7_io_output ? proc_6_io_next_header_36 : _GEN_4652; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4717 = 3'h6 == encoders_7_io_output ? proc_6_io_next_header_37 : _GEN_4653; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4718 = 3'h6 == encoders_7_io_output ? proc_6_io_next_header_38 : _GEN_4654; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4719 = 3'h6 == encoders_7_io_output ? proc_6_io_next_header_39 : _GEN_4655; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4720 = 3'h6 == encoders_7_io_output ? proc_6_io_next_header_40 : _GEN_4656; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4721 = 3'h6 == encoders_7_io_output ? proc_6_io_next_header_41 : _GEN_4657; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4722 = 3'h6 == encoders_7_io_output ? proc_6_io_next_header_42 : _GEN_4658; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4723 = 3'h6 == encoders_7_io_output ? proc_6_io_next_header_43 : _GEN_4659; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4724 = 3'h6 == encoders_7_io_output ? proc_6_io_next_header_44 : _GEN_4660; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4725 = 3'h6 == encoders_7_io_output ? proc_6_io_next_header_45 : _GEN_4661; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4726 = 3'h6 == encoders_7_io_output ? proc_6_io_next_header_46 : _GEN_4662; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4727 = 3'h6 == encoders_7_io_output ? proc_6_io_next_header_47 : _GEN_4663; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4728 = 3'h6 == encoders_7_io_output ? proc_6_io_next_header_48 : _GEN_4664; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4729 = 3'h6 == encoders_7_io_output ? proc_6_io_next_header_49 : _GEN_4665; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4730 = 3'h6 == encoders_7_io_output ? proc_6_io_next_header_50 : _GEN_4666; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4731 = 3'h6 == encoders_7_io_output ? proc_6_io_next_header_51 : _GEN_4667; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4732 = 3'h6 == encoders_7_io_output ? proc_6_io_next_header_52 : _GEN_4668; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4733 = 3'h6 == encoders_7_io_output ? proc_6_io_next_header_53 : _GEN_4669; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4734 = 3'h6 == encoders_7_io_output ? proc_6_io_next_header_54 : _GEN_4670; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4735 = 3'h6 == encoders_7_io_output ? proc_6_io_next_header_55 : _GEN_4671; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4736 = 3'h6 == encoders_7_io_output ? proc_6_io_next_header_56 : _GEN_4672; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4737 = 3'h6 == encoders_7_io_output ? proc_6_io_next_header_57 : _GEN_4673; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4738 = 3'h6 == encoders_7_io_output ? proc_6_io_next_header_58 : _GEN_4674; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4739 = 3'h6 == encoders_7_io_output ? proc_6_io_next_header_59 : _GEN_4675; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4740 = 3'h6 == encoders_7_io_output ? proc_6_io_next_header_60 : _GEN_4676; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4741 = 3'h6 == encoders_7_io_output ? proc_6_io_next_header_61 : _GEN_4677; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4742 = 3'h6 == encoders_7_io_output ? proc_6_io_next_header_62 : _GEN_4678; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4743 = 3'h6 == encoders_7_io_output ? proc_6_io_next_header_63 : _GEN_4679; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4744 = 3'h7 == encoders_7_io_output ? proc_7_io_next_header_0 : _GEN_4680; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4745 = 3'h7 == encoders_7_io_output ? proc_7_io_next_header_1 : _GEN_4681; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4746 = 3'h7 == encoders_7_io_output ? proc_7_io_next_header_2 : _GEN_4682; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4747 = 3'h7 == encoders_7_io_output ? proc_7_io_next_header_3 : _GEN_4683; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4748 = 3'h7 == encoders_7_io_output ? proc_7_io_next_header_4 : _GEN_4684; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4749 = 3'h7 == encoders_7_io_output ? proc_7_io_next_header_5 : _GEN_4685; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4750 = 3'h7 == encoders_7_io_output ? proc_7_io_next_header_6 : _GEN_4686; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4751 = 3'h7 == encoders_7_io_output ? proc_7_io_next_header_7 : _GEN_4687; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4752 = 3'h7 == encoders_7_io_output ? proc_7_io_next_header_8 : _GEN_4688; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4753 = 3'h7 == encoders_7_io_output ? proc_7_io_next_header_9 : _GEN_4689; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4754 = 3'h7 == encoders_7_io_output ? proc_7_io_next_header_10 : _GEN_4690; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4755 = 3'h7 == encoders_7_io_output ? proc_7_io_next_header_11 : _GEN_4691; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4756 = 3'h7 == encoders_7_io_output ? proc_7_io_next_header_12 : _GEN_4692; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4757 = 3'h7 == encoders_7_io_output ? proc_7_io_next_header_13 : _GEN_4693; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4758 = 3'h7 == encoders_7_io_output ? proc_7_io_next_header_14 : _GEN_4694; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4759 = 3'h7 == encoders_7_io_output ? proc_7_io_next_header_15 : _GEN_4695; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4760 = 3'h7 == encoders_7_io_output ? proc_7_io_next_header_16 : _GEN_4696; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4761 = 3'h7 == encoders_7_io_output ? proc_7_io_next_header_17 : _GEN_4697; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4762 = 3'h7 == encoders_7_io_output ? proc_7_io_next_header_18 : _GEN_4698; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4763 = 3'h7 == encoders_7_io_output ? proc_7_io_next_header_19 : _GEN_4699; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4764 = 3'h7 == encoders_7_io_output ? proc_7_io_next_header_20 : _GEN_4700; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4765 = 3'h7 == encoders_7_io_output ? proc_7_io_next_header_21 : _GEN_4701; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4766 = 3'h7 == encoders_7_io_output ? proc_7_io_next_header_22 : _GEN_4702; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4767 = 3'h7 == encoders_7_io_output ? proc_7_io_next_header_23 : _GEN_4703; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4768 = 3'h7 == encoders_7_io_output ? proc_7_io_next_header_24 : _GEN_4704; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4769 = 3'h7 == encoders_7_io_output ? proc_7_io_next_header_25 : _GEN_4705; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4770 = 3'h7 == encoders_7_io_output ? proc_7_io_next_header_26 : _GEN_4706; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4771 = 3'h7 == encoders_7_io_output ? proc_7_io_next_header_27 : _GEN_4707; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4772 = 3'h7 == encoders_7_io_output ? proc_7_io_next_header_28 : _GEN_4708; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4773 = 3'h7 == encoders_7_io_output ? proc_7_io_next_header_29 : _GEN_4709; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4774 = 3'h7 == encoders_7_io_output ? proc_7_io_next_header_30 : _GEN_4710; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4775 = 3'h7 == encoders_7_io_output ? proc_7_io_next_header_31 : _GEN_4711; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4776 = 3'h7 == encoders_7_io_output ? proc_7_io_next_header_32 : _GEN_4712; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4777 = 3'h7 == encoders_7_io_output ? proc_7_io_next_header_33 : _GEN_4713; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4778 = 3'h7 == encoders_7_io_output ? proc_7_io_next_header_34 : _GEN_4714; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4779 = 3'h7 == encoders_7_io_output ? proc_7_io_next_header_35 : _GEN_4715; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4780 = 3'h7 == encoders_7_io_output ? proc_7_io_next_header_36 : _GEN_4716; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4781 = 3'h7 == encoders_7_io_output ? proc_7_io_next_header_37 : _GEN_4717; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4782 = 3'h7 == encoders_7_io_output ? proc_7_io_next_header_38 : _GEN_4718; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4783 = 3'h7 == encoders_7_io_output ? proc_7_io_next_header_39 : _GEN_4719; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4784 = 3'h7 == encoders_7_io_output ? proc_7_io_next_header_40 : _GEN_4720; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4785 = 3'h7 == encoders_7_io_output ? proc_7_io_next_header_41 : _GEN_4721; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4786 = 3'h7 == encoders_7_io_output ? proc_7_io_next_header_42 : _GEN_4722; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4787 = 3'h7 == encoders_7_io_output ? proc_7_io_next_header_43 : _GEN_4723; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4788 = 3'h7 == encoders_7_io_output ? proc_7_io_next_header_44 : _GEN_4724; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4789 = 3'h7 == encoders_7_io_output ? proc_7_io_next_header_45 : _GEN_4725; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4790 = 3'h7 == encoders_7_io_output ? proc_7_io_next_header_46 : _GEN_4726; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4791 = 3'h7 == encoders_7_io_output ? proc_7_io_next_header_47 : _GEN_4727; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4792 = 3'h7 == encoders_7_io_output ? proc_7_io_next_header_48 : _GEN_4728; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4793 = 3'h7 == encoders_7_io_output ? proc_7_io_next_header_49 : _GEN_4729; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4794 = 3'h7 == encoders_7_io_output ? proc_7_io_next_header_50 : _GEN_4730; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4795 = 3'h7 == encoders_7_io_output ? proc_7_io_next_header_51 : _GEN_4731; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4796 = 3'h7 == encoders_7_io_output ? proc_7_io_next_header_52 : _GEN_4732; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4797 = 3'h7 == encoders_7_io_output ? proc_7_io_next_header_53 : _GEN_4733; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4798 = 3'h7 == encoders_7_io_output ? proc_7_io_next_header_54 : _GEN_4734; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4799 = 3'h7 == encoders_7_io_output ? proc_7_io_next_header_55 : _GEN_4735; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4800 = 3'h7 == encoders_7_io_output ? proc_7_io_next_header_56 : _GEN_4736; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4801 = 3'h7 == encoders_7_io_output ? proc_7_io_next_header_57 : _GEN_4737; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4802 = 3'h7 == encoders_7_io_output ? proc_7_io_next_header_58 : _GEN_4738; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4803 = 3'h7 == encoders_7_io_output ? proc_7_io_next_header_59 : _GEN_4739; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4804 = 3'h7 == encoders_7_io_output ? proc_7_io_next_header_60 : _GEN_4740; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4805 = 3'h7 == encoders_7_io_output ? proc_7_io_next_header_61 : _GEN_4741; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4806 = 3'h7 == encoders_7_io_output ? proc_7_io_next_header_62 : _GEN_4742; // @[controller.scala 94:46 controller.scala 95:46]
  wire [7:0] _GEN_4807 = 3'h7 == encoders_7_io_output ? proc_7_io_next_header_63 : _GEN_4743; // @[controller.scala 94:46 controller.scala 95:46]
  SRAM mem_0 ( // @[controller.scala 18:25]
    .clock(mem_0_clock),
    .io_mem_a_addr(mem_0_io_mem_a_addr),
    .io_mem_a_rdata(mem_0_io_mem_a_rdata),
    .io_mem_b_addr(mem_0_io_mem_b_addr),
    .io_mem_b_rdata(mem_0_io_mem_b_rdata)
  );
  SRAM mem_1 ( // @[controller.scala 18:25]
    .clock(mem_1_clock),
    .io_mem_a_addr(mem_1_io_mem_a_addr),
    .io_mem_a_rdata(mem_1_io_mem_a_rdata),
    .io_mem_b_addr(mem_1_io_mem_b_addr),
    .io_mem_b_rdata(mem_1_io_mem_b_rdata)
  );
  SRAM mem_2 ( // @[controller.scala 18:25]
    .clock(mem_2_clock),
    .io_mem_a_addr(mem_2_io_mem_a_addr),
    .io_mem_a_rdata(mem_2_io_mem_a_rdata),
    .io_mem_b_addr(mem_2_io_mem_b_addr),
    .io_mem_b_rdata(mem_2_io_mem_b_rdata)
  );
  SRAM mem_3 ( // @[controller.scala 18:25]
    .clock(mem_3_clock),
    .io_mem_a_addr(mem_3_io_mem_a_addr),
    .io_mem_a_rdata(mem_3_io_mem_a_rdata),
    .io_mem_b_addr(mem_3_io_mem_b_addr),
    .io_mem_b_rdata(mem_3_io_mem_b_rdata)
  );
  Encoder83 encoders_0 ( // @[controller.scala 23:25]
    .io_input(encoders_0_io_input),
    .io_output(encoders_0_io_output),
    .io_valid(encoders_0_io_valid)
  );
  Encoder83 encoders_1 ( // @[controller.scala 23:25]
    .io_input(encoders_1_io_input),
    .io_output(encoders_1_io_output),
    .io_valid(encoders_1_io_valid)
  );
  Encoder83 encoders_2 ( // @[controller.scala 23:25]
    .io_input(encoders_2_io_input),
    .io_output(encoders_2_io_output),
    .io_valid(encoders_2_io_valid)
  );
  Encoder83 encoders_3 ( // @[controller.scala 23:25]
    .io_input(encoders_3_io_input),
    .io_output(encoders_3_io_output),
    .io_valid(encoders_3_io_valid)
  );
  Encoder83 encoders_4 ( // @[controller.scala 23:25]
    .io_input(encoders_4_io_input),
    .io_output(encoders_4_io_output),
    .io_valid(encoders_4_io_valid)
  );
  Encoder83 encoders_5 ( // @[controller.scala 23:25]
    .io_input(encoders_5_io_input),
    .io_output(encoders_5_io_output),
    .io_valid(encoders_5_io_valid)
  );
  Encoder83 encoders_6 ( // @[controller.scala 23:25]
    .io_input(encoders_6_io_input),
    .io_output(encoders_6_io_output),
    .io_valid(encoders_6_io_valid)
  );
  Encoder83 encoders_7 ( // @[controller.scala 23:25]
    .io_input(encoders_7_io_input),
    .io_output(encoders_7_io_output),
    .io_valid(encoders_7_io_valid)
  );
  ProcessorController proc_0 ( // @[controller.scala 29:25]
    .clock(proc_0_clock),
    .reset(proc_0_reset),
    .io_update(proc_0_io_update),
    .io_packet_header_0(proc_0_io_packet_header_0),
    .io_packet_header_1(proc_0_io_packet_header_1),
    .io_packet_header_2(proc_0_io_packet_header_2),
    .io_packet_header_3(proc_0_io_packet_header_3),
    .io_packet_header_4(proc_0_io_packet_header_4),
    .io_packet_header_5(proc_0_io_packet_header_5),
    .io_packet_header_6(proc_0_io_packet_header_6),
    .io_packet_header_7(proc_0_io_packet_header_7),
    .io_packet_header_8(proc_0_io_packet_header_8),
    .io_packet_header_9(proc_0_io_packet_header_9),
    .io_packet_header_10(proc_0_io_packet_header_10),
    .io_packet_header_11(proc_0_io_packet_header_11),
    .io_packet_header_12(proc_0_io_packet_header_12),
    .io_packet_header_13(proc_0_io_packet_header_13),
    .io_packet_header_14(proc_0_io_packet_header_14),
    .io_packet_header_15(proc_0_io_packet_header_15),
    .io_packet_header_16(proc_0_io_packet_header_16),
    .io_packet_header_17(proc_0_io_packet_header_17),
    .io_packet_header_18(proc_0_io_packet_header_18),
    .io_packet_header_19(proc_0_io_packet_header_19),
    .io_packet_header_20(proc_0_io_packet_header_20),
    .io_packet_header_21(proc_0_io_packet_header_21),
    .io_packet_header_22(proc_0_io_packet_header_22),
    .io_packet_header_23(proc_0_io_packet_header_23),
    .io_packet_header_24(proc_0_io_packet_header_24),
    .io_packet_header_25(proc_0_io_packet_header_25),
    .io_packet_header_26(proc_0_io_packet_header_26),
    .io_packet_header_27(proc_0_io_packet_header_27),
    .io_packet_header_28(proc_0_io_packet_header_28),
    .io_packet_header_29(proc_0_io_packet_header_29),
    .io_packet_header_30(proc_0_io_packet_header_30),
    .io_packet_header_31(proc_0_io_packet_header_31),
    .io_packet_header_32(proc_0_io_packet_header_32),
    .io_packet_header_33(proc_0_io_packet_header_33),
    .io_packet_header_34(proc_0_io_packet_header_34),
    .io_packet_header_35(proc_0_io_packet_header_35),
    .io_packet_header_36(proc_0_io_packet_header_36),
    .io_packet_header_37(proc_0_io_packet_header_37),
    .io_packet_header_38(proc_0_io_packet_header_38),
    .io_packet_header_39(proc_0_io_packet_header_39),
    .io_packet_header_40(proc_0_io_packet_header_40),
    .io_packet_header_41(proc_0_io_packet_header_41),
    .io_packet_header_42(proc_0_io_packet_header_42),
    .io_packet_header_43(proc_0_io_packet_header_43),
    .io_packet_header_44(proc_0_io_packet_header_44),
    .io_packet_header_45(proc_0_io_packet_header_45),
    .io_packet_header_46(proc_0_io_packet_header_46),
    .io_packet_header_47(proc_0_io_packet_header_47),
    .io_packet_header_48(proc_0_io_packet_header_48),
    .io_packet_header_49(proc_0_io_packet_header_49),
    .io_packet_header_50(proc_0_io_packet_header_50),
    .io_packet_header_51(proc_0_io_packet_header_51),
    .io_packet_header_52(proc_0_io_packet_header_52),
    .io_packet_header_53(proc_0_io_packet_header_53),
    .io_packet_header_54(proc_0_io_packet_header_54),
    .io_packet_header_55(proc_0_io_packet_header_55),
    .io_packet_header_56(proc_0_io_packet_header_56),
    .io_packet_header_57(proc_0_io_packet_header_57),
    .io_packet_header_58(proc_0_io_packet_header_58),
    .io_packet_header_59(proc_0_io_packet_header_59),
    .io_packet_header_60(proc_0_io_packet_header_60),
    .io_packet_header_61(proc_0_io_packet_header_61),
    .io_packet_header_62(proc_0_io_packet_header_62),
    .io_packet_header_63(proc_0_io_packet_header_63),
    .io_end(proc_0_io_end),
    .io_mem_addr(proc_0_io_mem_addr),
    .io_mem_rdata(proc_0_io_mem_rdata),
    .io_ready(proc_0_io_ready),
    .io_mod_start(proc_0_io_mod_start),
    .io_mod_hit_action_addr(proc_0_io_mod_hit_action_addr),
    .io_mod_miss_action_addr(proc_0_io_mod_miss_action_addr),
    .io_mod_ps_mod_start(proc_0_io_mod_ps_mod_start),
    .io_mod_ps_mod_header_id(proc_0_io_mod_ps_mod_header_id),
    .io_mod_ps_mod_header_length(proc_0_io_mod_ps_mod_header_length),
    .io_mod_ps_mod_next_tag_start(proc_0_io_mod_ps_mod_next_tag_start),
    .io_mod_ps_mod_next_table_0(proc_0_io_mod_ps_mod_next_table_0),
    .io_mod_ps_mod_next_table_1(proc_0_io_mod_ps_mod_next_table_1),
    .io_mod_mt_mod_start(proc_0_io_mod_mt_mod_start),
    .io_mod_mt_mod_header_id(proc_0_io_mod_mt_mod_header_id),
    .io_mod_mt_mod_key_off(proc_0_io_mod_mt_mod_key_off),
    .io_mod_mt_mod_key_len(proc_0_io_mod_mt_mod_key_len),
    .io_mod_mt_mod_val_len(proc_0_io_mod_mt_mod_val_len),
    .io_mod_ex_mod_start(proc_0_io_mod_ex_mod_start),
    .io_mod_ex_mod_ops_0(proc_0_io_mod_ex_mod_ops_0),
    .io_mod_ex_mod_ops_1(proc_0_io_mod_ex_mod_ops_1),
    .io_mod_ex_mod_ops_2(proc_0_io_mod_ex_mod_ops_2),
    .io_mod_ex_mod_ops_3(proc_0_io_mod_ex_mod_ops_3),
    .io_mod_ex_mod_ops_4(proc_0_io_mod_ex_mod_ops_4),
    .io_mod_ex_mod_ops_5(proc_0_io_mod_ex_mod_ops_5),
    .io_mod_ex_mod_ops_6(proc_0_io_mod_ex_mod_ops_6),
    .io_mod_ex_mod_ops_7(proc_0_io_mod_ex_mod_ops_7),
    .io_mod_ex_mod_ops_8(proc_0_io_mod_ex_mod_ops_8),
    .io_mod_ex_mod_ops_9(proc_0_io_mod_ex_mod_ops_9),
    .io_mod_ex_mod_ops_10(proc_0_io_mod_ex_mod_ops_10),
    .io_mod_ex_mod_ops_11(proc_0_io_mod_ex_mod_ops_11),
    .io_mod_ex_mod_ops_12(proc_0_io_mod_ex_mod_ops_12),
    .io_mod_ex_mod_ops_13(proc_0_io_mod_ex_mod_ops_13),
    .io_mod_ex_mod_ops_14(proc_0_io_mod_ex_mod_ops_14),
    .io_mod_ex_mod_ops_15(proc_0_io_mod_ex_mod_ops_15),
    .io_next_en(proc_0_io_next_en),
    .io_next_header_0(proc_0_io_next_header_0),
    .io_next_header_1(proc_0_io_next_header_1),
    .io_next_header_2(proc_0_io_next_header_2),
    .io_next_header_3(proc_0_io_next_header_3),
    .io_next_header_4(proc_0_io_next_header_4),
    .io_next_header_5(proc_0_io_next_header_5),
    .io_next_header_6(proc_0_io_next_header_6),
    .io_next_header_7(proc_0_io_next_header_7),
    .io_next_header_8(proc_0_io_next_header_8),
    .io_next_header_9(proc_0_io_next_header_9),
    .io_next_header_10(proc_0_io_next_header_10),
    .io_next_header_11(proc_0_io_next_header_11),
    .io_next_header_12(proc_0_io_next_header_12),
    .io_next_header_13(proc_0_io_next_header_13),
    .io_next_header_14(proc_0_io_next_header_14),
    .io_next_header_15(proc_0_io_next_header_15),
    .io_next_header_16(proc_0_io_next_header_16),
    .io_next_header_17(proc_0_io_next_header_17),
    .io_next_header_18(proc_0_io_next_header_18),
    .io_next_header_19(proc_0_io_next_header_19),
    .io_next_header_20(proc_0_io_next_header_20),
    .io_next_header_21(proc_0_io_next_header_21),
    .io_next_header_22(proc_0_io_next_header_22),
    .io_next_header_23(proc_0_io_next_header_23),
    .io_next_header_24(proc_0_io_next_header_24),
    .io_next_header_25(proc_0_io_next_header_25),
    .io_next_header_26(proc_0_io_next_header_26),
    .io_next_header_27(proc_0_io_next_header_27),
    .io_next_header_28(proc_0_io_next_header_28),
    .io_next_header_29(proc_0_io_next_header_29),
    .io_next_header_30(proc_0_io_next_header_30),
    .io_next_header_31(proc_0_io_next_header_31),
    .io_next_header_32(proc_0_io_next_header_32),
    .io_next_header_33(proc_0_io_next_header_33),
    .io_next_header_34(proc_0_io_next_header_34),
    .io_next_header_35(proc_0_io_next_header_35),
    .io_next_header_36(proc_0_io_next_header_36),
    .io_next_header_37(proc_0_io_next_header_37),
    .io_next_header_38(proc_0_io_next_header_38),
    .io_next_header_39(proc_0_io_next_header_39),
    .io_next_header_40(proc_0_io_next_header_40),
    .io_next_header_41(proc_0_io_next_header_41),
    .io_next_header_42(proc_0_io_next_header_42),
    .io_next_header_43(proc_0_io_next_header_43),
    .io_next_header_44(proc_0_io_next_header_44),
    .io_next_header_45(proc_0_io_next_header_45),
    .io_next_header_46(proc_0_io_next_header_46),
    .io_next_header_47(proc_0_io_next_header_47),
    .io_next_header_48(proc_0_io_next_header_48),
    .io_next_header_49(proc_0_io_next_header_49),
    .io_next_header_50(proc_0_io_next_header_50),
    .io_next_header_51(proc_0_io_next_header_51),
    .io_next_header_52(proc_0_io_next_header_52),
    .io_next_header_53(proc_0_io_next_header_53),
    .io_next_header_54(proc_0_io_next_header_54),
    .io_next_header_55(proc_0_io_next_header_55),
    .io_next_header_56(proc_0_io_next_header_56),
    .io_next_header_57(proc_0_io_next_header_57),
    .io_next_header_58(proc_0_io_next_header_58),
    .io_next_header_59(proc_0_io_next_header_59),
    .io_next_header_60(proc_0_io_next_header_60),
    .io_next_header_61(proc_0_io_next_header_61),
    .io_next_header_62(proc_0_io_next_header_62),
    .io_next_header_63(proc_0_io_next_header_63),
    .io_next_proc(proc_0_io_next_proc)
  );
  ProcessorController proc_1 ( // @[controller.scala 29:25]
    .clock(proc_1_clock),
    .reset(proc_1_reset),
    .io_update(proc_1_io_update),
    .io_packet_header_0(proc_1_io_packet_header_0),
    .io_packet_header_1(proc_1_io_packet_header_1),
    .io_packet_header_2(proc_1_io_packet_header_2),
    .io_packet_header_3(proc_1_io_packet_header_3),
    .io_packet_header_4(proc_1_io_packet_header_4),
    .io_packet_header_5(proc_1_io_packet_header_5),
    .io_packet_header_6(proc_1_io_packet_header_6),
    .io_packet_header_7(proc_1_io_packet_header_7),
    .io_packet_header_8(proc_1_io_packet_header_8),
    .io_packet_header_9(proc_1_io_packet_header_9),
    .io_packet_header_10(proc_1_io_packet_header_10),
    .io_packet_header_11(proc_1_io_packet_header_11),
    .io_packet_header_12(proc_1_io_packet_header_12),
    .io_packet_header_13(proc_1_io_packet_header_13),
    .io_packet_header_14(proc_1_io_packet_header_14),
    .io_packet_header_15(proc_1_io_packet_header_15),
    .io_packet_header_16(proc_1_io_packet_header_16),
    .io_packet_header_17(proc_1_io_packet_header_17),
    .io_packet_header_18(proc_1_io_packet_header_18),
    .io_packet_header_19(proc_1_io_packet_header_19),
    .io_packet_header_20(proc_1_io_packet_header_20),
    .io_packet_header_21(proc_1_io_packet_header_21),
    .io_packet_header_22(proc_1_io_packet_header_22),
    .io_packet_header_23(proc_1_io_packet_header_23),
    .io_packet_header_24(proc_1_io_packet_header_24),
    .io_packet_header_25(proc_1_io_packet_header_25),
    .io_packet_header_26(proc_1_io_packet_header_26),
    .io_packet_header_27(proc_1_io_packet_header_27),
    .io_packet_header_28(proc_1_io_packet_header_28),
    .io_packet_header_29(proc_1_io_packet_header_29),
    .io_packet_header_30(proc_1_io_packet_header_30),
    .io_packet_header_31(proc_1_io_packet_header_31),
    .io_packet_header_32(proc_1_io_packet_header_32),
    .io_packet_header_33(proc_1_io_packet_header_33),
    .io_packet_header_34(proc_1_io_packet_header_34),
    .io_packet_header_35(proc_1_io_packet_header_35),
    .io_packet_header_36(proc_1_io_packet_header_36),
    .io_packet_header_37(proc_1_io_packet_header_37),
    .io_packet_header_38(proc_1_io_packet_header_38),
    .io_packet_header_39(proc_1_io_packet_header_39),
    .io_packet_header_40(proc_1_io_packet_header_40),
    .io_packet_header_41(proc_1_io_packet_header_41),
    .io_packet_header_42(proc_1_io_packet_header_42),
    .io_packet_header_43(proc_1_io_packet_header_43),
    .io_packet_header_44(proc_1_io_packet_header_44),
    .io_packet_header_45(proc_1_io_packet_header_45),
    .io_packet_header_46(proc_1_io_packet_header_46),
    .io_packet_header_47(proc_1_io_packet_header_47),
    .io_packet_header_48(proc_1_io_packet_header_48),
    .io_packet_header_49(proc_1_io_packet_header_49),
    .io_packet_header_50(proc_1_io_packet_header_50),
    .io_packet_header_51(proc_1_io_packet_header_51),
    .io_packet_header_52(proc_1_io_packet_header_52),
    .io_packet_header_53(proc_1_io_packet_header_53),
    .io_packet_header_54(proc_1_io_packet_header_54),
    .io_packet_header_55(proc_1_io_packet_header_55),
    .io_packet_header_56(proc_1_io_packet_header_56),
    .io_packet_header_57(proc_1_io_packet_header_57),
    .io_packet_header_58(proc_1_io_packet_header_58),
    .io_packet_header_59(proc_1_io_packet_header_59),
    .io_packet_header_60(proc_1_io_packet_header_60),
    .io_packet_header_61(proc_1_io_packet_header_61),
    .io_packet_header_62(proc_1_io_packet_header_62),
    .io_packet_header_63(proc_1_io_packet_header_63),
    .io_end(proc_1_io_end),
    .io_mem_addr(proc_1_io_mem_addr),
    .io_mem_rdata(proc_1_io_mem_rdata),
    .io_ready(proc_1_io_ready),
    .io_mod_start(proc_1_io_mod_start),
    .io_mod_hit_action_addr(proc_1_io_mod_hit_action_addr),
    .io_mod_miss_action_addr(proc_1_io_mod_miss_action_addr),
    .io_mod_ps_mod_start(proc_1_io_mod_ps_mod_start),
    .io_mod_ps_mod_header_id(proc_1_io_mod_ps_mod_header_id),
    .io_mod_ps_mod_header_length(proc_1_io_mod_ps_mod_header_length),
    .io_mod_ps_mod_next_tag_start(proc_1_io_mod_ps_mod_next_tag_start),
    .io_mod_ps_mod_next_table_0(proc_1_io_mod_ps_mod_next_table_0),
    .io_mod_ps_mod_next_table_1(proc_1_io_mod_ps_mod_next_table_1),
    .io_mod_mt_mod_start(proc_1_io_mod_mt_mod_start),
    .io_mod_mt_mod_header_id(proc_1_io_mod_mt_mod_header_id),
    .io_mod_mt_mod_key_off(proc_1_io_mod_mt_mod_key_off),
    .io_mod_mt_mod_key_len(proc_1_io_mod_mt_mod_key_len),
    .io_mod_mt_mod_val_len(proc_1_io_mod_mt_mod_val_len),
    .io_mod_ex_mod_start(proc_1_io_mod_ex_mod_start),
    .io_mod_ex_mod_ops_0(proc_1_io_mod_ex_mod_ops_0),
    .io_mod_ex_mod_ops_1(proc_1_io_mod_ex_mod_ops_1),
    .io_mod_ex_mod_ops_2(proc_1_io_mod_ex_mod_ops_2),
    .io_mod_ex_mod_ops_3(proc_1_io_mod_ex_mod_ops_3),
    .io_mod_ex_mod_ops_4(proc_1_io_mod_ex_mod_ops_4),
    .io_mod_ex_mod_ops_5(proc_1_io_mod_ex_mod_ops_5),
    .io_mod_ex_mod_ops_6(proc_1_io_mod_ex_mod_ops_6),
    .io_mod_ex_mod_ops_7(proc_1_io_mod_ex_mod_ops_7),
    .io_mod_ex_mod_ops_8(proc_1_io_mod_ex_mod_ops_8),
    .io_mod_ex_mod_ops_9(proc_1_io_mod_ex_mod_ops_9),
    .io_mod_ex_mod_ops_10(proc_1_io_mod_ex_mod_ops_10),
    .io_mod_ex_mod_ops_11(proc_1_io_mod_ex_mod_ops_11),
    .io_mod_ex_mod_ops_12(proc_1_io_mod_ex_mod_ops_12),
    .io_mod_ex_mod_ops_13(proc_1_io_mod_ex_mod_ops_13),
    .io_mod_ex_mod_ops_14(proc_1_io_mod_ex_mod_ops_14),
    .io_mod_ex_mod_ops_15(proc_1_io_mod_ex_mod_ops_15),
    .io_next_en(proc_1_io_next_en),
    .io_next_header_0(proc_1_io_next_header_0),
    .io_next_header_1(proc_1_io_next_header_1),
    .io_next_header_2(proc_1_io_next_header_2),
    .io_next_header_3(proc_1_io_next_header_3),
    .io_next_header_4(proc_1_io_next_header_4),
    .io_next_header_5(proc_1_io_next_header_5),
    .io_next_header_6(proc_1_io_next_header_6),
    .io_next_header_7(proc_1_io_next_header_7),
    .io_next_header_8(proc_1_io_next_header_8),
    .io_next_header_9(proc_1_io_next_header_9),
    .io_next_header_10(proc_1_io_next_header_10),
    .io_next_header_11(proc_1_io_next_header_11),
    .io_next_header_12(proc_1_io_next_header_12),
    .io_next_header_13(proc_1_io_next_header_13),
    .io_next_header_14(proc_1_io_next_header_14),
    .io_next_header_15(proc_1_io_next_header_15),
    .io_next_header_16(proc_1_io_next_header_16),
    .io_next_header_17(proc_1_io_next_header_17),
    .io_next_header_18(proc_1_io_next_header_18),
    .io_next_header_19(proc_1_io_next_header_19),
    .io_next_header_20(proc_1_io_next_header_20),
    .io_next_header_21(proc_1_io_next_header_21),
    .io_next_header_22(proc_1_io_next_header_22),
    .io_next_header_23(proc_1_io_next_header_23),
    .io_next_header_24(proc_1_io_next_header_24),
    .io_next_header_25(proc_1_io_next_header_25),
    .io_next_header_26(proc_1_io_next_header_26),
    .io_next_header_27(proc_1_io_next_header_27),
    .io_next_header_28(proc_1_io_next_header_28),
    .io_next_header_29(proc_1_io_next_header_29),
    .io_next_header_30(proc_1_io_next_header_30),
    .io_next_header_31(proc_1_io_next_header_31),
    .io_next_header_32(proc_1_io_next_header_32),
    .io_next_header_33(proc_1_io_next_header_33),
    .io_next_header_34(proc_1_io_next_header_34),
    .io_next_header_35(proc_1_io_next_header_35),
    .io_next_header_36(proc_1_io_next_header_36),
    .io_next_header_37(proc_1_io_next_header_37),
    .io_next_header_38(proc_1_io_next_header_38),
    .io_next_header_39(proc_1_io_next_header_39),
    .io_next_header_40(proc_1_io_next_header_40),
    .io_next_header_41(proc_1_io_next_header_41),
    .io_next_header_42(proc_1_io_next_header_42),
    .io_next_header_43(proc_1_io_next_header_43),
    .io_next_header_44(proc_1_io_next_header_44),
    .io_next_header_45(proc_1_io_next_header_45),
    .io_next_header_46(proc_1_io_next_header_46),
    .io_next_header_47(proc_1_io_next_header_47),
    .io_next_header_48(proc_1_io_next_header_48),
    .io_next_header_49(proc_1_io_next_header_49),
    .io_next_header_50(proc_1_io_next_header_50),
    .io_next_header_51(proc_1_io_next_header_51),
    .io_next_header_52(proc_1_io_next_header_52),
    .io_next_header_53(proc_1_io_next_header_53),
    .io_next_header_54(proc_1_io_next_header_54),
    .io_next_header_55(proc_1_io_next_header_55),
    .io_next_header_56(proc_1_io_next_header_56),
    .io_next_header_57(proc_1_io_next_header_57),
    .io_next_header_58(proc_1_io_next_header_58),
    .io_next_header_59(proc_1_io_next_header_59),
    .io_next_header_60(proc_1_io_next_header_60),
    .io_next_header_61(proc_1_io_next_header_61),
    .io_next_header_62(proc_1_io_next_header_62),
    .io_next_header_63(proc_1_io_next_header_63),
    .io_next_proc(proc_1_io_next_proc)
  );
  ProcessorController proc_2 ( // @[controller.scala 29:25]
    .clock(proc_2_clock),
    .reset(proc_2_reset),
    .io_update(proc_2_io_update),
    .io_packet_header_0(proc_2_io_packet_header_0),
    .io_packet_header_1(proc_2_io_packet_header_1),
    .io_packet_header_2(proc_2_io_packet_header_2),
    .io_packet_header_3(proc_2_io_packet_header_3),
    .io_packet_header_4(proc_2_io_packet_header_4),
    .io_packet_header_5(proc_2_io_packet_header_5),
    .io_packet_header_6(proc_2_io_packet_header_6),
    .io_packet_header_7(proc_2_io_packet_header_7),
    .io_packet_header_8(proc_2_io_packet_header_8),
    .io_packet_header_9(proc_2_io_packet_header_9),
    .io_packet_header_10(proc_2_io_packet_header_10),
    .io_packet_header_11(proc_2_io_packet_header_11),
    .io_packet_header_12(proc_2_io_packet_header_12),
    .io_packet_header_13(proc_2_io_packet_header_13),
    .io_packet_header_14(proc_2_io_packet_header_14),
    .io_packet_header_15(proc_2_io_packet_header_15),
    .io_packet_header_16(proc_2_io_packet_header_16),
    .io_packet_header_17(proc_2_io_packet_header_17),
    .io_packet_header_18(proc_2_io_packet_header_18),
    .io_packet_header_19(proc_2_io_packet_header_19),
    .io_packet_header_20(proc_2_io_packet_header_20),
    .io_packet_header_21(proc_2_io_packet_header_21),
    .io_packet_header_22(proc_2_io_packet_header_22),
    .io_packet_header_23(proc_2_io_packet_header_23),
    .io_packet_header_24(proc_2_io_packet_header_24),
    .io_packet_header_25(proc_2_io_packet_header_25),
    .io_packet_header_26(proc_2_io_packet_header_26),
    .io_packet_header_27(proc_2_io_packet_header_27),
    .io_packet_header_28(proc_2_io_packet_header_28),
    .io_packet_header_29(proc_2_io_packet_header_29),
    .io_packet_header_30(proc_2_io_packet_header_30),
    .io_packet_header_31(proc_2_io_packet_header_31),
    .io_packet_header_32(proc_2_io_packet_header_32),
    .io_packet_header_33(proc_2_io_packet_header_33),
    .io_packet_header_34(proc_2_io_packet_header_34),
    .io_packet_header_35(proc_2_io_packet_header_35),
    .io_packet_header_36(proc_2_io_packet_header_36),
    .io_packet_header_37(proc_2_io_packet_header_37),
    .io_packet_header_38(proc_2_io_packet_header_38),
    .io_packet_header_39(proc_2_io_packet_header_39),
    .io_packet_header_40(proc_2_io_packet_header_40),
    .io_packet_header_41(proc_2_io_packet_header_41),
    .io_packet_header_42(proc_2_io_packet_header_42),
    .io_packet_header_43(proc_2_io_packet_header_43),
    .io_packet_header_44(proc_2_io_packet_header_44),
    .io_packet_header_45(proc_2_io_packet_header_45),
    .io_packet_header_46(proc_2_io_packet_header_46),
    .io_packet_header_47(proc_2_io_packet_header_47),
    .io_packet_header_48(proc_2_io_packet_header_48),
    .io_packet_header_49(proc_2_io_packet_header_49),
    .io_packet_header_50(proc_2_io_packet_header_50),
    .io_packet_header_51(proc_2_io_packet_header_51),
    .io_packet_header_52(proc_2_io_packet_header_52),
    .io_packet_header_53(proc_2_io_packet_header_53),
    .io_packet_header_54(proc_2_io_packet_header_54),
    .io_packet_header_55(proc_2_io_packet_header_55),
    .io_packet_header_56(proc_2_io_packet_header_56),
    .io_packet_header_57(proc_2_io_packet_header_57),
    .io_packet_header_58(proc_2_io_packet_header_58),
    .io_packet_header_59(proc_2_io_packet_header_59),
    .io_packet_header_60(proc_2_io_packet_header_60),
    .io_packet_header_61(proc_2_io_packet_header_61),
    .io_packet_header_62(proc_2_io_packet_header_62),
    .io_packet_header_63(proc_2_io_packet_header_63),
    .io_end(proc_2_io_end),
    .io_mem_addr(proc_2_io_mem_addr),
    .io_mem_rdata(proc_2_io_mem_rdata),
    .io_ready(proc_2_io_ready),
    .io_mod_start(proc_2_io_mod_start),
    .io_mod_hit_action_addr(proc_2_io_mod_hit_action_addr),
    .io_mod_miss_action_addr(proc_2_io_mod_miss_action_addr),
    .io_mod_ps_mod_start(proc_2_io_mod_ps_mod_start),
    .io_mod_ps_mod_header_id(proc_2_io_mod_ps_mod_header_id),
    .io_mod_ps_mod_header_length(proc_2_io_mod_ps_mod_header_length),
    .io_mod_ps_mod_next_tag_start(proc_2_io_mod_ps_mod_next_tag_start),
    .io_mod_ps_mod_next_table_0(proc_2_io_mod_ps_mod_next_table_0),
    .io_mod_ps_mod_next_table_1(proc_2_io_mod_ps_mod_next_table_1),
    .io_mod_mt_mod_start(proc_2_io_mod_mt_mod_start),
    .io_mod_mt_mod_header_id(proc_2_io_mod_mt_mod_header_id),
    .io_mod_mt_mod_key_off(proc_2_io_mod_mt_mod_key_off),
    .io_mod_mt_mod_key_len(proc_2_io_mod_mt_mod_key_len),
    .io_mod_mt_mod_val_len(proc_2_io_mod_mt_mod_val_len),
    .io_mod_ex_mod_start(proc_2_io_mod_ex_mod_start),
    .io_mod_ex_mod_ops_0(proc_2_io_mod_ex_mod_ops_0),
    .io_mod_ex_mod_ops_1(proc_2_io_mod_ex_mod_ops_1),
    .io_mod_ex_mod_ops_2(proc_2_io_mod_ex_mod_ops_2),
    .io_mod_ex_mod_ops_3(proc_2_io_mod_ex_mod_ops_3),
    .io_mod_ex_mod_ops_4(proc_2_io_mod_ex_mod_ops_4),
    .io_mod_ex_mod_ops_5(proc_2_io_mod_ex_mod_ops_5),
    .io_mod_ex_mod_ops_6(proc_2_io_mod_ex_mod_ops_6),
    .io_mod_ex_mod_ops_7(proc_2_io_mod_ex_mod_ops_7),
    .io_mod_ex_mod_ops_8(proc_2_io_mod_ex_mod_ops_8),
    .io_mod_ex_mod_ops_9(proc_2_io_mod_ex_mod_ops_9),
    .io_mod_ex_mod_ops_10(proc_2_io_mod_ex_mod_ops_10),
    .io_mod_ex_mod_ops_11(proc_2_io_mod_ex_mod_ops_11),
    .io_mod_ex_mod_ops_12(proc_2_io_mod_ex_mod_ops_12),
    .io_mod_ex_mod_ops_13(proc_2_io_mod_ex_mod_ops_13),
    .io_mod_ex_mod_ops_14(proc_2_io_mod_ex_mod_ops_14),
    .io_mod_ex_mod_ops_15(proc_2_io_mod_ex_mod_ops_15),
    .io_next_en(proc_2_io_next_en),
    .io_next_header_0(proc_2_io_next_header_0),
    .io_next_header_1(proc_2_io_next_header_1),
    .io_next_header_2(proc_2_io_next_header_2),
    .io_next_header_3(proc_2_io_next_header_3),
    .io_next_header_4(proc_2_io_next_header_4),
    .io_next_header_5(proc_2_io_next_header_5),
    .io_next_header_6(proc_2_io_next_header_6),
    .io_next_header_7(proc_2_io_next_header_7),
    .io_next_header_8(proc_2_io_next_header_8),
    .io_next_header_9(proc_2_io_next_header_9),
    .io_next_header_10(proc_2_io_next_header_10),
    .io_next_header_11(proc_2_io_next_header_11),
    .io_next_header_12(proc_2_io_next_header_12),
    .io_next_header_13(proc_2_io_next_header_13),
    .io_next_header_14(proc_2_io_next_header_14),
    .io_next_header_15(proc_2_io_next_header_15),
    .io_next_header_16(proc_2_io_next_header_16),
    .io_next_header_17(proc_2_io_next_header_17),
    .io_next_header_18(proc_2_io_next_header_18),
    .io_next_header_19(proc_2_io_next_header_19),
    .io_next_header_20(proc_2_io_next_header_20),
    .io_next_header_21(proc_2_io_next_header_21),
    .io_next_header_22(proc_2_io_next_header_22),
    .io_next_header_23(proc_2_io_next_header_23),
    .io_next_header_24(proc_2_io_next_header_24),
    .io_next_header_25(proc_2_io_next_header_25),
    .io_next_header_26(proc_2_io_next_header_26),
    .io_next_header_27(proc_2_io_next_header_27),
    .io_next_header_28(proc_2_io_next_header_28),
    .io_next_header_29(proc_2_io_next_header_29),
    .io_next_header_30(proc_2_io_next_header_30),
    .io_next_header_31(proc_2_io_next_header_31),
    .io_next_header_32(proc_2_io_next_header_32),
    .io_next_header_33(proc_2_io_next_header_33),
    .io_next_header_34(proc_2_io_next_header_34),
    .io_next_header_35(proc_2_io_next_header_35),
    .io_next_header_36(proc_2_io_next_header_36),
    .io_next_header_37(proc_2_io_next_header_37),
    .io_next_header_38(proc_2_io_next_header_38),
    .io_next_header_39(proc_2_io_next_header_39),
    .io_next_header_40(proc_2_io_next_header_40),
    .io_next_header_41(proc_2_io_next_header_41),
    .io_next_header_42(proc_2_io_next_header_42),
    .io_next_header_43(proc_2_io_next_header_43),
    .io_next_header_44(proc_2_io_next_header_44),
    .io_next_header_45(proc_2_io_next_header_45),
    .io_next_header_46(proc_2_io_next_header_46),
    .io_next_header_47(proc_2_io_next_header_47),
    .io_next_header_48(proc_2_io_next_header_48),
    .io_next_header_49(proc_2_io_next_header_49),
    .io_next_header_50(proc_2_io_next_header_50),
    .io_next_header_51(proc_2_io_next_header_51),
    .io_next_header_52(proc_2_io_next_header_52),
    .io_next_header_53(proc_2_io_next_header_53),
    .io_next_header_54(proc_2_io_next_header_54),
    .io_next_header_55(proc_2_io_next_header_55),
    .io_next_header_56(proc_2_io_next_header_56),
    .io_next_header_57(proc_2_io_next_header_57),
    .io_next_header_58(proc_2_io_next_header_58),
    .io_next_header_59(proc_2_io_next_header_59),
    .io_next_header_60(proc_2_io_next_header_60),
    .io_next_header_61(proc_2_io_next_header_61),
    .io_next_header_62(proc_2_io_next_header_62),
    .io_next_header_63(proc_2_io_next_header_63),
    .io_next_proc(proc_2_io_next_proc)
  );
  ProcessorController proc_3 ( // @[controller.scala 29:25]
    .clock(proc_3_clock),
    .reset(proc_3_reset),
    .io_update(proc_3_io_update),
    .io_packet_header_0(proc_3_io_packet_header_0),
    .io_packet_header_1(proc_3_io_packet_header_1),
    .io_packet_header_2(proc_3_io_packet_header_2),
    .io_packet_header_3(proc_3_io_packet_header_3),
    .io_packet_header_4(proc_3_io_packet_header_4),
    .io_packet_header_5(proc_3_io_packet_header_5),
    .io_packet_header_6(proc_3_io_packet_header_6),
    .io_packet_header_7(proc_3_io_packet_header_7),
    .io_packet_header_8(proc_3_io_packet_header_8),
    .io_packet_header_9(proc_3_io_packet_header_9),
    .io_packet_header_10(proc_3_io_packet_header_10),
    .io_packet_header_11(proc_3_io_packet_header_11),
    .io_packet_header_12(proc_3_io_packet_header_12),
    .io_packet_header_13(proc_3_io_packet_header_13),
    .io_packet_header_14(proc_3_io_packet_header_14),
    .io_packet_header_15(proc_3_io_packet_header_15),
    .io_packet_header_16(proc_3_io_packet_header_16),
    .io_packet_header_17(proc_3_io_packet_header_17),
    .io_packet_header_18(proc_3_io_packet_header_18),
    .io_packet_header_19(proc_3_io_packet_header_19),
    .io_packet_header_20(proc_3_io_packet_header_20),
    .io_packet_header_21(proc_3_io_packet_header_21),
    .io_packet_header_22(proc_3_io_packet_header_22),
    .io_packet_header_23(proc_3_io_packet_header_23),
    .io_packet_header_24(proc_3_io_packet_header_24),
    .io_packet_header_25(proc_3_io_packet_header_25),
    .io_packet_header_26(proc_3_io_packet_header_26),
    .io_packet_header_27(proc_3_io_packet_header_27),
    .io_packet_header_28(proc_3_io_packet_header_28),
    .io_packet_header_29(proc_3_io_packet_header_29),
    .io_packet_header_30(proc_3_io_packet_header_30),
    .io_packet_header_31(proc_3_io_packet_header_31),
    .io_packet_header_32(proc_3_io_packet_header_32),
    .io_packet_header_33(proc_3_io_packet_header_33),
    .io_packet_header_34(proc_3_io_packet_header_34),
    .io_packet_header_35(proc_3_io_packet_header_35),
    .io_packet_header_36(proc_3_io_packet_header_36),
    .io_packet_header_37(proc_3_io_packet_header_37),
    .io_packet_header_38(proc_3_io_packet_header_38),
    .io_packet_header_39(proc_3_io_packet_header_39),
    .io_packet_header_40(proc_3_io_packet_header_40),
    .io_packet_header_41(proc_3_io_packet_header_41),
    .io_packet_header_42(proc_3_io_packet_header_42),
    .io_packet_header_43(proc_3_io_packet_header_43),
    .io_packet_header_44(proc_3_io_packet_header_44),
    .io_packet_header_45(proc_3_io_packet_header_45),
    .io_packet_header_46(proc_3_io_packet_header_46),
    .io_packet_header_47(proc_3_io_packet_header_47),
    .io_packet_header_48(proc_3_io_packet_header_48),
    .io_packet_header_49(proc_3_io_packet_header_49),
    .io_packet_header_50(proc_3_io_packet_header_50),
    .io_packet_header_51(proc_3_io_packet_header_51),
    .io_packet_header_52(proc_3_io_packet_header_52),
    .io_packet_header_53(proc_3_io_packet_header_53),
    .io_packet_header_54(proc_3_io_packet_header_54),
    .io_packet_header_55(proc_3_io_packet_header_55),
    .io_packet_header_56(proc_3_io_packet_header_56),
    .io_packet_header_57(proc_3_io_packet_header_57),
    .io_packet_header_58(proc_3_io_packet_header_58),
    .io_packet_header_59(proc_3_io_packet_header_59),
    .io_packet_header_60(proc_3_io_packet_header_60),
    .io_packet_header_61(proc_3_io_packet_header_61),
    .io_packet_header_62(proc_3_io_packet_header_62),
    .io_packet_header_63(proc_3_io_packet_header_63),
    .io_end(proc_3_io_end),
    .io_mem_addr(proc_3_io_mem_addr),
    .io_mem_rdata(proc_3_io_mem_rdata),
    .io_ready(proc_3_io_ready),
    .io_mod_start(proc_3_io_mod_start),
    .io_mod_hit_action_addr(proc_3_io_mod_hit_action_addr),
    .io_mod_miss_action_addr(proc_3_io_mod_miss_action_addr),
    .io_mod_ps_mod_start(proc_3_io_mod_ps_mod_start),
    .io_mod_ps_mod_header_id(proc_3_io_mod_ps_mod_header_id),
    .io_mod_ps_mod_header_length(proc_3_io_mod_ps_mod_header_length),
    .io_mod_ps_mod_next_tag_start(proc_3_io_mod_ps_mod_next_tag_start),
    .io_mod_ps_mod_next_table_0(proc_3_io_mod_ps_mod_next_table_0),
    .io_mod_ps_mod_next_table_1(proc_3_io_mod_ps_mod_next_table_1),
    .io_mod_mt_mod_start(proc_3_io_mod_mt_mod_start),
    .io_mod_mt_mod_header_id(proc_3_io_mod_mt_mod_header_id),
    .io_mod_mt_mod_key_off(proc_3_io_mod_mt_mod_key_off),
    .io_mod_mt_mod_key_len(proc_3_io_mod_mt_mod_key_len),
    .io_mod_mt_mod_val_len(proc_3_io_mod_mt_mod_val_len),
    .io_mod_ex_mod_start(proc_3_io_mod_ex_mod_start),
    .io_mod_ex_mod_ops_0(proc_3_io_mod_ex_mod_ops_0),
    .io_mod_ex_mod_ops_1(proc_3_io_mod_ex_mod_ops_1),
    .io_mod_ex_mod_ops_2(proc_3_io_mod_ex_mod_ops_2),
    .io_mod_ex_mod_ops_3(proc_3_io_mod_ex_mod_ops_3),
    .io_mod_ex_mod_ops_4(proc_3_io_mod_ex_mod_ops_4),
    .io_mod_ex_mod_ops_5(proc_3_io_mod_ex_mod_ops_5),
    .io_mod_ex_mod_ops_6(proc_3_io_mod_ex_mod_ops_6),
    .io_mod_ex_mod_ops_7(proc_3_io_mod_ex_mod_ops_7),
    .io_mod_ex_mod_ops_8(proc_3_io_mod_ex_mod_ops_8),
    .io_mod_ex_mod_ops_9(proc_3_io_mod_ex_mod_ops_9),
    .io_mod_ex_mod_ops_10(proc_3_io_mod_ex_mod_ops_10),
    .io_mod_ex_mod_ops_11(proc_3_io_mod_ex_mod_ops_11),
    .io_mod_ex_mod_ops_12(proc_3_io_mod_ex_mod_ops_12),
    .io_mod_ex_mod_ops_13(proc_3_io_mod_ex_mod_ops_13),
    .io_mod_ex_mod_ops_14(proc_3_io_mod_ex_mod_ops_14),
    .io_mod_ex_mod_ops_15(proc_3_io_mod_ex_mod_ops_15),
    .io_next_en(proc_3_io_next_en),
    .io_next_header_0(proc_3_io_next_header_0),
    .io_next_header_1(proc_3_io_next_header_1),
    .io_next_header_2(proc_3_io_next_header_2),
    .io_next_header_3(proc_3_io_next_header_3),
    .io_next_header_4(proc_3_io_next_header_4),
    .io_next_header_5(proc_3_io_next_header_5),
    .io_next_header_6(proc_3_io_next_header_6),
    .io_next_header_7(proc_3_io_next_header_7),
    .io_next_header_8(proc_3_io_next_header_8),
    .io_next_header_9(proc_3_io_next_header_9),
    .io_next_header_10(proc_3_io_next_header_10),
    .io_next_header_11(proc_3_io_next_header_11),
    .io_next_header_12(proc_3_io_next_header_12),
    .io_next_header_13(proc_3_io_next_header_13),
    .io_next_header_14(proc_3_io_next_header_14),
    .io_next_header_15(proc_3_io_next_header_15),
    .io_next_header_16(proc_3_io_next_header_16),
    .io_next_header_17(proc_3_io_next_header_17),
    .io_next_header_18(proc_3_io_next_header_18),
    .io_next_header_19(proc_3_io_next_header_19),
    .io_next_header_20(proc_3_io_next_header_20),
    .io_next_header_21(proc_3_io_next_header_21),
    .io_next_header_22(proc_3_io_next_header_22),
    .io_next_header_23(proc_3_io_next_header_23),
    .io_next_header_24(proc_3_io_next_header_24),
    .io_next_header_25(proc_3_io_next_header_25),
    .io_next_header_26(proc_3_io_next_header_26),
    .io_next_header_27(proc_3_io_next_header_27),
    .io_next_header_28(proc_3_io_next_header_28),
    .io_next_header_29(proc_3_io_next_header_29),
    .io_next_header_30(proc_3_io_next_header_30),
    .io_next_header_31(proc_3_io_next_header_31),
    .io_next_header_32(proc_3_io_next_header_32),
    .io_next_header_33(proc_3_io_next_header_33),
    .io_next_header_34(proc_3_io_next_header_34),
    .io_next_header_35(proc_3_io_next_header_35),
    .io_next_header_36(proc_3_io_next_header_36),
    .io_next_header_37(proc_3_io_next_header_37),
    .io_next_header_38(proc_3_io_next_header_38),
    .io_next_header_39(proc_3_io_next_header_39),
    .io_next_header_40(proc_3_io_next_header_40),
    .io_next_header_41(proc_3_io_next_header_41),
    .io_next_header_42(proc_3_io_next_header_42),
    .io_next_header_43(proc_3_io_next_header_43),
    .io_next_header_44(proc_3_io_next_header_44),
    .io_next_header_45(proc_3_io_next_header_45),
    .io_next_header_46(proc_3_io_next_header_46),
    .io_next_header_47(proc_3_io_next_header_47),
    .io_next_header_48(proc_3_io_next_header_48),
    .io_next_header_49(proc_3_io_next_header_49),
    .io_next_header_50(proc_3_io_next_header_50),
    .io_next_header_51(proc_3_io_next_header_51),
    .io_next_header_52(proc_3_io_next_header_52),
    .io_next_header_53(proc_3_io_next_header_53),
    .io_next_header_54(proc_3_io_next_header_54),
    .io_next_header_55(proc_3_io_next_header_55),
    .io_next_header_56(proc_3_io_next_header_56),
    .io_next_header_57(proc_3_io_next_header_57),
    .io_next_header_58(proc_3_io_next_header_58),
    .io_next_header_59(proc_3_io_next_header_59),
    .io_next_header_60(proc_3_io_next_header_60),
    .io_next_header_61(proc_3_io_next_header_61),
    .io_next_header_62(proc_3_io_next_header_62),
    .io_next_header_63(proc_3_io_next_header_63),
    .io_next_proc(proc_3_io_next_proc)
  );
  ProcessorController proc_4 ( // @[controller.scala 29:25]
    .clock(proc_4_clock),
    .reset(proc_4_reset),
    .io_update(proc_4_io_update),
    .io_packet_header_0(proc_4_io_packet_header_0),
    .io_packet_header_1(proc_4_io_packet_header_1),
    .io_packet_header_2(proc_4_io_packet_header_2),
    .io_packet_header_3(proc_4_io_packet_header_3),
    .io_packet_header_4(proc_4_io_packet_header_4),
    .io_packet_header_5(proc_4_io_packet_header_5),
    .io_packet_header_6(proc_4_io_packet_header_6),
    .io_packet_header_7(proc_4_io_packet_header_7),
    .io_packet_header_8(proc_4_io_packet_header_8),
    .io_packet_header_9(proc_4_io_packet_header_9),
    .io_packet_header_10(proc_4_io_packet_header_10),
    .io_packet_header_11(proc_4_io_packet_header_11),
    .io_packet_header_12(proc_4_io_packet_header_12),
    .io_packet_header_13(proc_4_io_packet_header_13),
    .io_packet_header_14(proc_4_io_packet_header_14),
    .io_packet_header_15(proc_4_io_packet_header_15),
    .io_packet_header_16(proc_4_io_packet_header_16),
    .io_packet_header_17(proc_4_io_packet_header_17),
    .io_packet_header_18(proc_4_io_packet_header_18),
    .io_packet_header_19(proc_4_io_packet_header_19),
    .io_packet_header_20(proc_4_io_packet_header_20),
    .io_packet_header_21(proc_4_io_packet_header_21),
    .io_packet_header_22(proc_4_io_packet_header_22),
    .io_packet_header_23(proc_4_io_packet_header_23),
    .io_packet_header_24(proc_4_io_packet_header_24),
    .io_packet_header_25(proc_4_io_packet_header_25),
    .io_packet_header_26(proc_4_io_packet_header_26),
    .io_packet_header_27(proc_4_io_packet_header_27),
    .io_packet_header_28(proc_4_io_packet_header_28),
    .io_packet_header_29(proc_4_io_packet_header_29),
    .io_packet_header_30(proc_4_io_packet_header_30),
    .io_packet_header_31(proc_4_io_packet_header_31),
    .io_packet_header_32(proc_4_io_packet_header_32),
    .io_packet_header_33(proc_4_io_packet_header_33),
    .io_packet_header_34(proc_4_io_packet_header_34),
    .io_packet_header_35(proc_4_io_packet_header_35),
    .io_packet_header_36(proc_4_io_packet_header_36),
    .io_packet_header_37(proc_4_io_packet_header_37),
    .io_packet_header_38(proc_4_io_packet_header_38),
    .io_packet_header_39(proc_4_io_packet_header_39),
    .io_packet_header_40(proc_4_io_packet_header_40),
    .io_packet_header_41(proc_4_io_packet_header_41),
    .io_packet_header_42(proc_4_io_packet_header_42),
    .io_packet_header_43(proc_4_io_packet_header_43),
    .io_packet_header_44(proc_4_io_packet_header_44),
    .io_packet_header_45(proc_4_io_packet_header_45),
    .io_packet_header_46(proc_4_io_packet_header_46),
    .io_packet_header_47(proc_4_io_packet_header_47),
    .io_packet_header_48(proc_4_io_packet_header_48),
    .io_packet_header_49(proc_4_io_packet_header_49),
    .io_packet_header_50(proc_4_io_packet_header_50),
    .io_packet_header_51(proc_4_io_packet_header_51),
    .io_packet_header_52(proc_4_io_packet_header_52),
    .io_packet_header_53(proc_4_io_packet_header_53),
    .io_packet_header_54(proc_4_io_packet_header_54),
    .io_packet_header_55(proc_4_io_packet_header_55),
    .io_packet_header_56(proc_4_io_packet_header_56),
    .io_packet_header_57(proc_4_io_packet_header_57),
    .io_packet_header_58(proc_4_io_packet_header_58),
    .io_packet_header_59(proc_4_io_packet_header_59),
    .io_packet_header_60(proc_4_io_packet_header_60),
    .io_packet_header_61(proc_4_io_packet_header_61),
    .io_packet_header_62(proc_4_io_packet_header_62),
    .io_packet_header_63(proc_4_io_packet_header_63),
    .io_end(proc_4_io_end),
    .io_mem_addr(proc_4_io_mem_addr),
    .io_mem_rdata(proc_4_io_mem_rdata),
    .io_ready(proc_4_io_ready),
    .io_mod_start(proc_4_io_mod_start),
    .io_mod_hit_action_addr(proc_4_io_mod_hit_action_addr),
    .io_mod_miss_action_addr(proc_4_io_mod_miss_action_addr),
    .io_mod_ps_mod_start(proc_4_io_mod_ps_mod_start),
    .io_mod_ps_mod_header_id(proc_4_io_mod_ps_mod_header_id),
    .io_mod_ps_mod_header_length(proc_4_io_mod_ps_mod_header_length),
    .io_mod_ps_mod_next_tag_start(proc_4_io_mod_ps_mod_next_tag_start),
    .io_mod_ps_mod_next_table_0(proc_4_io_mod_ps_mod_next_table_0),
    .io_mod_ps_mod_next_table_1(proc_4_io_mod_ps_mod_next_table_1),
    .io_mod_mt_mod_start(proc_4_io_mod_mt_mod_start),
    .io_mod_mt_mod_header_id(proc_4_io_mod_mt_mod_header_id),
    .io_mod_mt_mod_key_off(proc_4_io_mod_mt_mod_key_off),
    .io_mod_mt_mod_key_len(proc_4_io_mod_mt_mod_key_len),
    .io_mod_mt_mod_val_len(proc_4_io_mod_mt_mod_val_len),
    .io_mod_ex_mod_start(proc_4_io_mod_ex_mod_start),
    .io_mod_ex_mod_ops_0(proc_4_io_mod_ex_mod_ops_0),
    .io_mod_ex_mod_ops_1(proc_4_io_mod_ex_mod_ops_1),
    .io_mod_ex_mod_ops_2(proc_4_io_mod_ex_mod_ops_2),
    .io_mod_ex_mod_ops_3(proc_4_io_mod_ex_mod_ops_3),
    .io_mod_ex_mod_ops_4(proc_4_io_mod_ex_mod_ops_4),
    .io_mod_ex_mod_ops_5(proc_4_io_mod_ex_mod_ops_5),
    .io_mod_ex_mod_ops_6(proc_4_io_mod_ex_mod_ops_6),
    .io_mod_ex_mod_ops_7(proc_4_io_mod_ex_mod_ops_7),
    .io_mod_ex_mod_ops_8(proc_4_io_mod_ex_mod_ops_8),
    .io_mod_ex_mod_ops_9(proc_4_io_mod_ex_mod_ops_9),
    .io_mod_ex_mod_ops_10(proc_4_io_mod_ex_mod_ops_10),
    .io_mod_ex_mod_ops_11(proc_4_io_mod_ex_mod_ops_11),
    .io_mod_ex_mod_ops_12(proc_4_io_mod_ex_mod_ops_12),
    .io_mod_ex_mod_ops_13(proc_4_io_mod_ex_mod_ops_13),
    .io_mod_ex_mod_ops_14(proc_4_io_mod_ex_mod_ops_14),
    .io_mod_ex_mod_ops_15(proc_4_io_mod_ex_mod_ops_15),
    .io_next_en(proc_4_io_next_en),
    .io_next_header_0(proc_4_io_next_header_0),
    .io_next_header_1(proc_4_io_next_header_1),
    .io_next_header_2(proc_4_io_next_header_2),
    .io_next_header_3(proc_4_io_next_header_3),
    .io_next_header_4(proc_4_io_next_header_4),
    .io_next_header_5(proc_4_io_next_header_5),
    .io_next_header_6(proc_4_io_next_header_6),
    .io_next_header_7(proc_4_io_next_header_7),
    .io_next_header_8(proc_4_io_next_header_8),
    .io_next_header_9(proc_4_io_next_header_9),
    .io_next_header_10(proc_4_io_next_header_10),
    .io_next_header_11(proc_4_io_next_header_11),
    .io_next_header_12(proc_4_io_next_header_12),
    .io_next_header_13(proc_4_io_next_header_13),
    .io_next_header_14(proc_4_io_next_header_14),
    .io_next_header_15(proc_4_io_next_header_15),
    .io_next_header_16(proc_4_io_next_header_16),
    .io_next_header_17(proc_4_io_next_header_17),
    .io_next_header_18(proc_4_io_next_header_18),
    .io_next_header_19(proc_4_io_next_header_19),
    .io_next_header_20(proc_4_io_next_header_20),
    .io_next_header_21(proc_4_io_next_header_21),
    .io_next_header_22(proc_4_io_next_header_22),
    .io_next_header_23(proc_4_io_next_header_23),
    .io_next_header_24(proc_4_io_next_header_24),
    .io_next_header_25(proc_4_io_next_header_25),
    .io_next_header_26(proc_4_io_next_header_26),
    .io_next_header_27(proc_4_io_next_header_27),
    .io_next_header_28(proc_4_io_next_header_28),
    .io_next_header_29(proc_4_io_next_header_29),
    .io_next_header_30(proc_4_io_next_header_30),
    .io_next_header_31(proc_4_io_next_header_31),
    .io_next_header_32(proc_4_io_next_header_32),
    .io_next_header_33(proc_4_io_next_header_33),
    .io_next_header_34(proc_4_io_next_header_34),
    .io_next_header_35(proc_4_io_next_header_35),
    .io_next_header_36(proc_4_io_next_header_36),
    .io_next_header_37(proc_4_io_next_header_37),
    .io_next_header_38(proc_4_io_next_header_38),
    .io_next_header_39(proc_4_io_next_header_39),
    .io_next_header_40(proc_4_io_next_header_40),
    .io_next_header_41(proc_4_io_next_header_41),
    .io_next_header_42(proc_4_io_next_header_42),
    .io_next_header_43(proc_4_io_next_header_43),
    .io_next_header_44(proc_4_io_next_header_44),
    .io_next_header_45(proc_4_io_next_header_45),
    .io_next_header_46(proc_4_io_next_header_46),
    .io_next_header_47(proc_4_io_next_header_47),
    .io_next_header_48(proc_4_io_next_header_48),
    .io_next_header_49(proc_4_io_next_header_49),
    .io_next_header_50(proc_4_io_next_header_50),
    .io_next_header_51(proc_4_io_next_header_51),
    .io_next_header_52(proc_4_io_next_header_52),
    .io_next_header_53(proc_4_io_next_header_53),
    .io_next_header_54(proc_4_io_next_header_54),
    .io_next_header_55(proc_4_io_next_header_55),
    .io_next_header_56(proc_4_io_next_header_56),
    .io_next_header_57(proc_4_io_next_header_57),
    .io_next_header_58(proc_4_io_next_header_58),
    .io_next_header_59(proc_4_io_next_header_59),
    .io_next_header_60(proc_4_io_next_header_60),
    .io_next_header_61(proc_4_io_next_header_61),
    .io_next_header_62(proc_4_io_next_header_62),
    .io_next_header_63(proc_4_io_next_header_63),
    .io_next_proc(proc_4_io_next_proc)
  );
  ProcessorController proc_5 ( // @[controller.scala 29:25]
    .clock(proc_5_clock),
    .reset(proc_5_reset),
    .io_update(proc_5_io_update),
    .io_packet_header_0(proc_5_io_packet_header_0),
    .io_packet_header_1(proc_5_io_packet_header_1),
    .io_packet_header_2(proc_5_io_packet_header_2),
    .io_packet_header_3(proc_5_io_packet_header_3),
    .io_packet_header_4(proc_5_io_packet_header_4),
    .io_packet_header_5(proc_5_io_packet_header_5),
    .io_packet_header_6(proc_5_io_packet_header_6),
    .io_packet_header_7(proc_5_io_packet_header_7),
    .io_packet_header_8(proc_5_io_packet_header_8),
    .io_packet_header_9(proc_5_io_packet_header_9),
    .io_packet_header_10(proc_5_io_packet_header_10),
    .io_packet_header_11(proc_5_io_packet_header_11),
    .io_packet_header_12(proc_5_io_packet_header_12),
    .io_packet_header_13(proc_5_io_packet_header_13),
    .io_packet_header_14(proc_5_io_packet_header_14),
    .io_packet_header_15(proc_5_io_packet_header_15),
    .io_packet_header_16(proc_5_io_packet_header_16),
    .io_packet_header_17(proc_5_io_packet_header_17),
    .io_packet_header_18(proc_5_io_packet_header_18),
    .io_packet_header_19(proc_5_io_packet_header_19),
    .io_packet_header_20(proc_5_io_packet_header_20),
    .io_packet_header_21(proc_5_io_packet_header_21),
    .io_packet_header_22(proc_5_io_packet_header_22),
    .io_packet_header_23(proc_5_io_packet_header_23),
    .io_packet_header_24(proc_5_io_packet_header_24),
    .io_packet_header_25(proc_5_io_packet_header_25),
    .io_packet_header_26(proc_5_io_packet_header_26),
    .io_packet_header_27(proc_5_io_packet_header_27),
    .io_packet_header_28(proc_5_io_packet_header_28),
    .io_packet_header_29(proc_5_io_packet_header_29),
    .io_packet_header_30(proc_5_io_packet_header_30),
    .io_packet_header_31(proc_5_io_packet_header_31),
    .io_packet_header_32(proc_5_io_packet_header_32),
    .io_packet_header_33(proc_5_io_packet_header_33),
    .io_packet_header_34(proc_5_io_packet_header_34),
    .io_packet_header_35(proc_5_io_packet_header_35),
    .io_packet_header_36(proc_5_io_packet_header_36),
    .io_packet_header_37(proc_5_io_packet_header_37),
    .io_packet_header_38(proc_5_io_packet_header_38),
    .io_packet_header_39(proc_5_io_packet_header_39),
    .io_packet_header_40(proc_5_io_packet_header_40),
    .io_packet_header_41(proc_5_io_packet_header_41),
    .io_packet_header_42(proc_5_io_packet_header_42),
    .io_packet_header_43(proc_5_io_packet_header_43),
    .io_packet_header_44(proc_5_io_packet_header_44),
    .io_packet_header_45(proc_5_io_packet_header_45),
    .io_packet_header_46(proc_5_io_packet_header_46),
    .io_packet_header_47(proc_5_io_packet_header_47),
    .io_packet_header_48(proc_5_io_packet_header_48),
    .io_packet_header_49(proc_5_io_packet_header_49),
    .io_packet_header_50(proc_5_io_packet_header_50),
    .io_packet_header_51(proc_5_io_packet_header_51),
    .io_packet_header_52(proc_5_io_packet_header_52),
    .io_packet_header_53(proc_5_io_packet_header_53),
    .io_packet_header_54(proc_5_io_packet_header_54),
    .io_packet_header_55(proc_5_io_packet_header_55),
    .io_packet_header_56(proc_5_io_packet_header_56),
    .io_packet_header_57(proc_5_io_packet_header_57),
    .io_packet_header_58(proc_5_io_packet_header_58),
    .io_packet_header_59(proc_5_io_packet_header_59),
    .io_packet_header_60(proc_5_io_packet_header_60),
    .io_packet_header_61(proc_5_io_packet_header_61),
    .io_packet_header_62(proc_5_io_packet_header_62),
    .io_packet_header_63(proc_5_io_packet_header_63),
    .io_end(proc_5_io_end),
    .io_mem_addr(proc_5_io_mem_addr),
    .io_mem_rdata(proc_5_io_mem_rdata),
    .io_ready(proc_5_io_ready),
    .io_mod_start(proc_5_io_mod_start),
    .io_mod_hit_action_addr(proc_5_io_mod_hit_action_addr),
    .io_mod_miss_action_addr(proc_5_io_mod_miss_action_addr),
    .io_mod_ps_mod_start(proc_5_io_mod_ps_mod_start),
    .io_mod_ps_mod_header_id(proc_5_io_mod_ps_mod_header_id),
    .io_mod_ps_mod_header_length(proc_5_io_mod_ps_mod_header_length),
    .io_mod_ps_mod_next_tag_start(proc_5_io_mod_ps_mod_next_tag_start),
    .io_mod_ps_mod_next_table_0(proc_5_io_mod_ps_mod_next_table_0),
    .io_mod_ps_mod_next_table_1(proc_5_io_mod_ps_mod_next_table_1),
    .io_mod_mt_mod_start(proc_5_io_mod_mt_mod_start),
    .io_mod_mt_mod_header_id(proc_5_io_mod_mt_mod_header_id),
    .io_mod_mt_mod_key_off(proc_5_io_mod_mt_mod_key_off),
    .io_mod_mt_mod_key_len(proc_5_io_mod_mt_mod_key_len),
    .io_mod_mt_mod_val_len(proc_5_io_mod_mt_mod_val_len),
    .io_mod_ex_mod_start(proc_5_io_mod_ex_mod_start),
    .io_mod_ex_mod_ops_0(proc_5_io_mod_ex_mod_ops_0),
    .io_mod_ex_mod_ops_1(proc_5_io_mod_ex_mod_ops_1),
    .io_mod_ex_mod_ops_2(proc_5_io_mod_ex_mod_ops_2),
    .io_mod_ex_mod_ops_3(proc_5_io_mod_ex_mod_ops_3),
    .io_mod_ex_mod_ops_4(proc_5_io_mod_ex_mod_ops_4),
    .io_mod_ex_mod_ops_5(proc_5_io_mod_ex_mod_ops_5),
    .io_mod_ex_mod_ops_6(proc_5_io_mod_ex_mod_ops_6),
    .io_mod_ex_mod_ops_7(proc_5_io_mod_ex_mod_ops_7),
    .io_mod_ex_mod_ops_8(proc_5_io_mod_ex_mod_ops_8),
    .io_mod_ex_mod_ops_9(proc_5_io_mod_ex_mod_ops_9),
    .io_mod_ex_mod_ops_10(proc_5_io_mod_ex_mod_ops_10),
    .io_mod_ex_mod_ops_11(proc_5_io_mod_ex_mod_ops_11),
    .io_mod_ex_mod_ops_12(proc_5_io_mod_ex_mod_ops_12),
    .io_mod_ex_mod_ops_13(proc_5_io_mod_ex_mod_ops_13),
    .io_mod_ex_mod_ops_14(proc_5_io_mod_ex_mod_ops_14),
    .io_mod_ex_mod_ops_15(proc_5_io_mod_ex_mod_ops_15),
    .io_next_en(proc_5_io_next_en),
    .io_next_header_0(proc_5_io_next_header_0),
    .io_next_header_1(proc_5_io_next_header_1),
    .io_next_header_2(proc_5_io_next_header_2),
    .io_next_header_3(proc_5_io_next_header_3),
    .io_next_header_4(proc_5_io_next_header_4),
    .io_next_header_5(proc_5_io_next_header_5),
    .io_next_header_6(proc_5_io_next_header_6),
    .io_next_header_7(proc_5_io_next_header_7),
    .io_next_header_8(proc_5_io_next_header_8),
    .io_next_header_9(proc_5_io_next_header_9),
    .io_next_header_10(proc_5_io_next_header_10),
    .io_next_header_11(proc_5_io_next_header_11),
    .io_next_header_12(proc_5_io_next_header_12),
    .io_next_header_13(proc_5_io_next_header_13),
    .io_next_header_14(proc_5_io_next_header_14),
    .io_next_header_15(proc_5_io_next_header_15),
    .io_next_header_16(proc_5_io_next_header_16),
    .io_next_header_17(proc_5_io_next_header_17),
    .io_next_header_18(proc_5_io_next_header_18),
    .io_next_header_19(proc_5_io_next_header_19),
    .io_next_header_20(proc_5_io_next_header_20),
    .io_next_header_21(proc_5_io_next_header_21),
    .io_next_header_22(proc_5_io_next_header_22),
    .io_next_header_23(proc_5_io_next_header_23),
    .io_next_header_24(proc_5_io_next_header_24),
    .io_next_header_25(proc_5_io_next_header_25),
    .io_next_header_26(proc_5_io_next_header_26),
    .io_next_header_27(proc_5_io_next_header_27),
    .io_next_header_28(proc_5_io_next_header_28),
    .io_next_header_29(proc_5_io_next_header_29),
    .io_next_header_30(proc_5_io_next_header_30),
    .io_next_header_31(proc_5_io_next_header_31),
    .io_next_header_32(proc_5_io_next_header_32),
    .io_next_header_33(proc_5_io_next_header_33),
    .io_next_header_34(proc_5_io_next_header_34),
    .io_next_header_35(proc_5_io_next_header_35),
    .io_next_header_36(proc_5_io_next_header_36),
    .io_next_header_37(proc_5_io_next_header_37),
    .io_next_header_38(proc_5_io_next_header_38),
    .io_next_header_39(proc_5_io_next_header_39),
    .io_next_header_40(proc_5_io_next_header_40),
    .io_next_header_41(proc_5_io_next_header_41),
    .io_next_header_42(proc_5_io_next_header_42),
    .io_next_header_43(proc_5_io_next_header_43),
    .io_next_header_44(proc_5_io_next_header_44),
    .io_next_header_45(proc_5_io_next_header_45),
    .io_next_header_46(proc_5_io_next_header_46),
    .io_next_header_47(proc_5_io_next_header_47),
    .io_next_header_48(proc_5_io_next_header_48),
    .io_next_header_49(proc_5_io_next_header_49),
    .io_next_header_50(proc_5_io_next_header_50),
    .io_next_header_51(proc_5_io_next_header_51),
    .io_next_header_52(proc_5_io_next_header_52),
    .io_next_header_53(proc_5_io_next_header_53),
    .io_next_header_54(proc_5_io_next_header_54),
    .io_next_header_55(proc_5_io_next_header_55),
    .io_next_header_56(proc_5_io_next_header_56),
    .io_next_header_57(proc_5_io_next_header_57),
    .io_next_header_58(proc_5_io_next_header_58),
    .io_next_header_59(proc_5_io_next_header_59),
    .io_next_header_60(proc_5_io_next_header_60),
    .io_next_header_61(proc_5_io_next_header_61),
    .io_next_header_62(proc_5_io_next_header_62),
    .io_next_header_63(proc_5_io_next_header_63),
    .io_next_proc(proc_5_io_next_proc)
  );
  ProcessorController proc_6 ( // @[controller.scala 29:25]
    .clock(proc_6_clock),
    .reset(proc_6_reset),
    .io_update(proc_6_io_update),
    .io_packet_header_0(proc_6_io_packet_header_0),
    .io_packet_header_1(proc_6_io_packet_header_1),
    .io_packet_header_2(proc_6_io_packet_header_2),
    .io_packet_header_3(proc_6_io_packet_header_3),
    .io_packet_header_4(proc_6_io_packet_header_4),
    .io_packet_header_5(proc_6_io_packet_header_5),
    .io_packet_header_6(proc_6_io_packet_header_6),
    .io_packet_header_7(proc_6_io_packet_header_7),
    .io_packet_header_8(proc_6_io_packet_header_8),
    .io_packet_header_9(proc_6_io_packet_header_9),
    .io_packet_header_10(proc_6_io_packet_header_10),
    .io_packet_header_11(proc_6_io_packet_header_11),
    .io_packet_header_12(proc_6_io_packet_header_12),
    .io_packet_header_13(proc_6_io_packet_header_13),
    .io_packet_header_14(proc_6_io_packet_header_14),
    .io_packet_header_15(proc_6_io_packet_header_15),
    .io_packet_header_16(proc_6_io_packet_header_16),
    .io_packet_header_17(proc_6_io_packet_header_17),
    .io_packet_header_18(proc_6_io_packet_header_18),
    .io_packet_header_19(proc_6_io_packet_header_19),
    .io_packet_header_20(proc_6_io_packet_header_20),
    .io_packet_header_21(proc_6_io_packet_header_21),
    .io_packet_header_22(proc_6_io_packet_header_22),
    .io_packet_header_23(proc_6_io_packet_header_23),
    .io_packet_header_24(proc_6_io_packet_header_24),
    .io_packet_header_25(proc_6_io_packet_header_25),
    .io_packet_header_26(proc_6_io_packet_header_26),
    .io_packet_header_27(proc_6_io_packet_header_27),
    .io_packet_header_28(proc_6_io_packet_header_28),
    .io_packet_header_29(proc_6_io_packet_header_29),
    .io_packet_header_30(proc_6_io_packet_header_30),
    .io_packet_header_31(proc_6_io_packet_header_31),
    .io_packet_header_32(proc_6_io_packet_header_32),
    .io_packet_header_33(proc_6_io_packet_header_33),
    .io_packet_header_34(proc_6_io_packet_header_34),
    .io_packet_header_35(proc_6_io_packet_header_35),
    .io_packet_header_36(proc_6_io_packet_header_36),
    .io_packet_header_37(proc_6_io_packet_header_37),
    .io_packet_header_38(proc_6_io_packet_header_38),
    .io_packet_header_39(proc_6_io_packet_header_39),
    .io_packet_header_40(proc_6_io_packet_header_40),
    .io_packet_header_41(proc_6_io_packet_header_41),
    .io_packet_header_42(proc_6_io_packet_header_42),
    .io_packet_header_43(proc_6_io_packet_header_43),
    .io_packet_header_44(proc_6_io_packet_header_44),
    .io_packet_header_45(proc_6_io_packet_header_45),
    .io_packet_header_46(proc_6_io_packet_header_46),
    .io_packet_header_47(proc_6_io_packet_header_47),
    .io_packet_header_48(proc_6_io_packet_header_48),
    .io_packet_header_49(proc_6_io_packet_header_49),
    .io_packet_header_50(proc_6_io_packet_header_50),
    .io_packet_header_51(proc_6_io_packet_header_51),
    .io_packet_header_52(proc_6_io_packet_header_52),
    .io_packet_header_53(proc_6_io_packet_header_53),
    .io_packet_header_54(proc_6_io_packet_header_54),
    .io_packet_header_55(proc_6_io_packet_header_55),
    .io_packet_header_56(proc_6_io_packet_header_56),
    .io_packet_header_57(proc_6_io_packet_header_57),
    .io_packet_header_58(proc_6_io_packet_header_58),
    .io_packet_header_59(proc_6_io_packet_header_59),
    .io_packet_header_60(proc_6_io_packet_header_60),
    .io_packet_header_61(proc_6_io_packet_header_61),
    .io_packet_header_62(proc_6_io_packet_header_62),
    .io_packet_header_63(proc_6_io_packet_header_63),
    .io_end(proc_6_io_end),
    .io_mem_addr(proc_6_io_mem_addr),
    .io_mem_rdata(proc_6_io_mem_rdata),
    .io_ready(proc_6_io_ready),
    .io_mod_start(proc_6_io_mod_start),
    .io_mod_hit_action_addr(proc_6_io_mod_hit_action_addr),
    .io_mod_miss_action_addr(proc_6_io_mod_miss_action_addr),
    .io_mod_ps_mod_start(proc_6_io_mod_ps_mod_start),
    .io_mod_ps_mod_header_id(proc_6_io_mod_ps_mod_header_id),
    .io_mod_ps_mod_header_length(proc_6_io_mod_ps_mod_header_length),
    .io_mod_ps_mod_next_tag_start(proc_6_io_mod_ps_mod_next_tag_start),
    .io_mod_ps_mod_next_table_0(proc_6_io_mod_ps_mod_next_table_0),
    .io_mod_ps_mod_next_table_1(proc_6_io_mod_ps_mod_next_table_1),
    .io_mod_mt_mod_start(proc_6_io_mod_mt_mod_start),
    .io_mod_mt_mod_header_id(proc_6_io_mod_mt_mod_header_id),
    .io_mod_mt_mod_key_off(proc_6_io_mod_mt_mod_key_off),
    .io_mod_mt_mod_key_len(proc_6_io_mod_mt_mod_key_len),
    .io_mod_mt_mod_val_len(proc_6_io_mod_mt_mod_val_len),
    .io_mod_ex_mod_start(proc_6_io_mod_ex_mod_start),
    .io_mod_ex_mod_ops_0(proc_6_io_mod_ex_mod_ops_0),
    .io_mod_ex_mod_ops_1(proc_6_io_mod_ex_mod_ops_1),
    .io_mod_ex_mod_ops_2(proc_6_io_mod_ex_mod_ops_2),
    .io_mod_ex_mod_ops_3(proc_6_io_mod_ex_mod_ops_3),
    .io_mod_ex_mod_ops_4(proc_6_io_mod_ex_mod_ops_4),
    .io_mod_ex_mod_ops_5(proc_6_io_mod_ex_mod_ops_5),
    .io_mod_ex_mod_ops_6(proc_6_io_mod_ex_mod_ops_6),
    .io_mod_ex_mod_ops_7(proc_6_io_mod_ex_mod_ops_7),
    .io_mod_ex_mod_ops_8(proc_6_io_mod_ex_mod_ops_8),
    .io_mod_ex_mod_ops_9(proc_6_io_mod_ex_mod_ops_9),
    .io_mod_ex_mod_ops_10(proc_6_io_mod_ex_mod_ops_10),
    .io_mod_ex_mod_ops_11(proc_6_io_mod_ex_mod_ops_11),
    .io_mod_ex_mod_ops_12(proc_6_io_mod_ex_mod_ops_12),
    .io_mod_ex_mod_ops_13(proc_6_io_mod_ex_mod_ops_13),
    .io_mod_ex_mod_ops_14(proc_6_io_mod_ex_mod_ops_14),
    .io_mod_ex_mod_ops_15(proc_6_io_mod_ex_mod_ops_15),
    .io_next_en(proc_6_io_next_en),
    .io_next_header_0(proc_6_io_next_header_0),
    .io_next_header_1(proc_6_io_next_header_1),
    .io_next_header_2(proc_6_io_next_header_2),
    .io_next_header_3(proc_6_io_next_header_3),
    .io_next_header_4(proc_6_io_next_header_4),
    .io_next_header_5(proc_6_io_next_header_5),
    .io_next_header_6(proc_6_io_next_header_6),
    .io_next_header_7(proc_6_io_next_header_7),
    .io_next_header_8(proc_6_io_next_header_8),
    .io_next_header_9(proc_6_io_next_header_9),
    .io_next_header_10(proc_6_io_next_header_10),
    .io_next_header_11(proc_6_io_next_header_11),
    .io_next_header_12(proc_6_io_next_header_12),
    .io_next_header_13(proc_6_io_next_header_13),
    .io_next_header_14(proc_6_io_next_header_14),
    .io_next_header_15(proc_6_io_next_header_15),
    .io_next_header_16(proc_6_io_next_header_16),
    .io_next_header_17(proc_6_io_next_header_17),
    .io_next_header_18(proc_6_io_next_header_18),
    .io_next_header_19(proc_6_io_next_header_19),
    .io_next_header_20(proc_6_io_next_header_20),
    .io_next_header_21(proc_6_io_next_header_21),
    .io_next_header_22(proc_6_io_next_header_22),
    .io_next_header_23(proc_6_io_next_header_23),
    .io_next_header_24(proc_6_io_next_header_24),
    .io_next_header_25(proc_6_io_next_header_25),
    .io_next_header_26(proc_6_io_next_header_26),
    .io_next_header_27(proc_6_io_next_header_27),
    .io_next_header_28(proc_6_io_next_header_28),
    .io_next_header_29(proc_6_io_next_header_29),
    .io_next_header_30(proc_6_io_next_header_30),
    .io_next_header_31(proc_6_io_next_header_31),
    .io_next_header_32(proc_6_io_next_header_32),
    .io_next_header_33(proc_6_io_next_header_33),
    .io_next_header_34(proc_6_io_next_header_34),
    .io_next_header_35(proc_6_io_next_header_35),
    .io_next_header_36(proc_6_io_next_header_36),
    .io_next_header_37(proc_6_io_next_header_37),
    .io_next_header_38(proc_6_io_next_header_38),
    .io_next_header_39(proc_6_io_next_header_39),
    .io_next_header_40(proc_6_io_next_header_40),
    .io_next_header_41(proc_6_io_next_header_41),
    .io_next_header_42(proc_6_io_next_header_42),
    .io_next_header_43(proc_6_io_next_header_43),
    .io_next_header_44(proc_6_io_next_header_44),
    .io_next_header_45(proc_6_io_next_header_45),
    .io_next_header_46(proc_6_io_next_header_46),
    .io_next_header_47(proc_6_io_next_header_47),
    .io_next_header_48(proc_6_io_next_header_48),
    .io_next_header_49(proc_6_io_next_header_49),
    .io_next_header_50(proc_6_io_next_header_50),
    .io_next_header_51(proc_6_io_next_header_51),
    .io_next_header_52(proc_6_io_next_header_52),
    .io_next_header_53(proc_6_io_next_header_53),
    .io_next_header_54(proc_6_io_next_header_54),
    .io_next_header_55(proc_6_io_next_header_55),
    .io_next_header_56(proc_6_io_next_header_56),
    .io_next_header_57(proc_6_io_next_header_57),
    .io_next_header_58(proc_6_io_next_header_58),
    .io_next_header_59(proc_6_io_next_header_59),
    .io_next_header_60(proc_6_io_next_header_60),
    .io_next_header_61(proc_6_io_next_header_61),
    .io_next_header_62(proc_6_io_next_header_62),
    .io_next_header_63(proc_6_io_next_header_63),
    .io_next_proc(proc_6_io_next_proc)
  );
  ProcessorController proc_7 ( // @[controller.scala 29:25]
    .clock(proc_7_clock),
    .reset(proc_7_reset),
    .io_update(proc_7_io_update),
    .io_packet_header_0(proc_7_io_packet_header_0),
    .io_packet_header_1(proc_7_io_packet_header_1),
    .io_packet_header_2(proc_7_io_packet_header_2),
    .io_packet_header_3(proc_7_io_packet_header_3),
    .io_packet_header_4(proc_7_io_packet_header_4),
    .io_packet_header_5(proc_7_io_packet_header_5),
    .io_packet_header_6(proc_7_io_packet_header_6),
    .io_packet_header_7(proc_7_io_packet_header_7),
    .io_packet_header_8(proc_7_io_packet_header_8),
    .io_packet_header_9(proc_7_io_packet_header_9),
    .io_packet_header_10(proc_7_io_packet_header_10),
    .io_packet_header_11(proc_7_io_packet_header_11),
    .io_packet_header_12(proc_7_io_packet_header_12),
    .io_packet_header_13(proc_7_io_packet_header_13),
    .io_packet_header_14(proc_7_io_packet_header_14),
    .io_packet_header_15(proc_7_io_packet_header_15),
    .io_packet_header_16(proc_7_io_packet_header_16),
    .io_packet_header_17(proc_7_io_packet_header_17),
    .io_packet_header_18(proc_7_io_packet_header_18),
    .io_packet_header_19(proc_7_io_packet_header_19),
    .io_packet_header_20(proc_7_io_packet_header_20),
    .io_packet_header_21(proc_7_io_packet_header_21),
    .io_packet_header_22(proc_7_io_packet_header_22),
    .io_packet_header_23(proc_7_io_packet_header_23),
    .io_packet_header_24(proc_7_io_packet_header_24),
    .io_packet_header_25(proc_7_io_packet_header_25),
    .io_packet_header_26(proc_7_io_packet_header_26),
    .io_packet_header_27(proc_7_io_packet_header_27),
    .io_packet_header_28(proc_7_io_packet_header_28),
    .io_packet_header_29(proc_7_io_packet_header_29),
    .io_packet_header_30(proc_7_io_packet_header_30),
    .io_packet_header_31(proc_7_io_packet_header_31),
    .io_packet_header_32(proc_7_io_packet_header_32),
    .io_packet_header_33(proc_7_io_packet_header_33),
    .io_packet_header_34(proc_7_io_packet_header_34),
    .io_packet_header_35(proc_7_io_packet_header_35),
    .io_packet_header_36(proc_7_io_packet_header_36),
    .io_packet_header_37(proc_7_io_packet_header_37),
    .io_packet_header_38(proc_7_io_packet_header_38),
    .io_packet_header_39(proc_7_io_packet_header_39),
    .io_packet_header_40(proc_7_io_packet_header_40),
    .io_packet_header_41(proc_7_io_packet_header_41),
    .io_packet_header_42(proc_7_io_packet_header_42),
    .io_packet_header_43(proc_7_io_packet_header_43),
    .io_packet_header_44(proc_7_io_packet_header_44),
    .io_packet_header_45(proc_7_io_packet_header_45),
    .io_packet_header_46(proc_7_io_packet_header_46),
    .io_packet_header_47(proc_7_io_packet_header_47),
    .io_packet_header_48(proc_7_io_packet_header_48),
    .io_packet_header_49(proc_7_io_packet_header_49),
    .io_packet_header_50(proc_7_io_packet_header_50),
    .io_packet_header_51(proc_7_io_packet_header_51),
    .io_packet_header_52(proc_7_io_packet_header_52),
    .io_packet_header_53(proc_7_io_packet_header_53),
    .io_packet_header_54(proc_7_io_packet_header_54),
    .io_packet_header_55(proc_7_io_packet_header_55),
    .io_packet_header_56(proc_7_io_packet_header_56),
    .io_packet_header_57(proc_7_io_packet_header_57),
    .io_packet_header_58(proc_7_io_packet_header_58),
    .io_packet_header_59(proc_7_io_packet_header_59),
    .io_packet_header_60(proc_7_io_packet_header_60),
    .io_packet_header_61(proc_7_io_packet_header_61),
    .io_packet_header_62(proc_7_io_packet_header_62),
    .io_packet_header_63(proc_7_io_packet_header_63),
    .io_end(proc_7_io_end),
    .io_mem_addr(proc_7_io_mem_addr),
    .io_mem_rdata(proc_7_io_mem_rdata),
    .io_ready(proc_7_io_ready),
    .io_mod_start(proc_7_io_mod_start),
    .io_mod_hit_action_addr(proc_7_io_mod_hit_action_addr),
    .io_mod_miss_action_addr(proc_7_io_mod_miss_action_addr),
    .io_mod_ps_mod_start(proc_7_io_mod_ps_mod_start),
    .io_mod_ps_mod_header_id(proc_7_io_mod_ps_mod_header_id),
    .io_mod_ps_mod_header_length(proc_7_io_mod_ps_mod_header_length),
    .io_mod_ps_mod_next_tag_start(proc_7_io_mod_ps_mod_next_tag_start),
    .io_mod_ps_mod_next_table_0(proc_7_io_mod_ps_mod_next_table_0),
    .io_mod_ps_mod_next_table_1(proc_7_io_mod_ps_mod_next_table_1),
    .io_mod_mt_mod_start(proc_7_io_mod_mt_mod_start),
    .io_mod_mt_mod_header_id(proc_7_io_mod_mt_mod_header_id),
    .io_mod_mt_mod_key_off(proc_7_io_mod_mt_mod_key_off),
    .io_mod_mt_mod_key_len(proc_7_io_mod_mt_mod_key_len),
    .io_mod_mt_mod_val_len(proc_7_io_mod_mt_mod_val_len),
    .io_mod_ex_mod_start(proc_7_io_mod_ex_mod_start),
    .io_mod_ex_mod_ops_0(proc_7_io_mod_ex_mod_ops_0),
    .io_mod_ex_mod_ops_1(proc_7_io_mod_ex_mod_ops_1),
    .io_mod_ex_mod_ops_2(proc_7_io_mod_ex_mod_ops_2),
    .io_mod_ex_mod_ops_3(proc_7_io_mod_ex_mod_ops_3),
    .io_mod_ex_mod_ops_4(proc_7_io_mod_ex_mod_ops_4),
    .io_mod_ex_mod_ops_5(proc_7_io_mod_ex_mod_ops_5),
    .io_mod_ex_mod_ops_6(proc_7_io_mod_ex_mod_ops_6),
    .io_mod_ex_mod_ops_7(proc_7_io_mod_ex_mod_ops_7),
    .io_mod_ex_mod_ops_8(proc_7_io_mod_ex_mod_ops_8),
    .io_mod_ex_mod_ops_9(proc_7_io_mod_ex_mod_ops_9),
    .io_mod_ex_mod_ops_10(proc_7_io_mod_ex_mod_ops_10),
    .io_mod_ex_mod_ops_11(proc_7_io_mod_ex_mod_ops_11),
    .io_mod_ex_mod_ops_12(proc_7_io_mod_ex_mod_ops_12),
    .io_mod_ex_mod_ops_13(proc_7_io_mod_ex_mod_ops_13),
    .io_mod_ex_mod_ops_14(proc_7_io_mod_ex_mod_ops_14),
    .io_mod_ex_mod_ops_15(proc_7_io_mod_ex_mod_ops_15),
    .io_next_en(proc_7_io_next_en),
    .io_next_header_0(proc_7_io_next_header_0),
    .io_next_header_1(proc_7_io_next_header_1),
    .io_next_header_2(proc_7_io_next_header_2),
    .io_next_header_3(proc_7_io_next_header_3),
    .io_next_header_4(proc_7_io_next_header_4),
    .io_next_header_5(proc_7_io_next_header_5),
    .io_next_header_6(proc_7_io_next_header_6),
    .io_next_header_7(proc_7_io_next_header_7),
    .io_next_header_8(proc_7_io_next_header_8),
    .io_next_header_9(proc_7_io_next_header_9),
    .io_next_header_10(proc_7_io_next_header_10),
    .io_next_header_11(proc_7_io_next_header_11),
    .io_next_header_12(proc_7_io_next_header_12),
    .io_next_header_13(proc_7_io_next_header_13),
    .io_next_header_14(proc_7_io_next_header_14),
    .io_next_header_15(proc_7_io_next_header_15),
    .io_next_header_16(proc_7_io_next_header_16),
    .io_next_header_17(proc_7_io_next_header_17),
    .io_next_header_18(proc_7_io_next_header_18),
    .io_next_header_19(proc_7_io_next_header_19),
    .io_next_header_20(proc_7_io_next_header_20),
    .io_next_header_21(proc_7_io_next_header_21),
    .io_next_header_22(proc_7_io_next_header_22),
    .io_next_header_23(proc_7_io_next_header_23),
    .io_next_header_24(proc_7_io_next_header_24),
    .io_next_header_25(proc_7_io_next_header_25),
    .io_next_header_26(proc_7_io_next_header_26),
    .io_next_header_27(proc_7_io_next_header_27),
    .io_next_header_28(proc_7_io_next_header_28),
    .io_next_header_29(proc_7_io_next_header_29),
    .io_next_header_30(proc_7_io_next_header_30),
    .io_next_header_31(proc_7_io_next_header_31),
    .io_next_header_32(proc_7_io_next_header_32),
    .io_next_header_33(proc_7_io_next_header_33),
    .io_next_header_34(proc_7_io_next_header_34),
    .io_next_header_35(proc_7_io_next_header_35),
    .io_next_header_36(proc_7_io_next_header_36),
    .io_next_header_37(proc_7_io_next_header_37),
    .io_next_header_38(proc_7_io_next_header_38),
    .io_next_header_39(proc_7_io_next_header_39),
    .io_next_header_40(proc_7_io_next_header_40),
    .io_next_header_41(proc_7_io_next_header_41),
    .io_next_header_42(proc_7_io_next_header_42),
    .io_next_header_43(proc_7_io_next_header_43),
    .io_next_header_44(proc_7_io_next_header_44),
    .io_next_header_45(proc_7_io_next_header_45),
    .io_next_header_46(proc_7_io_next_header_46),
    .io_next_header_47(proc_7_io_next_header_47),
    .io_next_header_48(proc_7_io_next_header_48),
    .io_next_header_49(proc_7_io_next_header_49),
    .io_next_header_50(proc_7_io_next_header_50),
    .io_next_header_51(proc_7_io_next_header_51),
    .io_next_header_52(proc_7_io_next_header_52),
    .io_next_header_53(proc_7_io_next_header_53),
    .io_next_header_54(proc_7_io_next_header_54),
    .io_next_header_55(proc_7_io_next_header_55),
    .io_next_header_56(proc_7_io_next_header_56),
    .io_next_header_57(proc_7_io_next_header_57),
    .io_next_header_58(proc_7_io_next_header_58),
    .io_next_header_59(proc_7_io_next_header_59),
    .io_next_header_60(proc_7_io_next_header_60),
    .io_next_header_61(proc_7_io_next_header_61),
    .io_next_header_62(proc_7_io_next_header_62),
    .io_next_header_63(proc_7_io_next_header_63),
    .io_next_proc(proc_7_io_next_proc)
  );
  assign io_ready_0 = proc_0_io_ready; // @[controller.scala 99:21]
  assign io_ready_1 = proc_1_io_ready; // @[controller.scala 99:21]
  assign io_ready_2 = proc_2_io_ready; // @[controller.scala 99:21]
  assign io_ready_3 = proc_3_io_ready; // @[controller.scala 99:21]
  assign io_ready_4 = proc_4_io_ready; // @[controller.scala 99:21]
  assign io_ready_5 = proc_5_io_ready; // @[controller.scala 99:21]
  assign io_ready_6 = proc_6_io_ready; // @[controller.scala 99:21]
  assign io_ready_7 = proc_7_io_ready; // @[controller.scala 99:21]
  assign mem_0_clock = clock;
  assign mem_0_io_mem_a_addr = proc_0_io_mem_addr; // @[controller.scala 32:24]
  assign mem_0_io_mem_b_addr = proc_1_io_mem_addr; // @[controller.scala 34:24]
  assign mem_1_clock = clock;
  assign mem_1_io_mem_a_addr = proc_2_io_mem_addr; // @[controller.scala 32:24]
  assign mem_1_io_mem_b_addr = proc_3_io_mem_addr; // @[controller.scala 34:24]
  assign mem_2_clock = clock;
  assign mem_2_io_mem_a_addr = proc_4_io_mem_addr; // @[controller.scala 32:24]
  assign mem_2_io_mem_b_addr = proc_5_io_mem_addr; // @[controller.scala 34:24]
  assign mem_3_clock = clock;
  assign mem_3_io_mem_a_addr = proc_6_io_mem_addr; // @[controller.scala 32:24]
  assign mem_3_io_mem_b_addr = proc_7_io_mem_addr; // @[controller.scala 34:24]
  assign encoders_0_io_input = {next_table_hi,next_table_lo}; // @[Cat.scala 30:58]
  assign encoders_1_io_input = {next_table_hi_1,next_table_lo_1}; // @[Cat.scala 30:58]
  assign encoders_2_io_input = {next_table_hi_2,next_table_lo_2}; // @[Cat.scala 30:58]
  assign encoders_3_io_input = {next_table_hi_3,next_table_lo_3}; // @[Cat.scala 30:58]
  assign encoders_4_io_input = {next_table_hi_4,next_table_lo_4}; // @[Cat.scala 30:58]
  assign encoders_5_io_input = {next_table_hi_5,next_table_lo_5}; // @[Cat.scala 30:58]
  assign encoders_6_io_input = {next_table_hi_6,next_table_lo_6}; // @[Cat.scala 30:58]
  assign encoders_7_io_input = {next_table_hi_7,next_table_lo_7}; // @[Cat.scala 30:58]
  assign proc_0_clock = clock;
  assign proc_0_reset = reset;
  assign proc_0_io_update = encoders_0_io_valid & proc_0_io_ready | io_start & proc_0_io_ready; // @[controller.scala 89:57 controller.scala 91:31 controller.scala 37:27]
  assign proc_0_io_packet_header_0 = encoders_0_io_valid & proc_0_io_ready ? _GEN_704 : io_packet_header_0; // @[controller.scala 89:57 controller.scala 38:34]
  assign proc_0_io_packet_header_1 = encoders_0_io_valid & proc_0_io_ready ? _GEN_705 : io_packet_header_1; // @[controller.scala 89:57 controller.scala 38:34]
  assign proc_0_io_packet_header_2 = encoders_0_io_valid & proc_0_io_ready ? _GEN_706 : io_packet_header_2; // @[controller.scala 89:57 controller.scala 38:34]
  assign proc_0_io_packet_header_3 = encoders_0_io_valid & proc_0_io_ready ? _GEN_707 : io_packet_header_3; // @[controller.scala 89:57 controller.scala 38:34]
  assign proc_0_io_packet_header_4 = encoders_0_io_valid & proc_0_io_ready ? _GEN_708 : io_packet_header_4; // @[controller.scala 89:57 controller.scala 38:34]
  assign proc_0_io_packet_header_5 = encoders_0_io_valid & proc_0_io_ready ? _GEN_709 : io_packet_header_5; // @[controller.scala 89:57 controller.scala 38:34]
  assign proc_0_io_packet_header_6 = encoders_0_io_valid & proc_0_io_ready ? _GEN_710 : io_packet_header_6; // @[controller.scala 89:57 controller.scala 38:34]
  assign proc_0_io_packet_header_7 = encoders_0_io_valid & proc_0_io_ready ? _GEN_711 : io_packet_header_7; // @[controller.scala 89:57 controller.scala 38:34]
  assign proc_0_io_packet_header_8 = encoders_0_io_valid & proc_0_io_ready ? _GEN_712 : io_packet_header_8; // @[controller.scala 89:57 controller.scala 38:34]
  assign proc_0_io_packet_header_9 = encoders_0_io_valid & proc_0_io_ready ? _GEN_713 : io_packet_header_9; // @[controller.scala 89:57 controller.scala 38:34]
  assign proc_0_io_packet_header_10 = encoders_0_io_valid & proc_0_io_ready ? _GEN_714 : io_packet_header_10; // @[controller.scala 89:57 controller.scala 38:34]
  assign proc_0_io_packet_header_11 = encoders_0_io_valid & proc_0_io_ready ? _GEN_715 : io_packet_header_11; // @[controller.scala 89:57 controller.scala 38:34]
  assign proc_0_io_packet_header_12 = encoders_0_io_valid & proc_0_io_ready ? _GEN_716 : io_packet_header_12; // @[controller.scala 89:57 controller.scala 38:34]
  assign proc_0_io_packet_header_13 = encoders_0_io_valid & proc_0_io_ready ? _GEN_717 : io_packet_header_13; // @[controller.scala 89:57 controller.scala 38:34]
  assign proc_0_io_packet_header_14 = encoders_0_io_valid & proc_0_io_ready ? _GEN_718 : io_packet_header_14; // @[controller.scala 89:57 controller.scala 38:34]
  assign proc_0_io_packet_header_15 = encoders_0_io_valid & proc_0_io_ready ? _GEN_719 : io_packet_header_15; // @[controller.scala 89:57 controller.scala 38:34]
  assign proc_0_io_packet_header_16 = encoders_0_io_valid & proc_0_io_ready ? _GEN_720 : io_packet_header_16; // @[controller.scala 89:57 controller.scala 38:34]
  assign proc_0_io_packet_header_17 = encoders_0_io_valid & proc_0_io_ready ? _GEN_721 : io_packet_header_17; // @[controller.scala 89:57 controller.scala 38:34]
  assign proc_0_io_packet_header_18 = encoders_0_io_valid & proc_0_io_ready ? _GEN_722 : io_packet_header_18; // @[controller.scala 89:57 controller.scala 38:34]
  assign proc_0_io_packet_header_19 = encoders_0_io_valid & proc_0_io_ready ? _GEN_723 : io_packet_header_19; // @[controller.scala 89:57 controller.scala 38:34]
  assign proc_0_io_packet_header_20 = encoders_0_io_valid & proc_0_io_ready ? _GEN_724 : io_packet_header_20; // @[controller.scala 89:57 controller.scala 38:34]
  assign proc_0_io_packet_header_21 = encoders_0_io_valid & proc_0_io_ready ? _GEN_725 : io_packet_header_21; // @[controller.scala 89:57 controller.scala 38:34]
  assign proc_0_io_packet_header_22 = encoders_0_io_valid & proc_0_io_ready ? _GEN_726 : io_packet_header_22; // @[controller.scala 89:57 controller.scala 38:34]
  assign proc_0_io_packet_header_23 = encoders_0_io_valid & proc_0_io_ready ? _GEN_727 : io_packet_header_23; // @[controller.scala 89:57 controller.scala 38:34]
  assign proc_0_io_packet_header_24 = encoders_0_io_valid & proc_0_io_ready ? _GEN_728 : io_packet_header_24; // @[controller.scala 89:57 controller.scala 38:34]
  assign proc_0_io_packet_header_25 = encoders_0_io_valid & proc_0_io_ready ? _GEN_729 : io_packet_header_25; // @[controller.scala 89:57 controller.scala 38:34]
  assign proc_0_io_packet_header_26 = encoders_0_io_valid & proc_0_io_ready ? _GEN_730 : io_packet_header_26; // @[controller.scala 89:57 controller.scala 38:34]
  assign proc_0_io_packet_header_27 = encoders_0_io_valid & proc_0_io_ready ? _GEN_731 : io_packet_header_27; // @[controller.scala 89:57 controller.scala 38:34]
  assign proc_0_io_packet_header_28 = encoders_0_io_valid & proc_0_io_ready ? _GEN_732 : io_packet_header_28; // @[controller.scala 89:57 controller.scala 38:34]
  assign proc_0_io_packet_header_29 = encoders_0_io_valid & proc_0_io_ready ? _GEN_733 : io_packet_header_29; // @[controller.scala 89:57 controller.scala 38:34]
  assign proc_0_io_packet_header_30 = encoders_0_io_valid & proc_0_io_ready ? _GEN_734 : io_packet_header_30; // @[controller.scala 89:57 controller.scala 38:34]
  assign proc_0_io_packet_header_31 = encoders_0_io_valid & proc_0_io_ready ? _GEN_735 : io_packet_header_31; // @[controller.scala 89:57 controller.scala 38:34]
  assign proc_0_io_packet_header_32 = encoders_0_io_valid & proc_0_io_ready ? _GEN_736 : io_packet_header_32; // @[controller.scala 89:57 controller.scala 38:34]
  assign proc_0_io_packet_header_33 = encoders_0_io_valid & proc_0_io_ready ? _GEN_737 : io_packet_header_33; // @[controller.scala 89:57 controller.scala 38:34]
  assign proc_0_io_packet_header_34 = encoders_0_io_valid & proc_0_io_ready ? _GEN_738 : io_packet_header_34; // @[controller.scala 89:57 controller.scala 38:34]
  assign proc_0_io_packet_header_35 = encoders_0_io_valid & proc_0_io_ready ? _GEN_739 : io_packet_header_35; // @[controller.scala 89:57 controller.scala 38:34]
  assign proc_0_io_packet_header_36 = encoders_0_io_valid & proc_0_io_ready ? _GEN_740 : io_packet_header_36; // @[controller.scala 89:57 controller.scala 38:34]
  assign proc_0_io_packet_header_37 = encoders_0_io_valid & proc_0_io_ready ? _GEN_741 : io_packet_header_37; // @[controller.scala 89:57 controller.scala 38:34]
  assign proc_0_io_packet_header_38 = encoders_0_io_valid & proc_0_io_ready ? _GEN_742 : io_packet_header_38; // @[controller.scala 89:57 controller.scala 38:34]
  assign proc_0_io_packet_header_39 = encoders_0_io_valid & proc_0_io_ready ? _GEN_743 : io_packet_header_39; // @[controller.scala 89:57 controller.scala 38:34]
  assign proc_0_io_packet_header_40 = encoders_0_io_valid & proc_0_io_ready ? _GEN_744 : io_packet_header_40; // @[controller.scala 89:57 controller.scala 38:34]
  assign proc_0_io_packet_header_41 = encoders_0_io_valid & proc_0_io_ready ? _GEN_745 : io_packet_header_41; // @[controller.scala 89:57 controller.scala 38:34]
  assign proc_0_io_packet_header_42 = encoders_0_io_valid & proc_0_io_ready ? _GEN_746 : io_packet_header_42; // @[controller.scala 89:57 controller.scala 38:34]
  assign proc_0_io_packet_header_43 = encoders_0_io_valid & proc_0_io_ready ? _GEN_747 : io_packet_header_43; // @[controller.scala 89:57 controller.scala 38:34]
  assign proc_0_io_packet_header_44 = encoders_0_io_valid & proc_0_io_ready ? _GEN_748 : io_packet_header_44; // @[controller.scala 89:57 controller.scala 38:34]
  assign proc_0_io_packet_header_45 = encoders_0_io_valid & proc_0_io_ready ? _GEN_749 : io_packet_header_45; // @[controller.scala 89:57 controller.scala 38:34]
  assign proc_0_io_packet_header_46 = encoders_0_io_valid & proc_0_io_ready ? _GEN_750 : io_packet_header_46; // @[controller.scala 89:57 controller.scala 38:34]
  assign proc_0_io_packet_header_47 = encoders_0_io_valid & proc_0_io_ready ? _GEN_751 : io_packet_header_47; // @[controller.scala 89:57 controller.scala 38:34]
  assign proc_0_io_packet_header_48 = encoders_0_io_valid & proc_0_io_ready ? _GEN_752 : io_packet_header_48; // @[controller.scala 89:57 controller.scala 38:34]
  assign proc_0_io_packet_header_49 = encoders_0_io_valid & proc_0_io_ready ? _GEN_753 : io_packet_header_49; // @[controller.scala 89:57 controller.scala 38:34]
  assign proc_0_io_packet_header_50 = encoders_0_io_valid & proc_0_io_ready ? _GEN_754 : io_packet_header_50; // @[controller.scala 89:57 controller.scala 38:34]
  assign proc_0_io_packet_header_51 = encoders_0_io_valid & proc_0_io_ready ? _GEN_755 : io_packet_header_51; // @[controller.scala 89:57 controller.scala 38:34]
  assign proc_0_io_packet_header_52 = encoders_0_io_valid & proc_0_io_ready ? _GEN_756 : io_packet_header_52; // @[controller.scala 89:57 controller.scala 38:34]
  assign proc_0_io_packet_header_53 = encoders_0_io_valid & proc_0_io_ready ? _GEN_757 : io_packet_header_53; // @[controller.scala 89:57 controller.scala 38:34]
  assign proc_0_io_packet_header_54 = encoders_0_io_valid & proc_0_io_ready ? _GEN_758 : io_packet_header_54; // @[controller.scala 89:57 controller.scala 38:34]
  assign proc_0_io_packet_header_55 = encoders_0_io_valid & proc_0_io_ready ? _GEN_759 : io_packet_header_55; // @[controller.scala 89:57 controller.scala 38:34]
  assign proc_0_io_packet_header_56 = encoders_0_io_valid & proc_0_io_ready ? _GEN_760 : io_packet_header_56; // @[controller.scala 89:57 controller.scala 38:34]
  assign proc_0_io_packet_header_57 = encoders_0_io_valid & proc_0_io_ready ? _GEN_761 : io_packet_header_57; // @[controller.scala 89:57 controller.scala 38:34]
  assign proc_0_io_packet_header_58 = encoders_0_io_valid & proc_0_io_ready ? _GEN_762 : io_packet_header_58; // @[controller.scala 89:57 controller.scala 38:34]
  assign proc_0_io_packet_header_59 = encoders_0_io_valid & proc_0_io_ready ? _GEN_763 : io_packet_header_59; // @[controller.scala 89:57 controller.scala 38:34]
  assign proc_0_io_packet_header_60 = encoders_0_io_valid & proc_0_io_ready ? _GEN_764 : io_packet_header_60; // @[controller.scala 89:57 controller.scala 38:34]
  assign proc_0_io_packet_header_61 = encoders_0_io_valid & proc_0_io_ready ? _GEN_765 : io_packet_header_61; // @[controller.scala 89:57 controller.scala 38:34]
  assign proc_0_io_packet_header_62 = encoders_0_io_valid & proc_0_io_ready ? _GEN_766 : io_packet_header_62; // @[controller.scala 89:57 controller.scala 38:34]
  assign proc_0_io_packet_header_63 = encoders_0_io_valid & proc_0_io_ready ? _GEN_767 : io_packet_header_63; // @[controller.scala 89:57 controller.scala 38:34]
  assign proc_0_io_end = encoders_0_io_valid & proc_0_io_ready; // @[controller.scala 89:36]
  assign proc_0_io_mem_rdata = mem_0_io_mem_a_rdata; // @[controller.scala 32:24]
  assign proc_0_io_mod_start = io_mod_proc == 3'h0 & io_mod_start; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 52:34]
  assign proc_0_io_mod_hit_action_addr = io_mod_proc == 3'h0 ? io_mod_hit_action_addr : 32'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 53:44]
  assign proc_0_io_mod_miss_action_addr = io_mod_proc == 3'h0 ? io_mod_miss_action_addr : 32'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 54:45]
  assign proc_0_io_mod_ps_mod_start = io_mod_proc == 3'h0 & io_mod_ps_mod_start; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 55:41]
  assign proc_0_io_mod_ps_mod_header_id = io_mod_proc == 3'h0 & io_mod_ps_mod_header_id; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 56:45]
  assign proc_0_io_mod_ps_mod_header_length = io_mod_proc == 3'h0 ? io_mod_ps_mod_header_length : 32'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 57:49]
  assign proc_0_io_mod_ps_mod_next_tag_start = io_mod_proc == 3'h0 ? io_mod_ps_mod_next_tag_start : 32'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 58:50]
  assign proc_0_io_mod_ps_mod_next_table_0 = io_mod_proc == 3'h0 ? io_mod_ps_mod_next_table_0 : 32'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 61:53]
  assign proc_0_io_mod_ps_mod_next_table_1 = io_mod_proc == 3'h0 ? io_mod_ps_mod_next_table_1 : 32'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 61:53]
  assign proc_0_io_mod_mt_mod_start = io_mod_proc == 3'h0 & io_mod_mt_mod_start; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 63:41]
  assign proc_0_io_mod_mt_mod_header_id = io_mod_proc == 3'h0 ? io_mod_mt_mod_header_id : 4'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 64:45]
  assign proc_0_io_mod_mt_mod_key_off = io_mod_proc == 3'h0 ? io_mod_mt_mod_key_off : 6'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 65:43]
  assign proc_0_io_mod_mt_mod_key_len = io_mod_proc == 3'h0 ? io_mod_mt_mod_key_len : 6'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 66:43]
  assign proc_0_io_mod_mt_mod_val_len = io_mod_proc == 3'h0 ? io_mod_mt_mod_val_len : 6'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 67:43]
  assign proc_0_io_mod_ex_mod_start = io_mod_proc == 3'h0 & io_mod_ex_mod_start; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 68:41]
  assign proc_0_io_mod_ex_mod_ops_0 = io_mod_proc == 3'h0 ? io_mod_ex_mod_ops_0 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_0_io_mod_ex_mod_ops_1 = io_mod_proc == 3'h0 ? io_mod_ex_mod_ops_1 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_0_io_mod_ex_mod_ops_2 = io_mod_proc == 3'h0 ? io_mod_ex_mod_ops_2 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_0_io_mod_ex_mod_ops_3 = io_mod_proc == 3'h0 ? io_mod_ex_mod_ops_3 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_0_io_mod_ex_mod_ops_4 = io_mod_proc == 3'h0 ? io_mod_ex_mod_ops_4 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_0_io_mod_ex_mod_ops_5 = io_mod_proc == 3'h0 ? io_mod_ex_mod_ops_5 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_0_io_mod_ex_mod_ops_6 = io_mod_proc == 3'h0 ? io_mod_ex_mod_ops_6 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_0_io_mod_ex_mod_ops_7 = io_mod_proc == 3'h0 ? io_mod_ex_mod_ops_7 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_0_io_mod_ex_mod_ops_8 = io_mod_proc == 3'h0 ? io_mod_ex_mod_ops_8 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_0_io_mod_ex_mod_ops_9 = io_mod_proc == 3'h0 ? io_mod_ex_mod_ops_9 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_0_io_mod_ex_mod_ops_10 = io_mod_proc == 3'h0 ? io_mod_ex_mod_ops_10 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_0_io_mod_ex_mod_ops_11 = io_mod_proc == 3'h0 ? io_mod_ex_mod_ops_11 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_0_io_mod_ex_mod_ops_12 = io_mod_proc == 3'h0 ? io_mod_ex_mod_ops_12 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_0_io_mod_ex_mod_ops_13 = io_mod_proc == 3'h0 ? io_mod_ex_mod_ops_13 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_0_io_mod_ex_mod_ops_14 = io_mod_proc == 3'h0 ? io_mod_ex_mod_ops_14 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_0_io_mod_ex_mod_ops_15 = io_mod_proc == 3'h0 ? io_mod_ex_mod_ops_15 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_1_clock = clock;
  assign proc_1_reset = reset;
  assign proc_1_io_update = encoders_1_io_valid & proc_1_io_ready; // @[controller.scala 89:36]
  assign proc_1_io_packet_header_0 = encoders_1_io_valid & proc_1_io_ready ? _GEN_1282 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_1_io_packet_header_1 = encoders_1_io_valid & proc_1_io_ready ? _GEN_1283 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_1_io_packet_header_2 = encoders_1_io_valid & proc_1_io_ready ? _GEN_1284 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_1_io_packet_header_3 = encoders_1_io_valid & proc_1_io_ready ? _GEN_1285 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_1_io_packet_header_4 = encoders_1_io_valid & proc_1_io_ready ? _GEN_1286 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_1_io_packet_header_5 = encoders_1_io_valid & proc_1_io_ready ? _GEN_1287 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_1_io_packet_header_6 = encoders_1_io_valid & proc_1_io_ready ? _GEN_1288 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_1_io_packet_header_7 = encoders_1_io_valid & proc_1_io_ready ? _GEN_1289 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_1_io_packet_header_8 = encoders_1_io_valid & proc_1_io_ready ? _GEN_1290 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_1_io_packet_header_9 = encoders_1_io_valid & proc_1_io_ready ? _GEN_1291 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_1_io_packet_header_10 = encoders_1_io_valid & proc_1_io_ready ? _GEN_1292 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_1_io_packet_header_11 = encoders_1_io_valid & proc_1_io_ready ? _GEN_1293 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_1_io_packet_header_12 = encoders_1_io_valid & proc_1_io_ready ? _GEN_1294 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_1_io_packet_header_13 = encoders_1_io_valid & proc_1_io_ready ? _GEN_1295 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_1_io_packet_header_14 = encoders_1_io_valid & proc_1_io_ready ? _GEN_1296 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_1_io_packet_header_15 = encoders_1_io_valid & proc_1_io_ready ? _GEN_1297 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_1_io_packet_header_16 = encoders_1_io_valid & proc_1_io_ready ? _GEN_1298 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_1_io_packet_header_17 = encoders_1_io_valid & proc_1_io_ready ? _GEN_1299 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_1_io_packet_header_18 = encoders_1_io_valid & proc_1_io_ready ? _GEN_1300 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_1_io_packet_header_19 = encoders_1_io_valid & proc_1_io_ready ? _GEN_1301 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_1_io_packet_header_20 = encoders_1_io_valid & proc_1_io_ready ? _GEN_1302 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_1_io_packet_header_21 = encoders_1_io_valid & proc_1_io_ready ? _GEN_1303 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_1_io_packet_header_22 = encoders_1_io_valid & proc_1_io_ready ? _GEN_1304 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_1_io_packet_header_23 = encoders_1_io_valid & proc_1_io_ready ? _GEN_1305 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_1_io_packet_header_24 = encoders_1_io_valid & proc_1_io_ready ? _GEN_1306 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_1_io_packet_header_25 = encoders_1_io_valid & proc_1_io_ready ? _GEN_1307 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_1_io_packet_header_26 = encoders_1_io_valid & proc_1_io_ready ? _GEN_1308 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_1_io_packet_header_27 = encoders_1_io_valid & proc_1_io_ready ? _GEN_1309 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_1_io_packet_header_28 = encoders_1_io_valid & proc_1_io_ready ? _GEN_1310 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_1_io_packet_header_29 = encoders_1_io_valid & proc_1_io_ready ? _GEN_1311 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_1_io_packet_header_30 = encoders_1_io_valid & proc_1_io_ready ? _GEN_1312 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_1_io_packet_header_31 = encoders_1_io_valid & proc_1_io_ready ? _GEN_1313 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_1_io_packet_header_32 = encoders_1_io_valid & proc_1_io_ready ? _GEN_1314 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_1_io_packet_header_33 = encoders_1_io_valid & proc_1_io_ready ? _GEN_1315 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_1_io_packet_header_34 = encoders_1_io_valid & proc_1_io_ready ? _GEN_1316 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_1_io_packet_header_35 = encoders_1_io_valid & proc_1_io_ready ? _GEN_1317 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_1_io_packet_header_36 = encoders_1_io_valid & proc_1_io_ready ? _GEN_1318 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_1_io_packet_header_37 = encoders_1_io_valid & proc_1_io_ready ? _GEN_1319 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_1_io_packet_header_38 = encoders_1_io_valid & proc_1_io_ready ? _GEN_1320 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_1_io_packet_header_39 = encoders_1_io_valid & proc_1_io_ready ? _GEN_1321 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_1_io_packet_header_40 = encoders_1_io_valid & proc_1_io_ready ? _GEN_1322 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_1_io_packet_header_41 = encoders_1_io_valid & proc_1_io_ready ? _GEN_1323 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_1_io_packet_header_42 = encoders_1_io_valid & proc_1_io_ready ? _GEN_1324 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_1_io_packet_header_43 = encoders_1_io_valid & proc_1_io_ready ? _GEN_1325 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_1_io_packet_header_44 = encoders_1_io_valid & proc_1_io_ready ? _GEN_1326 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_1_io_packet_header_45 = encoders_1_io_valid & proc_1_io_ready ? _GEN_1327 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_1_io_packet_header_46 = encoders_1_io_valid & proc_1_io_ready ? _GEN_1328 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_1_io_packet_header_47 = encoders_1_io_valid & proc_1_io_ready ? _GEN_1329 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_1_io_packet_header_48 = encoders_1_io_valid & proc_1_io_ready ? _GEN_1330 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_1_io_packet_header_49 = encoders_1_io_valid & proc_1_io_ready ? _GEN_1331 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_1_io_packet_header_50 = encoders_1_io_valid & proc_1_io_ready ? _GEN_1332 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_1_io_packet_header_51 = encoders_1_io_valid & proc_1_io_ready ? _GEN_1333 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_1_io_packet_header_52 = encoders_1_io_valid & proc_1_io_ready ? _GEN_1334 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_1_io_packet_header_53 = encoders_1_io_valid & proc_1_io_ready ? _GEN_1335 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_1_io_packet_header_54 = encoders_1_io_valid & proc_1_io_ready ? _GEN_1336 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_1_io_packet_header_55 = encoders_1_io_valid & proc_1_io_ready ? _GEN_1337 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_1_io_packet_header_56 = encoders_1_io_valid & proc_1_io_ready ? _GEN_1338 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_1_io_packet_header_57 = encoders_1_io_valid & proc_1_io_ready ? _GEN_1339 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_1_io_packet_header_58 = encoders_1_io_valid & proc_1_io_ready ? _GEN_1340 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_1_io_packet_header_59 = encoders_1_io_valid & proc_1_io_ready ? _GEN_1341 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_1_io_packet_header_60 = encoders_1_io_valid & proc_1_io_ready ? _GEN_1342 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_1_io_packet_header_61 = encoders_1_io_valid & proc_1_io_ready ? _GEN_1343 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_1_io_packet_header_62 = encoders_1_io_valid & proc_1_io_ready ? _GEN_1344 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_1_io_packet_header_63 = encoders_1_io_valid & proc_1_io_ready ? _GEN_1345 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_1_io_end = encoders_1_io_valid & proc_1_io_ready; // @[controller.scala 89:36]
  assign proc_1_io_mem_rdata = mem_0_io_mem_b_rdata; // @[controller.scala 34:24]
  assign proc_1_io_mod_start = io_mod_proc == 3'h1 & io_mod_start; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 52:34]
  assign proc_1_io_mod_hit_action_addr = io_mod_proc == 3'h1 ? io_mod_hit_action_addr : 32'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 53:44]
  assign proc_1_io_mod_miss_action_addr = io_mod_proc == 3'h1 ? io_mod_miss_action_addr : 32'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 54:45]
  assign proc_1_io_mod_ps_mod_start = io_mod_proc == 3'h1 & io_mod_ps_mod_start; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 55:41]
  assign proc_1_io_mod_ps_mod_header_id = io_mod_proc == 3'h1 & io_mod_ps_mod_header_id; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 56:45]
  assign proc_1_io_mod_ps_mod_header_length = io_mod_proc == 3'h1 ? io_mod_ps_mod_header_length : 32'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 57:49]
  assign proc_1_io_mod_ps_mod_next_tag_start = io_mod_proc == 3'h1 ? io_mod_ps_mod_next_tag_start : 32'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 58:50]
  assign proc_1_io_mod_ps_mod_next_table_0 = io_mod_proc == 3'h1 ? io_mod_ps_mod_next_table_0 : 32'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 61:53]
  assign proc_1_io_mod_ps_mod_next_table_1 = io_mod_proc == 3'h1 ? io_mod_ps_mod_next_table_1 : 32'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 61:53]
  assign proc_1_io_mod_mt_mod_start = io_mod_proc == 3'h1 & io_mod_mt_mod_start; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 63:41]
  assign proc_1_io_mod_mt_mod_header_id = io_mod_proc == 3'h1 ? io_mod_mt_mod_header_id : 4'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 64:45]
  assign proc_1_io_mod_mt_mod_key_off = io_mod_proc == 3'h1 ? io_mod_mt_mod_key_off : 6'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 65:43]
  assign proc_1_io_mod_mt_mod_key_len = io_mod_proc == 3'h1 ? io_mod_mt_mod_key_len : 6'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 66:43]
  assign proc_1_io_mod_mt_mod_val_len = io_mod_proc == 3'h1 ? io_mod_mt_mod_val_len : 6'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 67:43]
  assign proc_1_io_mod_ex_mod_start = io_mod_proc == 3'h1 & io_mod_ex_mod_start; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 68:41]
  assign proc_1_io_mod_ex_mod_ops_0 = io_mod_proc == 3'h1 ? io_mod_ex_mod_ops_0 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_1_io_mod_ex_mod_ops_1 = io_mod_proc == 3'h1 ? io_mod_ex_mod_ops_1 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_1_io_mod_ex_mod_ops_2 = io_mod_proc == 3'h1 ? io_mod_ex_mod_ops_2 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_1_io_mod_ex_mod_ops_3 = io_mod_proc == 3'h1 ? io_mod_ex_mod_ops_3 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_1_io_mod_ex_mod_ops_4 = io_mod_proc == 3'h1 ? io_mod_ex_mod_ops_4 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_1_io_mod_ex_mod_ops_5 = io_mod_proc == 3'h1 ? io_mod_ex_mod_ops_5 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_1_io_mod_ex_mod_ops_6 = io_mod_proc == 3'h1 ? io_mod_ex_mod_ops_6 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_1_io_mod_ex_mod_ops_7 = io_mod_proc == 3'h1 ? io_mod_ex_mod_ops_7 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_1_io_mod_ex_mod_ops_8 = io_mod_proc == 3'h1 ? io_mod_ex_mod_ops_8 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_1_io_mod_ex_mod_ops_9 = io_mod_proc == 3'h1 ? io_mod_ex_mod_ops_9 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_1_io_mod_ex_mod_ops_10 = io_mod_proc == 3'h1 ? io_mod_ex_mod_ops_10 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_1_io_mod_ex_mod_ops_11 = io_mod_proc == 3'h1 ? io_mod_ex_mod_ops_11 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_1_io_mod_ex_mod_ops_12 = io_mod_proc == 3'h1 ? io_mod_ex_mod_ops_12 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_1_io_mod_ex_mod_ops_13 = io_mod_proc == 3'h1 ? io_mod_ex_mod_ops_13 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_1_io_mod_ex_mod_ops_14 = io_mod_proc == 3'h1 ? io_mod_ex_mod_ops_14 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_1_io_mod_ex_mod_ops_15 = io_mod_proc == 3'h1 ? io_mod_ex_mod_ops_15 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_2_clock = clock;
  assign proc_2_reset = reset;
  assign proc_2_io_update = encoders_2_io_valid & proc_2_io_ready; // @[controller.scala 89:36]
  assign proc_2_io_packet_header_0 = encoders_2_io_valid & proc_2_io_ready ? _GEN_1859 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_2_io_packet_header_1 = encoders_2_io_valid & proc_2_io_ready ? _GEN_1860 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_2_io_packet_header_2 = encoders_2_io_valid & proc_2_io_ready ? _GEN_1861 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_2_io_packet_header_3 = encoders_2_io_valid & proc_2_io_ready ? _GEN_1862 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_2_io_packet_header_4 = encoders_2_io_valid & proc_2_io_ready ? _GEN_1863 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_2_io_packet_header_5 = encoders_2_io_valid & proc_2_io_ready ? _GEN_1864 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_2_io_packet_header_6 = encoders_2_io_valid & proc_2_io_ready ? _GEN_1865 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_2_io_packet_header_7 = encoders_2_io_valid & proc_2_io_ready ? _GEN_1866 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_2_io_packet_header_8 = encoders_2_io_valid & proc_2_io_ready ? _GEN_1867 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_2_io_packet_header_9 = encoders_2_io_valid & proc_2_io_ready ? _GEN_1868 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_2_io_packet_header_10 = encoders_2_io_valid & proc_2_io_ready ? _GEN_1869 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_2_io_packet_header_11 = encoders_2_io_valid & proc_2_io_ready ? _GEN_1870 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_2_io_packet_header_12 = encoders_2_io_valid & proc_2_io_ready ? _GEN_1871 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_2_io_packet_header_13 = encoders_2_io_valid & proc_2_io_ready ? _GEN_1872 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_2_io_packet_header_14 = encoders_2_io_valid & proc_2_io_ready ? _GEN_1873 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_2_io_packet_header_15 = encoders_2_io_valid & proc_2_io_ready ? _GEN_1874 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_2_io_packet_header_16 = encoders_2_io_valid & proc_2_io_ready ? _GEN_1875 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_2_io_packet_header_17 = encoders_2_io_valid & proc_2_io_ready ? _GEN_1876 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_2_io_packet_header_18 = encoders_2_io_valid & proc_2_io_ready ? _GEN_1877 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_2_io_packet_header_19 = encoders_2_io_valid & proc_2_io_ready ? _GEN_1878 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_2_io_packet_header_20 = encoders_2_io_valid & proc_2_io_ready ? _GEN_1879 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_2_io_packet_header_21 = encoders_2_io_valid & proc_2_io_ready ? _GEN_1880 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_2_io_packet_header_22 = encoders_2_io_valid & proc_2_io_ready ? _GEN_1881 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_2_io_packet_header_23 = encoders_2_io_valid & proc_2_io_ready ? _GEN_1882 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_2_io_packet_header_24 = encoders_2_io_valid & proc_2_io_ready ? _GEN_1883 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_2_io_packet_header_25 = encoders_2_io_valid & proc_2_io_ready ? _GEN_1884 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_2_io_packet_header_26 = encoders_2_io_valid & proc_2_io_ready ? _GEN_1885 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_2_io_packet_header_27 = encoders_2_io_valid & proc_2_io_ready ? _GEN_1886 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_2_io_packet_header_28 = encoders_2_io_valid & proc_2_io_ready ? _GEN_1887 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_2_io_packet_header_29 = encoders_2_io_valid & proc_2_io_ready ? _GEN_1888 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_2_io_packet_header_30 = encoders_2_io_valid & proc_2_io_ready ? _GEN_1889 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_2_io_packet_header_31 = encoders_2_io_valid & proc_2_io_ready ? _GEN_1890 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_2_io_packet_header_32 = encoders_2_io_valid & proc_2_io_ready ? _GEN_1891 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_2_io_packet_header_33 = encoders_2_io_valid & proc_2_io_ready ? _GEN_1892 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_2_io_packet_header_34 = encoders_2_io_valid & proc_2_io_ready ? _GEN_1893 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_2_io_packet_header_35 = encoders_2_io_valid & proc_2_io_ready ? _GEN_1894 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_2_io_packet_header_36 = encoders_2_io_valid & proc_2_io_ready ? _GEN_1895 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_2_io_packet_header_37 = encoders_2_io_valid & proc_2_io_ready ? _GEN_1896 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_2_io_packet_header_38 = encoders_2_io_valid & proc_2_io_ready ? _GEN_1897 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_2_io_packet_header_39 = encoders_2_io_valid & proc_2_io_ready ? _GEN_1898 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_2_io_packet_header_40 = encoders_2_io_valid & proc_2_io_ready ? _GEN_1899 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_2_io_packet_header_41 = encoders_2_io_valid & proc_2_io_ready ? _GEN_1900 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_2_io_packet_header_42 = encoders_2_io_valid & proc_2_io_ready ? _GEN_1901 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_2_io_packet_header_43 = encoders_2_io_valid & proc_2_io_ready ? _GEN_1902 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_2_io_packet_header_44 = encoders_2_io_valid & proc_2_io_ready ? _GEN_1903 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_2_io_packet_header_45 = encoders_2_io_valid & proc_2_io_ready ? _GEN_1904 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_2_io_packet_header_46 = encoders_2_io_valid & proc_2_io_ready ? _GEN_1905 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_2_io_packet_header_47 = encoders_2_io_valid & proc_2_io_ready ? _GEN_1906 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_2_io_packet_header_48 = encoders_2_io_valid & proc_2_io_ready ? _GEN_1907 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_2_io_packet_header_49 = encoders_2_io_valid & proc_2_io_ready ? _GEN_1908 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_2_io_packet_header_50 = encoders_2_io_valid & proc_2_io_ready ? _GEN_1909 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_2_io_packet_header_51 = encoders_2_io_valid & proc_2_io_ready ? _GEN_1910 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_2_io_packet_header_52 = encoders_2_io_valid & proc_2_io_ready ? _GEN_1911 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_2_io_packet_header_53 = encoders_2_io_valid & proc_2_io_ready ? _GEN_1912 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_2_io_packet_header_54 = encoders_2_io_valid & proc_2_io_ready ? _GEN_1913 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_2_io_packet_header_55 = encoders_2_io_valid & proc_2_io_ready ? _GEN_1914 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_2_io_packet_header_56 = encoders_2_io_valid & proc_2_io_ready ? _GEN_1915 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_2_io_packet_header_57 = encoders_2_io_valid & proc_2_io_ready ? _GEN_1916 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_2_io_packet_header_58 = encoders_2_io_valid & proc_2_io_ready ? _GEN_1917 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_2_io_packet_header_59 = encoders_2_io_valid & proc_2_io_ready ? _GEN_1918 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_2_io_packet_header_60 = encoders_2_io_valid & proc_2_io_ready ? _GEN_1919 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_2_io_packet_header_61 = encoders_2_io_valid & proc_2_io_ready ? _GEN_1920 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_2_io_packet_header_62 = encoders_2_io_valid & proc_2_io_ready ? _GEN_1921 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_2_io_packet_header_63 = encoders_2_io_valid & proc_2_io_ready ? _GEN_1922 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_2_io_end = encoders_2_io_valid & proc_2_io_ready; // @[controller.scala 89:36]
  assign proc_2_io_mem_rdata = mem_1_io_mem_a_rdata; // @[controller.scala 32:24]
  assign proc_2_io_mod_start = io_mod_proc == 3'h2 & io_mod_start; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 52:34]
  assign proc_2_io_mod_hit_action_addr = io_mod_proc == 3'h2 ? io_mod_hit_action_addr : 32'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 53:44]
  assign proc_2_io_mod_miss_action_addr = io_mod_proc == 3'h2 ? io_mod_miss_action_addr : 32'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 54:45]
  assign proc_2_io_mod_ps_mod_start = io_mod_proc == 3'h2 & io_mod_ps_mod_start; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 55:41]
  assign proc_2_io_mod_ps_mod_header_id = io_mod_proc == 3'h2 & io_mod_ps_mod_header_id; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 56:45]
  assign proc_2_io_mod_ps_mod_header_length = io_mod_proc == 3'h2 ? io_mod_ps_mod_header_length : 32'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 57:49]
  assign proc_2_io_mod_ps_mod_next_tag_start = io_mod_proc == 3'h2 ? io_mod_ps_mod_next_tag_start : 32'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 58:50]
  assign proc_2_io_mod_ps_mod_next_table_0 = io_mod_proc == 3'h2 ? io_mod_ps_mod_next_table_0 : 32'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 61:53]
  assign proc_2_io_mod_ps_mod_next_table_1 = io_mod_proc == 3'h2 ? io_mod_ps_mod_next_table_1 : 32'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 61:53]
  assign proc_2_io_mod_mt_mod_start = io_mod_proc == 3'h2 & io_mod_mt_mod_start; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 63:41]
  assign proc_2_io_mod_mt_mod_header_id = io_mod_proc == 3'h2 ? io_mod_mt_mod_header_id : 4'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 64:45]
  assign proc_2_io_mod_mt_mod_key_off = io_mod_proc == 3'h2 ? io_mod_mt_mod_key_off : 6'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 65:43]
  assign proc_2_io_mod_mt_mod_key_len = io_mod_proc == 3'h2 ? io_mod_mt_mod_key_len : 6'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 66:43]
  assign proc_2_io_mod_mt_mod_val_len = io_mod_proc == 3'h2 ? io_mod_mt_mod_val_len : 6'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 67:43]
  assign proc_2_io_mod_ex_mod_start = io_mod_proc == 3'h2 & io_mod_ex_mod_start; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 68:41]
  assign proc_2_io_mod_ex_mod_ops_0 = io_mod_proc == 3'h2 ? io_mod_ex_mod_ops_0 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_2_io_mod_ex_mod_ops_1 = io_mod_proc == 3'h2 ? io_mod_ex_mod_ops_1 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_2_io_mod_ex_mod_ops_2 = io_mod_proc == 3'h2 ? io_mod_ex_mod_ops_2 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_2_io_mod_ex_mod_ops_3 = io_mod_proc == 3'h2 ? io_mod_ex_mod_ops_3 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_2_io_mod_ex_mod_ops_4 = io_mod_proc == 3'h2 ? io_mod_ex_mod_ops_4 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_2_io_mod_ex_mod_ops_5 = io_mod_proc == 3'h2 ? io_mod_ex_mod_ops_5 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_2_io_mod_ex_mod_ops_6 = io_mod_proc == 3'h2 ? io_mod_ex_mod_ops_6 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_2_io_mod_ex_mod_ops_7 = io_mod_proc == 3'h2 ? io_mod_ex_mod_ops_7 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_2_io_mod_ex_mod_ops_8 = io_mod_proc == 3'h2 ? io_mod_ex_mod_ops_8 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_2_io_mod_ex_mod_ops_9 = io_mod_proc == 3'h2 ? io_mod_ex_mod_ops_9 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_2_io_mod_ex_mod_ops_10 = io_mod_proc == 3'h2 ? io_mod_ex_mod_ops_10 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_2_io_mod_ex_mod_ops_11 = io_mod_proc == 3'h2 ? io_mod_ex_mod_ops_11 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_2_io_mod_ex_mod_ops_12 = io_mod_proc == 3'h2 ? io_mod_ex_mod_ops_12 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_2_io_mod_ex_mod_ops_13 = io_mod_proc == 3'h2 ? io_mod_ex_mod_ops_13 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_2_io_mod_ex_mod_ops_14 = io_mod_proc == 3'h2 ? io_mod_ex_mod_ops_14 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_2_io_mod_ex_mod_ops_15 = io_mod_proc == 3'h2 ? io_mod_ex_mod_ops_15 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_3_clock = clock;
  assign proc_3_reset = reset;
  assign proc_3_io_update = encoders_3_io_valid & proc_3_io_ready; // @[controller.scala 89:36]
  assign proc_3_io_packet_header_0 = encoders_3_io_valid & proc_3_io_ready ? _GEN_2436 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_3_io_packet_header_1 = encoders_3_io_valid & proc_3_io_ready ? _GEN_2437 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_3_io_packet_header_2 = encoders_3_io_valid & proc_3_io_ready ? _GEN_2438 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_3_io_packet_header_3 = encoders_3_io_valid & proc_3_io_ready ? _GEN_2439 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_3_io_packet_header_4 = encoders_3_io_valid & proc_3_io_ready ? _GEN_2440 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_3_io_packet_header_5 = encoders_3_io_valid & proc_3_io_ready ? _GEN_2441 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_3_io_packet_header_6 = encoders_3_io_valid & proc_3_io_ready ? _GEN_2442 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_3_io_packet_header_7 = encoders_3_io_valid & proc_3_io_ready ? _GEN_2443 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_3_io_packet_header_8 = encoders_3_io_valid & proc_3_io_ready ? _GEN_2444 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_3_io_packet_header_9 = encoders_3_io_valid & proc_3_io_ready ? _GEN_2445 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_3_io_packet_header_10 = encoders_3_io_valid & proc_3_io_ready ? _GEN_2446 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_3_io_packet_header_11 = encoders_3_io_valid & proc_3_io_ready ? _GEN_2447 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_3_io_packet_header_12 = encoders_3_io_valid & proc_3_io_ready ? _GEN_2448 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_3_io_packet_header_13 = encoders_3_io_valid & proc_3_io_ready ? _GEN_2449 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_3_io_packet_header_14 = encoders_3_io_valid & proc_3_io_ready ? _GEN_2450 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_3_io_packet_header_15 = encoders_3_io_valid & proc_3_io_ready ? _GEN_2451 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_3_io_packet_header_16 = encoders_3_io_valid & proc_3_io_ready ? _GEN_2452 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_3_io_packet_header_17 = encoders_3_io_valid & proc_3_io_ready ? _GEN_2453 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_3_io_packet_header_18 = encoders_3_io_valid & proc_3_io_ready ? _GEN_2454 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_3_io_packet_header_19 = encoders_3_io_valid & proc_3_io_ready ? _GEN_2455 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_3_io_packet_header_20 = encoders_3_io_valid & proc_3_io_ready ? _GEN_2456 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_3_io_packet_header_21 = encoders_3_io_valid & proc_3_io_ready ? _GEN_2457 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_3_io_packet_header_22 = encoders_3_io_valid & proc_3_io_ready ? _GEN_2458 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_3_io_packet_header_23 = encoders_3_io_valid & proc_3_io_ready ? _GEN_2459 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_3_io_packet_header_24 = encoders_3_io_valid & proc_3_io_ready ? _GEN_2460 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_3_io_packet_header_25 = encoders_3_io_valid & proc_3_io_ready ? _GEN_2461 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_3_io_packet_header_26 = encoders_3_io_valid & proc_3_io_ready ? _GEN_2462 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_3_io_packet_header_27 = encoders_3_io_valid & proc_3_io_ready ? _GEN_2463 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_3_io_packet_header_28 = encoders_3_io_valid & proc_3_io_ready ? _GEN_2464 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_3_io_packet_header_29 = encoders_3_io_valid & proc_3_io_ready ? _GEN_2465 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_3_io_packet_header_30 = encoders_3_io_valid & proc_3_io_ready ? _GEN_2466 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_3_io_packet_header_31 = encoders_3_io_valid & proc_3_io_ready ? _GEN_2467 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_3_io_packet_header_32 = encoders_3_io_valid & proc_3_io_ready ? _GEN_2468 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_3_io_packet_header_33 = encoders_3_io_valid & proc_3_io_ready ? _GEN_2469 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_3_io_packet_header_34 = encoders_3_io_valid & proc_3_io_ready ? _GEN_2470 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_3_io_packet_header_35 = encoders_3_io_valid & proc_3_io_ready ? _GEN_2471 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_3_io_packet_header_36 = encoders_3_io_valid & proc_3_io_ready ? _GEN_2472 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_3_io_packet_header_37 = encoders_3_io_valid & proc_3_io_ready ? _GEN_2473 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_3_io_packet_header_38 = encoders_3_io_valid & proc_3_io_ready ? _GEN_2474 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_3_io_packet_header_39 = encoders_3_io_valid & proc_3_io_ready ? _GEN_2475 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_3_io_packet_header_40 = encoders_3_io_valid & proc_3_io_ready ? _GEN_2476 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_3_io_packet_header_41 = encoders_3_io_valid & proc_3_io_ready ? _GEN_2477 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_3_io_packet_header_42 = encoders_3_io_valid & proc_3_io_ready ? _GEN_2478 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_3_io_packet_header_43 = encoders_3_io_valid & proc_3_io_ready ? _GEN_2479 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_3_io_packet_header_44 = encoders_3_io_valid & proc_3_io_ready ? _GEN_2480 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_3_io_packet_header_45 = encoders_3_io_valid & proc_3_io_ready ? _GEN_2481 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_3_io_packet_header_46 = encoders_3_io_valid & proc_3_io_ready ? _GEN_2482 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_3_io_packet_header_47 = encoders_3_io_valid & proc_3_io_ready ? _GEN_2483 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_3_io_packet_header_48 = encoders_3_io_valid & proc_3_io_ready ? _GEN_2484 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_3_io_packet_header_49 = encoders_3_io_valid & proc_3_io_ready ? _GEN_2485 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_3_io_packet_header_50 = encoders_3_io_valid & proc_3_io_ready ? _GEN_2486 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_3_io_packet_header_51 = encoders_3_io_valid & proc_3_io_ready ? _GEN_2487 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_3_io_packet_header_52 = encoders_3_io_valid & proc_3_io_ready ? _GEN_2488 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_3_io_packet_header_53 = encoders_3_io_valid & proc_3_io_ready ? _GEN_2489 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_3_io_packet_header_54 = encoders_3_io_valid & proc_3_io_ready ? _GEN_2490 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_3_io_packet_header_55 = encoders_3_io_valid & proc_3_io_ready ? _GEN_2491 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_3_io_packet_header_56 = encoders_3_io_valid & proc_3_io_ready ? _GEN_2492 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_3_io_packet_header_57 = encoders_3_io_valid & proc_3_io_ready ? _GEN_2493 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_3_io_packet_header_58 = encoders_3_io_valid & proc_3_io_ready ? _GEN_2494 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_3_io_packet_header_59 = encoders_3_io_valid & proc_3_io_ready ? _GEN_2495 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_3_io_packet_header_60 = encoders_3_io_valid & proc_3_io_ready ? _GEN_2496 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_3_io_packet_header_61 = encoders_3_io_valid & proc_3_io_ready ? _GEN_2497 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_3_io_packet_header_62 = encoders_3_io_valid & proc_3_io_ready ? _GEN_2498 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_3_io_packet_header_63 = encoders_3_io_valid & proc_3_io_ready ? _GEN_2499 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_3_io_end = encoders_3_io_valid & proc_3_io_ready; // @[controller.scala 89:36]
  assign proc_3_io_mem_rdata = mem_1_io_mem_b_rdata; // @[controller.scala 34:24]
  assign proc_3_io_mod_start = io_mod_proc == 3'h3 & io_mod_start; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 52:34]
  assign proc_3_io_mod_hit_action_addr = io_mod_proc == 3'h3 ? io_mod_hit_action_addr : 32'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 53:44]
  assign proc_3_io_mod_miss_action_addr = io_mod_proc == 3'h3 ? io_mod_miss_action_addr : 32'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 54:45]
  assign proc_3_io_mod_ps_mod_start = io_mod_proc == 3'h3 & io_mod_ps_mod_start; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 55:41]
  assign proc_3_io_mod_ps_mod_header_id = io_mod_proc == 3'h3 & io_mod_ps_mod_header_id; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 56:45]
  assign proc_3_io_mod_ps_mod_header_length = io_mod_proc == 3'h3 ? io_mod_ps_mod_header_length : 32'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 57:49]
  assign proc_3_io_mod_ps_mod_next_tag_start = io_mod_proc == 3'h3 ? io_mod_ps_mod_next_tag_start : 32'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 58:50]
  assign proc_3_io_mod_ps_mod_next_table_0 = io_mod_proc == 3'h3 ? io_mod_ps_mod_next_table_0 : 32'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 61:53]
  assign proc_3_io_mod_ps_mod_next_table_1 = io_mod_proc == 3'h3 ? io_mod_ps_mod_next_table_1 : 32'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 61:53]
  assign proc_3_io_mod_mt_mod_start = io_mod_proc == 3'h3 & io_mod_mt_mod_start; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 63:41]
  assign proc_3_io_mod_mt_mod_header_id = io_mod_proc == 3'h3 ? io_mod_mt_mod_header_id : 4'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 64:45]
  assign proc_3_io_mod_mt_mod_key_off = io_mod_proc == 3'h3 ? io_mod_mt_mod_key_off : 6'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 65:43]
  assign proc_3_io_mod_mt_mod_key_len = io_mod_proc == 3'h3 ? io_mod_mt_mod_key_len : 6'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 66:43]
  assign proc_3_io_mod_mt_mod_val_len = io_mod_proc == 3'h3 ? io_mod_mt_mod_val_len : 6'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 67:43]
  assign proc_3_io_mod_ex_mod_start = io_mod_proc == 3'h3 & io_mod_ex_mod_start; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 68:41]
  assign proc_3_io_mod_ex_mod_ops_0 = io_mod_proc == 3'h3 ? io_mod_ex_mod_ops_0 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_3_io_mod_ex_mod_ops_1 = io_mod_proc == 3'h3 ? io_mod_ex_mod_ops_1 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_3_io_mod_ex_mod_ops_2 = io_mod_proc == 3'h3 ? io_mod_ex_mod_ops_2 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_3_io_mod_ex_mod_ops_3 = io_mod_proc == 3'h3 ? io_mod_ex_mod_ops_3 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_3_io_mod_ex_mod_ops_4 = io_mod_proc == 3'h3 ? io_mod_ex_mod_ops_4 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_3_io_mod_ex_mod_ops_5 = io_mod_proc == 3'h3 ? io_mod_ex_mod_ops_5 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_3_io_mod_ex_mod_ops_6 = io_mod_proc == 3'h3 ? io_mod_ex_mod_ops_6 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_3_io_mod_ex_mod_ops_7 = io_mod_proc == 3'h3 ? io_mod_ex_mod_ops_7 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_3_io_mod_ex_mod_ops_8 = io_mod_proc == 3'h3 ? io_mod_ex_mod_ops_8 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_3_io_mod_ex_mod_ops_9 = io_mod_proc == 3'h3 ? io_mod_ex_mod_ops_9 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_3_io_mod_ex_mod_ops_10 = io_mod_proc == 3'h3 ? io_mod_ex_mod_ops_10 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_3_io_mod_ex_mod_ops_11 = io_mod_proc == 3'h3 ? io_mod_ex_mod_ops_11 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_3_io_mod_ex_mod_ops_12 = io_mod_proc == 3'h3 ? io_mod_ex_mod_ops_12 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_3_io_mod_ex_mod_ops_13 = io_mod_proc == 3'h3 ? io_mod_ex_mod_ops_13 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_3_io_mod_ex_mod_ops_14 = io_mod_proc == 3'h3 ? io_mod_ex_mod_ops_14 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_3_io_mod_ex_mod_ops_15 = io_mod_proc == 3'h3 ? io_mod_ex_mod_ops_15 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_4_clock = clock;
  assign proc_4_reset = reset;
  assign proc_4_io_update = encoders_4_io_valid & proc_4_io_ready; // @[controller.scala 89:36]
  assign proc_4_io_packet_header_0 = encoders_4_io_valid & proc_4_io_ready ? _GEN_3013 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_4_io_packet_header_1 = encoders_4_io_valid & proc_4_io_ready ? _GEN_3014 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_4_io_packet_header_2 = encoders_4_io_valid & proc_4_io_ready ? _GEN_3015 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_4_io_packet_header_3 = encoders_4_io_valid & proc_4_io_ready ? _GEN_3016 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_4_io_packet_header_4 = encoders_4_io_valid & proc_4_io_ready ? _GEN_3017 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_4_io_packet_header_5 = encoders_4_io_valid & proc_4_io_ready ? _GEN_3018 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_4_io_packet_header_6 = encoders_4_io_valid & proc_4_io_ready ? _GEN_3019 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_4_io_packet_header_7 = encoders_4_io_valid & proc_4_io_ready ? _GEN_3020 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_4_io_packet_header_8 = encoders_4_io_valid & proc_4_io_ready ? _GEN_3021 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_4_io_packet_header_9 = encoders_4_io_valid & proc_4_io_ready ? _GEN_3022 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_4_io_packet_header_10 = encoders_4_io_valid & proc_4_io_ready ? _GEN_3023 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_4_io_packet_header_11 = encoders_4_io_valid & proc_4_io_ready ? _GEN_3024 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_4_io_packet_header_12 = encoders_4_io_valid & proc_4_io_ready ? _GEN_3025 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_4_io_packet_header_13 = encoders_4_io_valid & proc_4_io_ready ? _GEN_3026 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_4_io_packet_header_14 = encoders_4_io_valid & proc_4_io_ready ? _GEN_3027 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_4_io_packet_header_15 = encoders_4_io_valid & proc_4_io_ready ? _GEN_3028 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_4_io_packet_header_16 = encoders_4_io_valid & proc_4_io_ready ? _GEN_3029 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_4_io_packet_header_17 = encoders_4_io_valid & proc_4_io_ready ? _GEN_3030 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_4_io_packet_header_18 = encoders_4_io_valid & proc_4_io_ready ? _GEN_3031 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_4_io_packet_header_19 = encoders_4_io_valid & proc_4_io_ready ? _GEN_3032 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_4_io_packet_header_20 = encoders_4_io_valid & proc_4_io_ready ? _GEN_3033 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_4_io_packet_header_21 = encoders_4_io_valid & proc_4_io_ready ? _GEN_3034 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_4_io_packet_header_22 = encoders_4_io_valid & proc_4_io_ready ? _GEN_3035 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_4_io_packet_header_23 = encoders_4_io_valid & proc_4_io_ready ? _GEN_3036 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_4_io_packet_header_24 = encoders_4_io_valid & proc_4_io_ready ? _GEN_3037 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_4_io_packet_header_25 = encoders_4_io_valid & proc_4_io_ready ? _GEN_3038 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_4_io_packet_header_26 = encoders_4_io_valid & proc_4_io_ready ? _GEN_3039 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_4_io_packet_header_27 = encoders_4_io_valid & proc_4_io_ready ? _GEN_3040 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_4_io_packet_header_28 = encoders_4_io_valid & proc_4_io_ready ? _GEN_3041 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_4_io_packet_header_29 = encoders_4_io_valid & proc_4_io_ready ? _GEN_3042 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_4_io_packet_header_30 = encoders_4_io_valid & proc_4_io_ready ? _GEN_3043 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_4_io_packet_header_31 = encoders_4_io_valid & proc_4_io_ready ? _GEN_3044 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_4_io_packet_header_32 = encoders_4_io_valid & proc_4_io_ready ? _GEN_3045 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_4_io_packet_header_33 = encoders_4_io_valid & proc_4_io_ready ? _GEN_3046 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_4_io_packet_header_34 = encoders_4_io_valid & proc_4_io_ready ? _GEN_3047 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_4_io_packet_header_35 = encoders_4_io_valid & proc_4_io_ready ? _GEN_3048 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_4_io_packet_header_36 = encoders_4_io_valid & proc_4_io_ready ? _GEN_3049 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_4_io_packet_header_37 = encoders_4_io_valid & proc_4_io_ready ? _GEN_3050 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_4_io_packet_header_38 = encoders_4_io_valid & proc_4_io_ready ? _GEN_3051 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_4_io_packet_header_39 = encoders_4_io_valid & proc_4_io_ready ? _GEN_3052 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_4_io_packet_header_40 = encoders_4_io_valid & proc_4_io_ready ? _GEN_3053 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_4_io_packet_header_41 = encoders_4_io_valid & proc_4_io_ready ? _GEN_3054 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_4_io_packet_header_42 = encoders_4_io_valid & proc_4_io_ready ? _GEN_3055 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_4_io_packet_header_43 = encoders_4_io_valid & proc_4_io_ready ? _GEN_3056 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_4_io_packet_header_44 = encoders_4_io_valid & proc_4_io_ready ? _GEN_3057 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_4_io_packet_header_45 = encoders_4_io_valid & proc_4_io_ready ? _GEN_3058 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_4_io_packet_header_46 = encoders_4_io_valid & proc_4_io_ready ? _GEN_3059 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_4_io_packet_header_47 = encoders_4_io_valid & proc_4_io_ready ? _GEN_3060 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_4_io_packet_header_48 = encoders_4_io_valid & proc_4_io_ready ? _GEN_3061 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_4_io_packet_header_49 = encoders_4_io_valid & proc_4_io_ready ? _GEN_3062 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_4_io_packet_header_50 = encoders_4_io_valid & proc_4_io_ready ? _GEN_3063 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_4_io_packet_header_51 = encoders_4_io_valid & proc_4_io_ready ? _GEN_3064 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_4_io_packet_header_52 = encoders_4_io_valid & proc_4_io_ready ? _GEN_3065 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_4_io_packet_header_53 = encoders_4_io_valid & proc_4_io_ready ? _GEN_3066 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_4_io_packet_header_54 = encoders_4_io_valid & proc_4_io_ready ? _GEN_3067 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_4_io_packet_header_55 = encoders_4_io_valid & proc_4_io_ready ? _GEN_3068 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_4_io_packet_header_56 = encoders_4_io_valid & proc_4_io_ready ? _GEN_3069 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_4_io_packet_header_57 = encoders_4_io_valid & proc_4_io_ready ? _GEN_3070 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_4_io_packet_header_58 = encoders_4_io_valid & proc_4_io_ready ? _GEN_3071 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_4_io_packet_header_59 = encoders_4_io_valid & proc_4_io_ready ? _GEN_3072 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_4_io_packet_header_60 = encoders_4_io_valid & proc_4_io_ready ? _GEN_3073 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_4_io_packet_header_61 = encoders_4_io_valid & proc_4_io_ready ? _GEN_3074 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_4_io_packet_header_62 = encoders_4_io_valid & proc_4_io_ready ? _GEN_3075 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_4_io_packet_header_63 = encoders_4_io_valid & proc_4_io_ready ? _GEN_3076 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_4_io_end = encoders_4_io_valid & proc_4_io_ready; // @[controller.scala 89:36]
  assign proc_4_io_mem_rdata = mem_2_io_mem_a_rdata; // @[controller.scala 32:24]
  assign proc_4_io_mod_start = io_mod_proc == 3'h4 & io_mod_start; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 52:34]
  assign proc_4_io_mod_hit_action_addr = io_mod_proc == 3'h4 ? io_mod_hit_action_addr : 32'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 53:44]
  assign proc_4_io_mod_miss_action_addr = io_mod_proc == 3'h4 ? io_mod_miss_action_addr : 32'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 54:45]
  assign proc_4_io_mod_ps_mod_start = io_mod_proc == 3'h4 & io_mod_ps_mod_start; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 55:41]
  assign proc_4_io_mod_ps_mod_header_id = io_mod_proc == 3'h4 & io_mod_ps_mod_header_id; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 56:45]
  assign proc_4_io_mod_ps_mod_header_length = io_mod_proc == 3'h4 ? io_mod_ps_mod_header_length : 32'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 57:49]
  assign proc_4_io_mod_ps_mod_next_tag_start = io_mod_proc == 3'h4 ? io_mod_ps_mod_next_tag_start : 32'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 58:50]
  assign proc_4_io_mod_ps_mod_next_table_0 = io_mod_proc == 3'h4 ? io_mod_ps_mod_next_table_0 : 32'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 61:53]
  assign proc_4_io_mod_ps_mod_next_table_1 = io_mod_proc == 3'h4 ? io_mod_ps_mod_next_table_1 : 32'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 61:53]
  assign proc_4_io_mod_mt_mod_start = io_mod_proc == 3'h4 & io_mod_mt_mod_start; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 63:41]
  assign proc_4_io_mod_mt_mod_header_id = io_mod_proc == 3'h4 ? io_mod_mt_mod_header_id : 4'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 64:45]
  assign proc_4_io_mod_mt_mod_key_off = io_mod_proc == 3'h4 ? io_mod_mt_mod_key_off : 6'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 65:43]
  assign proc_4_io_mod_mt_mod_key_len = io_mod_proc == 3'h4 ? io_mod_mt_mod_key_len : 6'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 66:43]
  assign proc_4_io_mod_mt_mod_val_len = io_mod_proc == 3'h4 ? io_mod_mt_mod_val_len : 6'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 67:43]
  assign proc_4_io_mod_ex_mod_start = io_mod_proc == 3'h4 & io_mod_ex_mod_start; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 68:41]
  assign proc_4_io_mod_ex_mod_ops_0 = io_mod_proc == 3'h4 ? io_mod_ex_mod_ops_0 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_4_io_mod_ex_mod_ops_1 = io_mod_proc == 3'h4 ? io_mod_ex_mod_ops_1 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_4_io_mod_ex_mod_ops_2 = io_mod_proc == 3'h4 ? io_mod_ex_mod_ops_2 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_4_io_mod_ex_mod_ops_3 = io_mod_proc == 3'h4 ? io_mod_ex_mod_ops_3 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_4_io_mod_ex_mod_ops_4 = io_mod_proc == 3'h4 ? io_mod_ex_mod_ops_4 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_4_io_mod_ex_mod_ops_5 = io_mod_proc == 3'h4 ? io_mod_ex_mod_ops_5 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_4_io_mod_ex_mod_ops_6 = io_mod_proc == 3'h4 ? io_mod_ex_mod_ops_6 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_4_io_mod_ex_mod_ops_7 = io_mod_proc == 3'h4 ? io_mod_ex_mod_ops_7 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_4_io_mod_ex_mod_ops_8 = io_mod_proc == 3'h4 ? io_mod_ex_mod_ops_8 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_4_io_mod_ex_mod_ops_9 = io_mod_proc == 3'h4 ? io_mod_ex_mod_ops_9 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_4_io_mod_ex_mod_ops_10 = io_mod_proc == 3'h4 ? io_mod_ex_mod_ops_10 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_4_io_mod_ex_mod_ops_11 = io_mod_proc == 3'h4 ? io_mod_ex_mod_ops_11 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_4_io_mod_ex_mod_ops_12 = io_mod_proc == 3'h4 ? io_mod_ex_mod_ops_12 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_4_io_mod_ex_mod_ops_13 = io_mod_proc == 3'h4 ? io_mod_ex_mod_ops_13 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_4_io_mod_ex_mod_ops_14 = io_mod_proc == 3'h4 ? io_mod_ex_mod_ops_14 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_4_io_mod_ex_mod_ops_15 = io_mod_proc == 3'h4 ? io_mod_ex_mod_ops_15 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_5_clock = clock;
  assign proc_5_reset = reset;
  assign proc_5_io_update = encoders_5_io_valid & proc_5_io_ready; // @[controller.scala 89:36]
  assign proc_5_io_packet_header_0 = encoders_5_io_valid & proc_5_io_ready ? _GEN_3590 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_5_io_packet_header_1 = encoders_5_io_valid & proc_5_io_ready ? _GEN_3591 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_5_io_packet_header_2 = encoders_5_io_valid & proc_5_io_ready ? _GEN_3592 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_5_io_packet_header_3 = encoders_5_io_valid & proc_5_io_ready ? _GEN_3593 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_5_io_packet_header_4 = encoders_5_io_valid & proc_5_io_ready ? _GEN_3594 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_5_io_packet_header_5 = encoders_5_io_valid & proc_5_io_ready ? _GEN_3595 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_5_io_packet_header_6 = encoders_5_io_valid & proc_5_io_ready ? _GEN_3596 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_5_io_packet_header_7 = encoders_5_io_valid & proc_5_io_ready ? _GEN_3597 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_5_io_packet_header_8 = encoders_5_io_valid & proc_5_io_ready ? _GEN_3598 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_5_io_packet_header_9 = encoders_5_io_valid & proc_5_io_ready ? _GEN_3599 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_5_io_packet_header_10 = encoders_5_io_valid & proc_5_io_ready ? _GEN_3600 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_5_io_packet_header_11 = encoders_5_io_valid & proc_5_io_ready ? _GEN_3601 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_5_io_packet_header_12 = encoders_5_io_valid & proc_5_io_ready ? _GEN_3602 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_5_io_packet_header_13 = encoders_5_io_valid & proc_5_io_ready ? _GEN_3603 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_5_io_packet_header_14 = encoders_5_io_valid & proc_5_io_ready ? _GEN_3604 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_5_io_packet_header_15 = encoders_5_io_valid & proc_5_io_ready ? _GEN_3605 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_5_io_packet_header_16 = encoders_5_io_valid & proc_5_io_ready ? _GEN_3606 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_5_io_packet_header_17 = encoders_5_io_valid & proc_5_io_ready ? _GEN_3607 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_5_io_packet_header_18 = encoders_5_io_valid & proc_5_io_ready ? _GEN_3608 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_5_io_packet_header_19 = encoders_5_io_valid & proc_5_io_ready ? _GEN_3609 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_5_io_packet_header_20 = encoders_5_io_valid & proc_5_io_ready ? _GEN_3610 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_5_io_packet_header_21 = encoders_5_io_valid & proc_5_io_ready ? _GEN_3611 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_5_io_packet_header_22 = encoders_5_io_valid & proc_5_io_ready ? _GEN_3612 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_5_io_packet_header_23 = encoders_5_io_valid & proc_5_io_ready ? _GEN_3613 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_5_io_packet_header_24 = encoders_5_io_valid & proc_5_io_ready ? _GEN_3614 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_5_io_packet_header_25 = encoders_5_io_valid & proc_5_io_ready ? _GEN_3615 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_5_io_packet_header_26 = encoders_5_io_valid & proc_5_io_ready ? _GEN_3616 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_5_io_packet_header_27 = encoders_5_io_valid & proc_5_io_ready ? _GEN_3617 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_5_io_packet_header_28 = encoders_5_io_valid & proc_5_io_ready ? _GEN_3618 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_5_io_packet_header_29 = encoders_5_io_valid & proc_5_io_ready ? _GEN_3619 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_5_io_packet_header_30 = encoders_5_io_valid & proc_5_io_ready ? _GEN_3620 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_5_io_packet_header_31 = encoders_5_io_valid & proc_5_io_ready ? _GEN_3621 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_5_io_packet_header_32 = encoders_5_io_valid & proc_5_io_ready ? _GEN_3622 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_5_io_packet_header_33 = encoders_5_io_valid & proc_5_io_ready ? _GEN_3623 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_5_io_packet_header_34 = encoders_5_io_valid & proc_5_io_ready ? _GEN_3624 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_5_io_packet_header_35 = encoders_5_io_valid & proc_5_io_ready ? _GEN_3625 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_5_io_packet_header_36 = encoders_5_io_valid & proc_5_io_ready ? _GEN_3626 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_5_io_packet_header_37 = encoders_5_io_valid & proc_5_io_ready ? _GEN_3627 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_5_io_packet_header_38 = encoders_5_io_valid & proc_5_io_ready ? _GEN_3628 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_5_io_packet_header_39 = encoders_5_io_valid & proc_5_io_ready ? _GEN_3629 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_5_io_packet_header_40 = encoders_5_io_valid & proc_5_io_ready ? _GEN_3630 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_5_io_packet_header_41 = encoders_5_io_valid & proc_5_io_ready ? _GEN_3631 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_5_io_packet_header_42 = encoders_5_io_valid & proc_5_io_ready ? _GEN_3632 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_5_io_packet_header_43 = encoders_5_io_valid & proc_5_io_ready ? _GEN_3633 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_5_io_packet_header_44 = encoders_5_io_valid & proc_5_io_ready ? _GEN_3634 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_5_io_packet_header_45 = encoders_5_io_valid & proc_5_io_ready ? _GEN_3635 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_5_io_packet_header_46 = encoders_5_io_valid & proc_5_io_ready ? _GEN_3636 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_5_io_packet_header_47 = encoders_5_io_valid & proc_5_io_ready ? _GEN_3637 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_5_io_packet_header_48 = encoders_5_io_valid & proc_5_io_ready ? _GEN_3638 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_5_io_packet_header_49 = encoders_5_io_valid & proc_5_io_ready ? _GEN_3639 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_5_io_packet_header_50 = encoders_5_io_valid & proc_5_io_ready ? _GEN_3640 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_5_io_packet_header_51 = encoders_5_io_valid & proc_5_io_ready ? _GEN_3641 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_5_io_packet_header_52 = encoders_5_io_valid & proc_5_io_ready ? _GEN_3642 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_5_io_packet_header_53 = encoders_5_io_valid & proc_5_io_ready ? _GEN_3643 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_5_io_packet_header_54 = encoders_5_io_valid & proc_5_io_ready ? _GEN_3644 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_5_io_packet_header_55 = encoders_5_io_valid & proc_5_io_ready ? _GEN_3645 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_5_io_packet_header_56 = encoders_5_io_valid & proc_5_io_ready ? _GEN_3646 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_5_io_packet_header_57 = encoders_5_io_valid & proc_5_io_ready ? _GEN_3647 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_5_io_packet_header_58 = encoders_5_io_valid & proc_5_io_ready ? _GEN_3648 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_5_io_packet_header_59 = encoders_5_io_valid & proc_5_io_ready ? _GEN_3649 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_5_io_packet_header_60 = encoders_5_io_valid & proc_5_io_ready ? _GEN_3650 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_5_io_packet_header_61 = encoders_5_io_valid & proc_5_io_ready ? _GEN_3651 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_5_io_packet_header_62 = encoders_5_io_valid & proc_5_io_ready ? _GEN_3652 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_5_io_packet_header_63 = encoders_5_io_valid & proc_5_io_ready ? _GEN_3653 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_5_io_end = encoders_5_io_valid & proc_5_io_ready; // @[controller.scala 89:36]
  assign proc_5_io_mem_rdata = mem_2_io_mem_b_rdata; // @[controller.scala 34:24]
  assign proc_5_io_mod_start = io_mod_proc == 3'h5 & io_mod_start; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 52:34]
  assign proc_5_io_mod_hit_action_addr = io_mod_proc == 3'h5 ? io_mod_hit_action_addr : 32'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 53:44]
  assign proc_5_io_mod_miss_action_addr = io_mod_proc == 3'h5 ? io_mod_miss_action_addr : 32'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 54:45]
  assign proc_5_io_mod_ps_mod_start = io_mod_proc == 3'h5 & io_mod_ps_mod_start; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 55:41]
  assign proc_5_io_mod_ps_mod_header_id = io_mod_proc == 3'h5 & io_mod_ps_mod_header_id; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 56:45]
  assign proc_5_io_mod_ps_mod_header_length = io_mod_proc == 3'h5 ? io_mod_ps_mod_header_length : 32'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 57:49]
  assign proc_5_io_mod_ps_mod_next_tag_start = io_mod_proc == 3'h5 ? io_mod_ps_mod_next_tag_start : 32'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 58:50]
  assign proc_5_io_mod_ps_mod_next_table_0 = io_mod_proc == 3'h5 ? io_mod_ps_mod_next_table_0 : 32'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 61:53]
  assign proc_5_io_mod_ps_mod_next_table_1 = io_mod_proc == 3'h5 ? io_mod_ps_mod_next_table_1 : 32'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 61:53]
  assign proc_5_io_mod_mt_mod_start = io_mod_proc == 3'h5 & io_mod_mt_mod_start; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 63:41]
  assign proc_5_io_mod_mt_mod_header_id = io_mod_proc == 3'h5 ? io_mod_mt_mod_header_id : 4'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 64:45]
  assign proc_5_io_mod_mt_mod_key_off = io_mod_proc == 3'h5 ? io_mod_mt_mod_key_off : 6'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 65:43]
  assign proc_5_io_mod_mt_mod_key_len = io_mod_proc == 3'h5 ? io_mod_mt_mod_key_len : 6'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 66:43]
  assign proc_5_io_mod_mt_mod_val_len = io_mod_proc == 3'h5 ? io_mod_mt_mod_val_len : 6'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 67:43]
  assign proc_5_io_mod_ex_mod_start = io_mod_proc == 3'h5 & io_mod_ex_mod_start; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 68:41]
  assign proc_5_io_mod_ex_mod_ops_0 = io_mod_proc == 3'h5 ? io_mod_ex_mod_ops_0 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_5_io_mod_ex_mod_ops_1 = io_mod_proc == 3'h5 ? io_mod_ex_mod_ops_1 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_5_io_mod_ex_mod_ops_2 = io_mod_proc == 3'h5 ? io_mod_ex_mod_ops_2 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_5_io_mod_ex_mod_ops_3 = io_mod_proc == 3'h5 ? io_mod_ex_mod_ops_3 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_5_io_mod_ex_mod_ops_4 = io_mod_proc == 3'h5 ? io_mod_ex_mod_ops_4 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_5_io_mod_ex_mod_ops_5 = io_mod_proc == 3'h5 ? io_mod_ex_mod_ops_5 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_5_io_mod_ex_mod_ops_6 = io_mod_proc == 3'h5 ? io_mod_ex_mod_ops_6 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_5_io_mod_ex_mod_ops_7 = io_mod_proc == 3'h5 ? io_mod_ex_mod_ops_7 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_5_io_mod_ex_mod_ops_8 = io_mod_proc == 3'h5 ? io_mod_ex_mod_ops_8 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_5_io_mod_ex_mod_ops_9 = io_mod_proc == 3'h5 ? io_mod_ex_mod_ops_9 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_5_io_mod_ex_mod_ops_10 = io_mod_proc == 3'h5 ? io_mod_ex_mod_ops_10 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_5_io_mod_ex_mod_ops_11 = io_mod_proc == 3'h5 ? io_mod_ex_mod_ops_11 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_5_io_mod_ex_mod_ops_12 = io_mod_proc == 3'h5 ? io_mod_ex_mod_ops_12 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_5_io_mod_ex_mod_ops_13 = io_mod_proc == 3'h5 ? io_mod_ex_mod_ops_13 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_5_io_mod_ex_mod_ops_14 = io_mod_proc == 3'h5 ? io_mod_ex_mod_ops_14 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_5_io_mod_ex_mod_ops_15 = io_mod_proc == 3'h5 ? io_mod_ex_mod_ops_15 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_6_clock = clock;
  assign proc_6_reset = reset;
  assign proc_6_io_update = encoders_6_io_valid & proc_6_io_ready; // @[controller.scala 89:36]
  assign proc_6_io_packet_header_0 = encoders_6_io_valid & proc_6_io_ready ? _GEN_4167 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_6_io_packet_header_1 = encoders_6_io_valid & proc_6_io_ready ? _GEN_4168 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_6_io_packet_header_2 = encoders_6_io_valid & proc_6_io_ready ? _GEN_4169 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_6_io_packet_header_3 = encoders_6_io_valid & proc_6_io_ready ? _GEN_4170 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_6_io_packet_header_4 = encoders_6_io_valid & proc_6_io_ready ? _GEN_4171 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_6_io_packet_header_5 = encoders_6_io_valid & proc_6_io_ready ? _GEN_4172 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_6_io_packet_header_6 = encoders_6_io_valid & proc_6_io_ready ? _GEN_4173 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_6_io_packet_header_7 = encoders_6_io_valid & proc_6_io_ready ? _GEN_4174 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_6_io_packet_header_8 = encoders_6_io_valid & proc_6_io_ready ? _GEN_4175 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_6_io_packet_header_9 = encoders_6_io_valid & proc_6_io_ready ? _GEN_4176 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_6_io_packet_header_10 = encoders_6_io_valid & proc_6_io_ready ? _GEN_4177 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_6_io_packet_header_11 = encoders_6_io_valid & proc_6_io_ready ? _GEN_4178 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_6_io_packet_header_12 = encoders_6_io_valid & proc_6_io_ready ? _GEN_4179 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_6_io_packet_header_13 = encoders_6_io_valid & proc_6_io_ready ? _GEN_4180 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_6_io_packet_header_14 = encoders_6_io_valid & proc_6_io_ready ? _GEN_4181 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_6_io_packet_header_15 = encoders_6_io_valid & proc_6_io_ready ? _GEN_4182 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_6_io_packet_header_16 = encoders_6_io_valid & proc_6_io_ready ? _GEN_4183 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_6_io_packet_header_17 = encoders_6_io_valid & proc_6_io_ready ? _GEN_4184 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_6_io_packet_header_18 = encoders_6_io_valid & proc_6_io_ready ? _GEN_4185 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_6_io_packet_header_19 = encoders_6_io_valid & proc_6_io_ready ? _GEN_4186 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_6_io_packet_header_20 = encoders_6_io_valid & proc_6_io_ready ? _GEN_4187 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_6_io_packet_header_21 = encoders_6_io_valid & proc_6_io_ready ? _GEN_4188 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_6_io_packet_header_22 = encoders_6_io_valid & proc_6_io_ready ? _GEN_4189 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_6_io_packet_header_23 = encoders_6_io_valid & proc_6_io_ready ? _GEN_4190 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_6_io_packet_header_24 = encoders_6_io_valid & proc_6_io_ready ? _GEN_4191 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_6_io_packet_header_25 = encoders_6_io_valid & proc_6_io_ready ? _GEN_4192 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_6_io_packet_header_26 = encoders_6_io_valid & proc_6_io_ready ? _GEN_4193 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_6_io_packet_header_27 = encoders_6_io_valid & proc_6_io_ready ? _GEN_4194 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_6_io_packet_header_28 = encoders_6_io_valid & proc_6_io_ready ? _GEN_4195 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_6_io_packet_header_29 = encoders_6_io_valid & proc_6_io_ready ? _GEN_4196 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_6_io_packet_header_30 = encoders_6_io_valid & proc_6_io_ready ? _GEN_4197 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_6_io_packet_header_31 = encoders_6_io_valid & proc_6_io_ready ? _GEN_4198 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_6_io_packet_header_32 = encoders_6_io_valid & proc_6_io_ready ? _GEN_4199 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_6_io_packet_header_33 = encoders_6_io_valid & proc_6_io_ready ? _GEN_4200 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_6_io_packet_header_34 = encoders_6_io_valid & proc_6_io_ready ? _GEN_4201 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_6_io_packet_header_35 = encoders_6_io_valid & proc_6_io_ready ? _GEN_4202 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_6_io_packet_header_36 = encoders_6_io_valid & proc_6_io_ready ? _GEN_4203 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_6_io_packet_header_37 = encoders_6_io_valid & proc_6_io_ready ? _GEN_4204 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_6_io_packet_header_38 = encoders_6_io_valid & proc_6_io_ready ? _GEN_4205 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_6_io_packet_header_39 = encoders_6_io_valid & proc_6_io_ready ? _GEN_4206 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_6_io_packet_header_40 = encoders_6_io_valid & proc_6_io_ready ? _GEN_4207 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_6_io_packet_header_41 = encoders_6_io_valid & proc_6_io_ready ? _GEN_4208 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_6_io_packet_header_42 = encoders_6_io_valid & proc_6_io_ready ? _GEN_4209 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_6_io_packet_header_43 = encoders_6_io_valid & proc_6_io_ready ? _GEN_4210 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_6_io_packet_header_44 = encoders_6_io_valid & proc_6_io_ready ? _GEN_4211 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_6_io_packet_header_45 = encoders_6_io_valid & proc_6_io_ready ? _GEN_4212 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_6_io_packet_header_46 = encoders_6_io_valid & proc_6_io_ready ? _GEN_4213 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_6_io_packet_header_47 = encoders_6_io_valid & proc_6_io_ready ? _GEN_4214 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_6_io_packet_header_48 = encoders_6_io_valid & proc_6_io_ready ? _GEN_4215 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_6_io_packet_header_49 = encoders_6_io_valid & proc_6_io_ready ? _GEN_4216 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_6_io_packet_header_50 = encoders_6_io_valid & proc_6_io_ready ? _GEN_4217 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_6_io_packet_header_51 = encoders_6_io_valid & proc_6_io_ready ? _GEN_4218 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_6_io_packet_header_52 = encoders_6_io_valid & proc_6_io_ready ? _GEN_4219 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_6_io_packet_header_53 = encoders_6_io_valid & proc_6_io_ready ? _GEN_4220 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_6_io_packet_header_54 = encoders_6_io_valid & proc_6_io_ready ? _GEN_4221 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_6_io_packet_header_55 = encoders_6_io_valid & proc_6_io_ready ? _GEN_4222 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_6_io_packet_header_56 = encoders_6_io_valid & proc_6_io_ready ? _GEN_4223 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_6_io_packet_header_57 = encoders_6_io_valid & proc_6_io_ready ? _GEN_4224 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_6_io_packet_header_58 = encoders_6_io_valid & proc_6_io_ready ? _GEN_4225 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_6_io_packet_header_59 = encoders_6_io_valid & proc_6_io_ready ? _GEN_4226 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_6_io_packet_header_60 = encoders_6_io_valid & proc_6_io_ready ? _GEN_4227 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_6_io_packet_header_61 = encoders_6_io_valid & proc_6_io_ready ? _GEN_4228 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_6_io_packet_header_62 = encoders_6_io_valid & proc_6_io_ready ? _GEN_4229 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_6_io_packet_header_63 = encoders_6_io_valid & proc_6_io_ready ? _GEN_4230 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_6_io_end = encoders_6_io_valid & proc_6_io_ready; // @[controller.scala 89:36]
  assign proc_6_io_mem_rdata = mem_3_io_mem_a_rdata; // @[controller.scala 32:24]
  assign proc_6_io_mod_start = io_mod_proc == 3'h6 & io_mod_start; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 52:34]
  assign proc_6_io_mod_hit_action_addr = io_mod_proc == 3'h6 ? io_mod_hit_action_addr : 32'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 53:44]
  assign proc_6_io_mod_miss_action_addr = io_mod_proc == 3'h6 ? io_mod_miss_action_addr : 32'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 54:45]
  assign proc_6_io_mod_ps_mod_start = io_mod_proc == 3'h6 & io_mod_ps_mod_start; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 55:41]
  assign proc_6_io_mod_ps_mod_header_id = io_mod_proc == 3'h6 & io_mod_ps_mod_header_id; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 56:45]
  assign proc_6_io_mod_ps_mod_header_length = io_mod_proc == 3'h6 ? io_mod_ps_mod_header_length : 32'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 57:49]
  assign proc_6_io_mod_ps_mod_next_tag_start = io_mod_proc == 3'h6 ? io_mod_ps_mod_next_tag_start : 32'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 58:50]
  assign proc_6_io_mod_ps_mod_next_table_0 = io_mod_proc == 3'h6 ? io_mod_ps_mod_next_table_0 : 32'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 61:53]
  assign proc_6_io_mod_ps_mod_next_table_1 = io_mod_proc == 3'h6 ? io_mod_ps_mod_next_table_1 : 32'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 61:53]
  assign proc_6_io_mod_mt_mod_start = io_mod_proc == 3'h6 & io_mod_mt_mod_start; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 63:41]
  assign proc_6_io_mod_mt_mod_header_id = io_mod_proc == 3'h6 ? io_mod_mt_mod_header_id : 4'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 64:45]
  assign proc_6_io_mod_mt_mod_key_off = io_mod_proc == 3'h6 ? io_mod_mt_mod_key_off : 6'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 65:43]
  assign proc_6_io_mod_mt_mod_key_len = io_mod_proc == 3'h6 ? io_mod_mt_mod_key_len : 6'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 66:43]
  assign proc_6_io_mod_mt_mod_val_len = io_mod_proc == 3'h6 ? io_mod_mt_mod_val_len : 6'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 67:43]
  assign proc_6_io_mod_ex_mod_start = io_mod_proc == 3'h6 & io_mod_ex_mod_start; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 68:41]
  assign proc_6_io_mod_ex_mod_ops_0 = io_mod_proc == 3'h6 ? io_mod_ex_mod_ops_0 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_6_io_mod_ex_mod_ops_1 = io_mod_proc == 3'h6 ? io_mod_ex_mod_ops_1 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_6_io_mod_ex_mod_ops_2 = io_mod_proc == 3'h6 ? io_mod_ex_mod_ops_2 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_6_io_mod_ex_mod_ops_3 = io_mod_proc == 3'h6 ? io_mod_ex_mod_ops_3 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_6_io_mod_ex_mod_ops_4 = io_mod_proc == 3'h6 ? io_mod_ex_mod_ops_4 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_6_io_mod_ex_mod_ops_5 = io_mod_proc == 3'h6 ? io_mod_ex_mod_ops_5 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_6_io_mod_ex_mod_ops_6 = io_mod_proc == 3'h6 ? io_mod_ex_mod_ops_6 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_6_io_mod_ex_mod_ops_7 = io_mod_proc == 3'h6 ? io_mod_ex_mod_ops_7 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_6_io_mod_ex_mod_ops_8 = io_mod_proc == 3'h6 ? io_mod_ex_mod_ops_8 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_6_io_mod_ex_mod_ops_9 = io_mod_proc == 3'h6 ? io_mod_ex_mod_ops_9 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_6_io_mod_ex_mod_ops_10 = io_mod_proc == 3'h6 ? io_mod_ex_mod_ops_10 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_6_io_mod_ex_mod_ops_11 = io_mod_proc == 3'h6 ? io_mod_ex_mod_ops_11 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_6_io_mod_ex_mod_ops_12 = io_mod_proc == 3'h6 ? io_mod_ex_mod_ops_12 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_6_io_mod_ex_mod_ops_13 = io_mod_proc == 3'h6 ? io_mod_ex_mod_ops_13 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_6_io_mod_ex_mod_ops_14 = io_mod_proc == 3'h6 ? io_mod_ex_mod_ops_14 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_6_io_mod_ex_mod_ops_15 = io_mod_proc == 3'h6 ? io_mod_ex_mod_ops_15 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_7_clock = clock;
  assign proc_7_reset = reset;
  assign proc_7_io_update = encoders_7_io_valid & proc_7_io_ready; // @[controller.scala 89:36]
  assign proc_7_io_packet_header_0 = encoders_7_io_valid & proc_7_io_ready ? _GEN_4744 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_7_io_packet_header_1 = encoders_7_io_valid & proc_7_io_ready ? _GEN_4745 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_7_io_packet_header_2 = encoders_7_io_valid & proc_7_io_ready ? _GEN_4746 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_7_io_packet_header_3 = encoders_7_io_valid & proc_7_io_ready ? _GEN_4747 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_7_io_packet_header_4 = encoders_7_io_valid & proc_7_io_ready ? _GEN_4748 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_7_io_packet_header_5 = encoders_7_io_valid & proc_7_io_ready ? _GEN_4749 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_7_io_packet_header_6 = encoders_7_io_valid & proc_7_io_ready ? _GEN_4750 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_7_io_packet_header_7 = encoders_7_io_valid & proc_7_io_ready ? _GEN_4751 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_7_io_packet_header_8 = encoders_7_io_valid & proc_7_io_ready ? _GEN_4752 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_7_io_packet_header_9 = encoders_7_io_valid & proc_7_io_ready ? _GEN_4753 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_7_io_packet_header_10 = encoders_7_io_valid & proc_7_io_ready ? _GEN_4754 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_7_io_packet_header_11 = encoders_7_io_valid & proc_7_io_ready ? _GEN_4755 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_7_io_packet_header_12 = encoders_7_io_valid & proc_7_io_ready ? _GEN_4756 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_7_io_packet_header_13 = encoders_7_io_valid & proc_7_io_ready ? _GEN_4757 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_7_io_packet_header_14 = encoders_7_io_valid & proc_7_io_ready ? _GEN_4758 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_7_io_packet_header_15 = encoders_7_io_valid & proc_7_io_ready ? _GEN_4759 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_7_io_packet_header_16 = encoders_7_io_valid & proc_7_io_ready ? _GEN_4760 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_7_io_packet_header_17 = encoders_7_io_valid & proc_7_io_ready ? _GEN_4761 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_7_io_packet_header_18 = encoders_7_io_valid & proc_7_io_ready ? _GEN_4762 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_7_io_packet_header_19 = encoders_7_io_valid & proc_7_io_ready ? _GEN_4763 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_7_io_packet_header_20 = encoders_7_io_valid & proc_7_io_ready ? _GEN_4764 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_7_io_packet_header_21 = encoders_7_io_valid & proc_7_io_ready ? _GEN_4765 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_7_io_packet_header_22 = encoders_7_io_valid & proc_7_io_ready ? _GEN_4766 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_7_io_packet_header_23 = encoders_7_io_valid & proc_7_io_ready ? _GEN_4767 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_7_io_packet_header_24 = encoders_7_io_valid & proc_7_io_ready ? _GEN_4768 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_7_io_packet_header_25 = encoders_7_io_valid & proc_7_io_ready ? _GEN_4769 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_7_io_packet_header_26 = encoders_7_io_valid & proc_7_io_ready ? _GEN_4770 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_7_io_packet_header_27 = encoders_7_io_valid & proc_7_io_ready ? _GEN_4771 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_7_io_packet_header_28 = encoders_7_io_valid & proc_7_io_ready ? _GEN_4772 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_7_io_packet_header_29 = encoders_7_io_valid & proc_7_io_ready ? _GEN_4773 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_7_io_packet_header_30 = encoders_7_io_valid & proc_7_io_ready ? _GEN_4774 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_7_io_packet_header_31 = encoders_7_io_valid & proc_7_io_ready ? _GEN_4775 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_7_io_packet_header_32 = encoders_7_io_valid & proc_7_io_ready ? _GEN_4776 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_7_io_packet_header_33 = encoders_7_io_valid & proc_7_io_ready ? _GEN_4777 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_7_io_packet_header_34 = encoders_7_io_valid & proc_7_io_ready ? _GEN_4778 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_7_io_packet_header_35 = encoders_7_io_valid & proc_7_io_ready ? _GEN_4779 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_7_io_packet_header_36 = encoders_7_io_valid & proc_7_io_ready ? _GEN_4780 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_7_io_packet_header_37 = encoders_7_io_valid & proc_7_io_ready ? _GEN_4781 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_7_io_packet_header_38 = encoders_7_io_valid & proc_7_io_ready ? _GEN_4782 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_7_io_packet_header_39 = encoders_7_io_valid & proc_7_io_ready ? _GEN_4783 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_7_io_packet_header_40 = encoders_7_io_valid & proc_7_io_ready ? _GEN_4784 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_7_io_packet_header_41 = encoders_7_io_valid & proc_7_io_ready ? _GEN_4785 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_7_io_packet_header_42 = encoders_7_io_valid & proc_7_io_ready ? _GEN_4786 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_7_io_packet_header_43 = encoders_7_io_valid & proc_7_io_ready ? _GEN_4787 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_7_io_packet_header_44 = encoders_7_io_valid & proc_7_io_ready ? _GEN_4788 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_7_io_packet_header_45 = encoders_7_io_valid & proc_7_io_ready ? _GEN_4789 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_7_io_packet_header_46 = encoders_7_io_valid & proc_7_io_ready ? _GEN_4790 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_7_io_packet_header_47 = encoders_7_io_valid & proc_7_io_ready ? _GEN_4791 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_7_io_packet_header_48 = encoders_7_io_valid & proc_7_io_ready ? _GEN_4792 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_7_io_packet_header_49 = encoders_7_io_valid & proc_7_io_ready ? _GEN_4793 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_7_io_packet_header_50 = encoders_7_io_valid & proc_7_io_ready ? _GEN_4794 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_7_io_packet_header_51 = encoders_7_io_valid & proc_7_io_ready ? _GEN_4795 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_7_io_packet_header_52 = encoders_7_io_valid & proc_7_io_ready ? _GEN_4796 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_7_io_packet_header_53 = encoders_7_io_valid & proc_7_io_ready ? _GEN_4797 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_7_io_packet_header_54 = encoders_7_io_valid & proc_7_io_ready ? _GEN_4798 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_7_io_packet_header_55 = encoders_7_io_valid & proc_7_io_ready ? _GEN_4799 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_7_io_packet_header_56 = encoders_7_io_valid & proc_7_io_ready ? _GEN_4800 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_7_io_packet_header_57 = encoders_7_io_valid & proc_7_io_ready ? _GEN_4801 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_7_io_packet_header_58 = encoders_7_io_valid & proc_7_io_ready ? _GEN_4802 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_7_io_packet_header_59 = encoders_7_io_valid & proc_7_io_ready ? _GEN_4803 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_7_io_packet_header_60 = encoders_7_io_valid & proc_7_io_ready ? _GEN_4804 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_7_io_packet_header_61 = encoders_7_io_valid & proc_7_io_ready ? _GEN_4805 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_7_io_packet_header_62 = encoders_7_io_valid & proc_7_io_ready ? _GEN_4806 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_7_io_packet_header_63 = encoders_7_io_valid & proc_7_io_ready ? _GEN_4807 : 8'h0; // @[controller.scala 89:57 controller.scala 42:41]
  assign proc_7_io_end = encoders_7_io_valid & proc_7_io_ready; // @[controller.scala 89:36]
  assign proc_7_io_mem_rdata = mem_3_io_mem_b_rdata; // @[controller.scala 34:24]
  assign proc_7_io_mod_start = io_mod_proc == 3'h7 & io_mod_start; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 52:34]
  assign proc_7_io_mod_hit_action_addr = io_mod_proc == 3'h7 ? io_mod_hit_action_addr : 32'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 53:44]
  assign proc_7_io_mod_miss_action_addr = io_mod_proc == 3'h7 ? io_mod_miss_action_addr : 32'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 54:45]
  assign proc_7_io_mod_ps_mod_start = io_mod_proc == 3'h7 & io_mod_ps_mod_start; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 55:41]
  assign proc_7_io_mod_ps_mod_header_id = io_mod_proc == 3'h7 & io_mod_ps_mod_header_id; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 56:45]
  assign proc_7_io_mod_ps_mod_header_length = io_mod_proc == 3'h7 ? io_mod_ps_mod_header_length : 32'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 57:49]
  assign proc_7_io_mod_ps_mod_next_tag_start = io_mod_proc == 3'h7 ? io_mod_ps_mod_next_tag_start : 32'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 58:50]
  assign proc_7_io_mod_ps_mod_next_table_0 = io_mod_proc == 3'h7 ? io_mod_ps_mod_next_table_0 : 32'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 61:53]
  assign proc_7_io_mod_ps_mod_next_table_1 = io_mod_proc == 3'h7 ? io_mod_ps_mod_next_table_1 : 32'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 61:53]
  assign proc_7_io_mod_mt_mod_start = io_mod_proc == 3'h7 & io_mod_mt_mod_start; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 63:41]
  assign proc_7_io_mod_mt_mod_header_id = io_mod_proc == 3'h7 ? io_mod_mt_mod_header_id : 4'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 64:45]
  assign proc_7_io_mod_mt_mod_key_off = io_mod_proc == 3'h7 ? io_mod_mt_mod_key_off : 6'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 65:43]
  assign proc_7_io_mod_mt_mod_key_len = io_mod_proc == 3'h7 ? io_mod_mt_mod_key_len : 6'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 66:43]
  assign proc_7_io_mod_mt_mod_val_len = io_mod_proc == 3'h7 ? io_mod_mt_mod_val_len : 6'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 67:43]
  assign proc_7_io_mod_ex_mod_start = io_mod_proc == 3'h7 & io_mod_ex_mod_start; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 68:41]
  assign proc_7_io_mod_ex_mod_ops_0 = io_mod_proc == 3'h7 ? io_mod_ex_mod_ops_0 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_7_io_mod_ex_mod_ops_1 = io_mod_proc == 3'h7 ? io_mod_ex_mod_ops_1 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_7_io_mod_ex_mod_ops_2 = io_mod_proc == 3'h7 ? io_mod_ex_mod_ops_2 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_7_io_mod_ex_mod_ops_3 = io_mod_proc == 3'h7 ? io_mod_ex_mod_ops_3 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_7_io_mod_ex_mod_ops_4 = io_mod_proc == 3'h7 ? io_mod_ex_mod_ops_4 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_7_io_mod_ex_mod_ops_5 = io_mod_proc == 3'h7 ? io_mod_ex_mod_ops_5 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_7_io_mod_ex_mod_ops_6 = io_mod_proc == 3'h7 ? io_mod_ex_mod_ops_6 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_7_io_mod_ex_mod_ops_7 = io_mod_proc == 3'h7 ? io_mod_ex_mod_ops_7 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_7_io_mod_ex_mod_ops_8 = io_mod_proc == 3'h7 ? io_mod_ex_mod_ops_8 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_7_io_mod_ex_mod_ops_9 = io_mod_proc == 3'h7 ? io_mod_ex_mod_ops_9 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_7_io_mod_ex_mod_ops_10 = io_mod_proc == 3'h7 ? io_mod_ex_mod_ops_10 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_7_io_mod_ex_mod_ops_11 = io_mod_proc == 3'h7 ? io_mod_ex_mod_ops_11 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_7_io_mod_ex_mod_ops_12 = io_mod_proc == 3'h7 ? io_mod_ex_mod_ops_12 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_7_io_mod_ex_mod_ops_13 = io_mod_proc == 3'h7 ? io_mod_ex_mod_ops_13 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_7_io_mod_ex_mod_ops_14 = io_mod_proc == 3'h7 ? io_mod_ex_mod_ops_14 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
  assign proc_7_io_mod_ex_mod_ops_15 = io_mod_proc == 3'h7 ? io_mod_ex_mod_ops_15 : 64'h0; // @[controller.scala 49:41 controller.scala 50:28 controller.scala 70:46]
endmodule
